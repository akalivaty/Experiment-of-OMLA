//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 1 1 1 0 0 0 1 0 0 1 1 1 1 1 0 1 0 0 1 1 1 1 0 1 0 0 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n775, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G22gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(G228gat), .A2(G233gat), .ZN(new_n206));
  INV_X1    g005(.A(G141gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT78), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT78), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G141gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n210), .A3(G148gat), .ZN(new_n211));
  INV_X1    g010(.A(G148gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT79), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT79), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G148gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n215), .A3(G141gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n211), .A2(new_n216), .ZN(new_n217));
  AND2_X1   g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219));
  OAI21_X1  g018(.A(KEYINPUT80), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G155gat), .ZN(new_n221));
  INV_X1    g020(.A(G162gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT80), .ZN(new_n224));
  NAND2_X1  g023(.A1(G155gat), .A2(G162gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n220), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT2), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n218), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n217), .A2(new_n227), .A3(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT77), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n225), .B1(new_n219), .B2(new_n232), .ZN(new_n233));
  NOR3_X1   g032(.A1(KEYINPUT77), .A2(G155gat), .A3(G162gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n207), .A2(G148gat), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n212), .A2(G141gat), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n228), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT81), .B(KEYINPUT3), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n231), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT29), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(G211gat), .ZN(new_n244));
  INV_X1    g043(.A(G218gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(G211gat), .A2(G218gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT22), .ZN(new_n249));
  INV_X1    g048(.A(G197gat), .ZN(new_n250));
  INV_X1    g049(.A(G204gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(G197gat), .A2(G204gat), .ZN(new_n253));
  AOI221_X4 g052(.A(KEYINPUT74), .B1(new_n247), .B2(new_n249), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT74), .ZN(new_n255));
  XNOR2_X1  g054(.A(G197gat), .B(G204gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n247), .A2(new_n249), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n248), .B1(new_n254), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n256), .A2(new_n255), .A3(new_n257), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n260), .A2(new_n247), .A3(new_n246), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n243), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT29), .B1(new_n231), .B2(new_n239), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n231), .A2(new_n239), .ZN(new_n266));
  INV_X1    g065(.A(new_n240), .ZN(new_n267));
  AOI22_X1  g066(.A1(new_n265), .A2(new_n262), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n264), .B1(new_n268), .B2(KEYINPUT84), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n265), .A2(new_n262), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n266), .A2(new_n267), .ZN(new_n271));
  AND3_X1   g070(.A1(new_n270), .A2(KEYINPUT84), .A3(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n206), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n266), .A2(KEYINPUT3), .ZN(new_n274));
  INV_X1    g073(.A(new_n206), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n264), .A2(new_n274), .A3(new_n275), .A4(new_n270), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n205), .B1(new_n273), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT85), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n204), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n262), .B1(new_n242), .B2(new_n241), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n270), .A2(new_n271), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT84), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT84), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n275), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n276), .ZN(new_n286));
  OAI21_X1  g085(.A(G22gat), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n273), .A2(new_n205), .A3(new_n276), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n279), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n287), .A2(new_n278), .A3(new_n288), .A4(new_n204), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(G226gat), .ZN(new_n294));
  INV_X1    g093(.A(G233gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(G183gat), .A2(G190gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT26), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(G169gat), .A2(G176gat), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT66), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n298), .B1(new_n301), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G183gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT27), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT27), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G183gat), .ZN(new_n312));
  INV_X1    g111(.A(G190gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n310), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT68), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT28), .ZN(new_n316));
  AND3_X1   g115(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n315), .B1(new_n314), .B2(new_n316), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n310), .A2(new_n312), .A3(KEYINPUT28), .A4(new_n313), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT69), .ZN(new_n321));
  XNOR2_X1  g120(.A(KEYINPUT27), .B(G183gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT69), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n322), .A2(new_n323), .A3(KEYINPUT28), .A4(new_n313), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n308), .B1(new_n319), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G169gat), .ZN(new_n327));
  INV_X1    g126(.A(G176gat), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT23), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n327), .A2(new_n328), .B1(new_n329), .B2(KEYINPUT65), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT65), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT23), .ZN(new_n332));
  AOI22_X1  g131(.A1(new_n330), .A2(new_n332), .B1(new_n304), .B2(new_n305), .ZN(new_n333));
  NOR4_X1   g132(.A1(new_n329), .A2(KEYINPUT64), .A3(G169gat), .A4(G176gat), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT64), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n335), .B1(new_n299), .B2(KEYINPUT23), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT24), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n298), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n309), .A2(new_n313), .ZN(new_n340));
  NAND3_X1  g139(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n333), .A2(new_n337), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT25), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT67), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n298), .B1(new_n345), .B2(KEYINPUT24), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n338), .A2(KEYINPUT67), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n340), .B(new_n341), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n327), .A2(new_n328), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n329), .A2(KEYINPUT65), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(new_n332), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n344), .B1(new_n299), .B2(KEYINPUT23), .ZN(new_n352));
  AND3_X1   g151(.A1(new_n351), .A2(new_n306), .A3(new_n352), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n343), .A2(new_n344), .B1(new_n348), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT75), .B1(new_n326), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT64), .B1(new_n349), .B2(new_n329), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n299), .A2(new_n335), .A3(KEYINPUT23), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n342), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n351), .A2(new_n306), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n344), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n353), .A2(new_n348), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT75), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n321), .A2(new_n324), .ZN(new_n364));
  NOR3_X1   g163(.A1(new_n364), .A2(new_n317), .A3(new_n318), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n362), .B(new_n363), .C1(new_n365), .C2(new_n308), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n297), .B1(new_n355), .B2(new_n366), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n296), .A2(KEYINPUT29), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT76), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n370), .B1(new_n326), .B2(new_n354), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n362), .B(KEYINPUT76), .C1(new_n365), .C2(new_n308), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n369), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n262), .B1(new_n367), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n355), .A2(new_n366), .A3(new_n368), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n371), .A2(new_n296), .A3(new_n372), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(new_n376), .A3(new_n263), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G8gat), .B(G36gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(G64gat), .B(G92gat), .ZN(new_n380));
  XOR2_X1   g179(.A(new_n379), .B(new_n380), .Z(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n374), .A2(new_n377), .A3(new_n381), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(new_n384), .A3(KEYINPUT30), .ZN(new_n385));
  OR3_X1    g184(.A1(new_n378), .A2(KEYINPUT30), .A3(new_n382), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  XOR2_X1   g186(.A(G127gat), .B(G134gat), .Z(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT70), .ZN(new_n389));
  XNOR2_X1  g188(.A(G127gat), .B(G134gat), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT70), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(G113gat), .ZN(new_n393));
  INV_X1    g192(.A(G120gat), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT1), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n396), .B1(G113gat), .B2(G120gat), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n389), .A2(new_n392), .A3(new_n398), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n390), .B(new_n391), .C1(new_n395), .C2(new_n397), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n229), .B1(new_n211), .B2(new_n216), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n402), .A2(new_n227), .B1(new_n238), .B2(new_n235), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n401), .A2(new_n403), .A3(KEYINPUT4), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT4), .B1(new_n401), .B2(new_n403), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(G225gat), .A2(G233gat), .ZN(new_n408));
  AND2_X1   g207(.A1(new_n399), .A2(new_n400), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n274), .A2(new_n409), .A3(new_n241), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n407), .A2(KEYINPUT5), .A3(new_n408), .A4(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n406), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n410), .A2(new_n412), .A3(new_n404), .ZN(new_n413));
  INV_X1    g212(.A(new_n408), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT5), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n401), .B(new_n403), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n416), .B1(new_n417), .B2(new_n414), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n411), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(G1gat), .B(G29gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n420), .B(KEYINPUT0), .ZN(new_n421));
  XNOR2_X1  g220(.A(G57gat), .B(G85gat), .ZN(new_n422));
  XOR2_X1   g221(.A(new_n421), .B(new_n422), .Z(new_n423));
  AOI21_X1  g222(.A(KEYINPUT6), .B1(new_n419), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n418), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n425), .B1(new_n414), .B2(new_n413), .ZN(new_n426));
  INV_X1    g225(.A(new_n423), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n426), .A2(KEYINPUT82), .A3(new_n427), .A4(new_n411), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n411), .B(new_n427), .C1(new_n415), .C2(new_n418), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT82), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n424), .A2(new_n428), .A3(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT6), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT83), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n387), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n437), .B1(new_n387), .B2(new_n436), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n293), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n401), .B1(new_n326), .B2(new_n354), .ZN(new_n442));
  INV_X1    g241(.A(G227gat), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n443), .A2(new_n295), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n362), .B(new_n409), .C1(new_n365), .C2(new_n308), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n442), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT71), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT71), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n442), .A2(new_n445), .A3(new_n448), .A4(new_n444), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XOR2_X1   g249(.A(G15gat), .B(G43gat), .Z(new_n451));
  XNOR2_X1  g250(.A(new_n451), .B(KEYINPUT72), .ZN(new_n452));
  XNOR2_X1  g251(.A(G71gat), .B(G99gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n452), .B(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT33), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT32), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT73), .B1(new_n450), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT73), .ZN(new_n459));
  AOI211_X1 g258(.A(new_n459), .B(new_n456), .C1(new_n447), .C2(new_n449), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT32), .ZN(new_n461));
  AOI22_X1  g260(.A1(new_n447), .A2(new_n449), .B1(new_n461), .B2(KEYINPUT33), .ZN(new_n462));
  OAI22_X1  g261(.A1(new_n458), .A2(new_n460), .B1(new_n462), .B2(new_n454), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT34), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n442), .A2(new_n445), .ZN(new_n465));
  INV_X1    g264(.A(new_n444), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI211_X1 g266(.A(KEYINPUT34), .B(new_n444), .C1(new_n442), .C2(new_n445), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n463), .A2(new_n470), .ZN(new_n471));
  OAI221_X1 g270(.A(new_n469), .B1(new_n462), .B2(new_n454), .C1(new_n458), .C2(new_n460), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT36), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n471), .A2(new_n472), .A3(KEYINPUT36), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n441), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT86), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n423), .B1(new_n419), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n481), .B1(new_n480), .B2(new_n419), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n434), .B1(new_n482), .B2(new_n424), .ZN(new_n483));
  XNOR2_X1  g282(.A(KEYINPUT87), .B(KEYINPUT37), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n382), .B1(new_n378), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n263), .B1(new_n367), .B2(new_n373), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n375), .A2(new_n376), .A3(new_n262), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n486), .A2(KEYINPUT37), .A3(new_n487), .ZN(new_n488));
  OR3_X1    g287(.A1(new_n485), .A2(new_n488), .A3(KEYINPUT38), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n378), .A2(KEYINPUT37), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT38), .B1(new_n490), .B2(new_n485), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n483), .A2(new_n489), .A3(new_n491), .A4(new_n384), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n413), .A2(new_n414), .ZN(new_n493));
  OR2_X1    g292(.A1(new_n493), .A2(KEYINPUT39), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n493), .B(KEYINPUT39), .C1(new_n414), .C2(new_n417), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n494), .A2(new_n495), .A3(new_n423), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n496), .B(KEYINPUT40), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n497), .A2(new_n482), .A3(new_n385), .A4(new_n386), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n492), .A2(new_n292), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT88), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n492), .A2(KEYINPUT88), .A3(new_n292), .A4(new_n498), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n292), .A2(new_n471), .A3(new_n472), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT90), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n387), .A2(new_n436), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(KEYINPUT83), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT90), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n292), .A2(new_n471), .A3(new_n472), .A4(new_n508), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n505), .A2(new_n507), .A3(new_n438), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT35), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n471), .A2(new_n472), .A3(KEYINPUT89), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT89), .B1(new_n471), .B2(new_n472), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT35), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n387), .A2(new_n515), .ZN(new_n516));
  NOR3_X1   g315(.A1(new_n516), .A2(new_n293), .A3(new_n483), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  AOI22_X1  g317(.A1(new_n479), .A2(new_n503), .B1(new_n511), .B2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(G15gat), .B(G22gat), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT16), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n520), .B1(new_n521), .B2(G1gat), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n522), .B(KEYINPUT94), .C1(G1gat), .C2(new_n520), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(G8gat), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n526));
  NOR2_X1   g325(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n527));
  INV_X1    g326(.A(G36gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n529), .A2(KEYINPUT92), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT92), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n531), .B1(new_n527), .B2(new_n528), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n526), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G29gat), .A2(G36gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(G43gat), .B(G50gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT15), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n535), .A2(KEYINPUT15), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n533), .A2(new_n534), .A3(new_n536), .A4(new_n537), .ZN(new_n538));
  AOI22_X1  g337(.A1(new_n529), .A2(new_n526), .B1(G29gat), .B2(G36gat), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n539), .A2(new_n536), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT93), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT17), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT17), .ZN(new_n544));
  AOI211_X1 g343(.A(KEYINPUT93), .B(new_n544), .C1(new_n538), .C2(new_n540), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n525), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(G229gat), .A2(G233gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n524), .A2(new_n541), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT18), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n546), .A2(KEYINPUT18), .A3(new_n547), .A4(new_n548), .ZN(new_n552));
  INV_X1    g351(.A(new_n541), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n525), .A2(KEYINPUT95), .A3(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT95), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(new_n524), .B2(new_n541), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n554), .A2(new_n548), .A3(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n547), .B(KEYINPUT13), .Z(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n551), .A2(new_n552), .A3(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(G113gat), .B(G141gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(KEYINPUT91), .B(G197gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(KEYINPUT11), .B(G169gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT12), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n560), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n551), .A2(new_n552), .A3(new_n559), .A4(new_n566), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  AND2_X1   g370(.A1(G232gat), .A2(G233gat), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n572), .A2(KEYINPUT41), .ZN(new_n573));
  XNOR2_X1  g372(.A(G134gat), .B(G162gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n572), .A2(KEYINPUT41), .ZN(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT99), .B(G92gat), .ZN(new_n578));
  INV_X1    g377(.A(G85gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(G99gat), .A2(G106gat), .ZN(new_n580));
  AOI22_X1  g379(.A1(new_n578), .A2(new_n579), .B1(KEYINPUT8), .B2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT98), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n582), .A2(G85gat), .A3(G92gat), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT7), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OR2_X1    g384(.A1(new_n583), .A2(new_n584), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n581), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(G99gat), .B(G106gat), .Z(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n587), .B(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(new_n541), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(KEYINPUT100), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n543), .A2(new_n545), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n577), .B(new_n591), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G190gat), .B(G218gat), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n595), .B(KEYINPUT101), .Z(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n594), .A2(new_n596), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n576), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(G57gat), .B(G64gat), .Z(new_n601));
  NAND2_X1  g400(.A1(G71gat), .A2(G78gat), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT9), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT96), .ZN(new_n606));
  OR2_X1    g405(.A1(G71gat), .A2(G78gat), .ZN(new_n607));
  AOI22_X1  g406(.A1(new_n606), .A2(new_n604), .B1(new_n607), .B2(new_n602), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  AND2_X1   g408(.A1(new_n607), .A2(new_n602), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n604), .B(new_n601), .C1(new_n610), .C2(new_n606), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n612), .A2(KEYINPUT21), .ZN(new_n613));
  XOR2_X1   g412(.A(G127gat), .B(G155gat), .Z(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n524), .B1(KEYINPUT21), .B2(new_n612), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(G231gat), .A2(G233gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT97), .ZN(new_n619));
  XOR2_X1   g418(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G183gat), .B(G211gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n617), .B(new_n623), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n594), .A2(new_n596), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n625), .A2(new_n597), .A3(new_n575), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n600), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT102), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n600), .A2(new_n626), .A3(new_n624), .A4(KEYINPUT102), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n609), .A2(new_n611), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n588), .A2(KEYINPUT104), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n631), .B1(new_n587), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n633), .B1(new_n587), .B2(new_n632), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT103), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n635), .B1(new_n590), .B2(new_n612), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n587), .B(new_n588), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n637), .A2(KEYINPUT103), .A3(new_n631), .ZN(new_n638));
  XOR2_X1   g437(.A(KEYINPUT105), .B(KEYINPUT10), .Z(new_n639));
  NAND4_X1  g438(.A1(new_n634), .A2(new_n636), .A3(new_n638), .A4(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n590), .A2(KEYINPUT10), .A3(new_n612), .ZN(new_n641));
  AOI21_X1  g440(.A(KEYINPUT106), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(G230gat), .A2(G233gat), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  AND3_X1   g444(.A1(new_n640), .A2(KEYINPUT106), .A3(new_n641), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n634), .A2(new_n636), .A3(new_n638), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(new_n644), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT107), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n649), .A2(KEYINPUT107), .A3(new_n644), .ZN(new_n653));
  XNOR2_X1  g452(.A(G120gat), .B(G148gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(G176gat), .B(G204gat), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n654), .B(new_n655), .Z(new_n656));
  AND3_X1   g455(.A1(new_n652), .A2(new_n653), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n648), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT108), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n640), .A2(new_n641), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(new_n643), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n661), .A2(new_n653), .A3(new_n652), .ZN(new_n662));
  INV_X1    g461(.A(new_n656), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AND3_X1   g463(.A1(new_n658), .A2(new_n659), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n659), .B1(new_n658), .B2(new_n664), .ZN(new_n666));
  OAI211_X1 g465(.A(new_n629), .B(new_n630), .C1(new_n665), .C2(new_n666), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n519), .A2(new_n571), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n436), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(G1gat), .ZN(G1324gat));
  INV_X1    g470(.A(new_n387), .ZN(new_n672));
  XOR2_X1   g471(.A(KEYINPUT16), .B(G8gat), .Z(new_n673));
  NAND3_X1  g472(.A1(new_n668), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n668), .ZN(new_n675));
  OAI21_X1  g474(.A(G8gat), .B1(new_n675), .B2(new_n387), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(new_n674), .ZN(new_n677));
  MUX2_X1   g476(.A(new_n674), .B(new_n677), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g477(.A(G15gat), .B1(new_n675), .B2(new_n477), .ZN(new_n679));
  INV_X1    g478(.A(new_n514), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n680), .A2(G15gat), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n679), .B1(new_n675), .B2(new_n681), .ZN(G1326gat));
  NAND2_X1  g481(.A1(new_n479), .A2(new_n503), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n511), .A2(new_n518), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n685), .A2(new_n293), .A3(new_n570), .ZN(new_n686));
  OR3_X1    g485(.A1(new_n686), .A2(KEYINPUT109), .A3(new_n667), .ZN(new_n687));
  OAI21_X1  g486(.A(KEYINPUT109), .B1(new_n686), .B2(new_n667), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT43), .B(G22gat), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(G1327gat));
  NAND2_X1  g490(.A1(new_n600), .A2(new_n626), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n662), .A2(new_n663), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n646), .A2(new_n642), .A3(new_n644), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n652), .A2(new_n653), .A3(new_n656), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(KEYINPUT108), .B1(new_n694), .B2(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n658), .A2(new_n659), .A3(new_n664), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n701), .A2(new_n624), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(new_n570), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n519), .A2(new_n693), .A3(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n705), .A2(G29gat), .A3(new_n436), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n706), .B(KEYINPUT45), .Z(new_n707));
  INV_X1    g506(.A(KEYINPUT112), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT110), .ZN(new_n709));
  AOI221_X4 g508(.A(new_n709), .B1(new_n514), .B2(new_n517), .C1(new_n510), .C2(KEYINPUT35), .ZN(new_n710));
  AOI21_X1  g509(.A(KEYINPUT110), .B1(new_n511), .B2(new_n518), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n683), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  XOR2_X1   g511(.A(KEYINPUT111), .B(KEYINPUT44), .Z(new_n713));
  NOR2_X1   g512(.A1(new_n693), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(KEYINPUT44), .B1(new_n519), .B2(new_n693), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n703), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n708), .B1(new_n719), .B2(new_n436), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n703), .B1(new_n715), .B2(new_n716), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n721), .A2(KEYINPUT112), .A3(new_n669), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n720), .A2(G29gat), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n723), .ZN(G1328gat));
  OAI21_X1  g523(.A(G36gat), .B1(new_n719), .B2(new_n387), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n672), .A2(new_n528), .ZN(new_n726));
  OAI21_X1  g525(.A(KEYINPUT46), .B1(new_n705), .B2(new_n726), .ZN(new_n727));
  OR3_X1    g526(.A1(new_n705), .A2(KEYINPUT46), .A3(new_n726), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n725), .A2(new_n727), .A3(new_n728), .ZN(G1329gat));
  OAI21_X1  g528(.A(G43gat), .B1(new_n719), .B2(new_n477), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n680), .A2(G43gat), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n685), .A2(new_n692), .A3(new_n718), .A4(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT113), .ZN(new_n734));
  AOI21_X1  g533(.A(KEYINPUT47), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT114), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT114), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n735), .B(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n739), .A2(new_n730), .A3(new_n732), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n737), .A2(new_n740), .ZN(G1330gat));
  OAI21_X1  g540(.A(G50gat), .B1(new_n719), .B2(new_n292), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT48), .ZN(new_n743));
  INV_X1    g542(.A(G50gat), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n702), .A2(new_n744), .A3(new_n692), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n686), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n742), .A2(KEYINPUT115), .A3(new_n743), .A4(new_n747), .ZN(new_n748));
  OR2_X1    g547(.A1(new_n743), .A2(KEYINPUT115), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n743), .A2(KEYINPUT115), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n744), .B1(new_n721), .B2(new_n293), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n749), .B(new_n750), .C1(new_n751), .C2(new_n746), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n748), .A2(new_n752), .ZN(G1331gat));
  AOI21_X1  g552(.A(new_n478), .B1(new_n501), .B2(new_n502), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n684), .A2(new_n709), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n511), .A2(KEYINPUT110), .A3(new_n518), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n629), .A2(new_n630), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n701), .A2(new_n758), .A3(new_n571), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n669), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n672), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n763), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n764));
  XOR2_X1   g563(.A(KEYINPUT49), .B(G64gat), .Z(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(new_n763), .B2(new_n765), .ZN(G1333gat));
  XNOR2_X1  g565(.A(new_n514), .B(KEYINPUT116), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(G71gat), .B1(new_n760), .B2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n477), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n770), .A2(G71gat), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n769), .B1(new_n760), .B2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT50), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n772), .B(new_n773), .ZN(G1334gat));
  NAND2_X1  g573(.A1(new_n760), .A2(new_n293), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g575(.A1(new_n570), .A2(new_n624), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n700), .A2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n780), .B1(new_n715), .B2(new_n716), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(G85gat), .B1(new_n782), .B2(new_n436), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT51), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n778), .A2(new_n693), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n784), .B1(new_n757), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n712), .A2(KEYINPUT51), .A3(new_n785), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n701), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n669), .A2(new_n579), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n783), .B1(new_n790), .B2(new_n791), .ZN(G1336gat));
  AOI21_X1  g591(.A(new_n578), .B1(new_n781), .B2(new_n672), .ZN(new_n793));
  OR3_X1    g592(.A1(new_n700), .A2(G92gat), .A3(new_n387), .ZN(new_n794));
  XOR2_X1   g593(.A(new_n794), .B(KEYINPUT117), .Z(new_n795));
  AOI21_X1  g594(.A(new_n793), .B1(new_n789), .B2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n797));
  INV_X1    g596(.A(new_n789), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n797), .B1(new_n798), .B2(new_n794), .ZN(new_n799));
  OAI22_X1  g598(.A1(new_n796), .A2(new_n797), .B1(new_n799), .B2(new_n793), .ZN(G1337gat));
  OAI21_X1  g599(.A(G99gat), .B1(new_n782), .B2(new_n477), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n680), .A2(G99gat), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n801), .B1(new_n790), .B2(new_n802), .ZN(G1338gat));
  INV_X1    g602(.A(KEYINPUT118), .ZN(new_n804));
  OR2_X1    g603(.A1(new_n804), .A2(KEYINPUT53), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(KEYINPUT53), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n292), .A2(G106gat), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  AOI211_X1 g607(.A(new_n700), .B(new_n808), .C1(new_n787), .C2(new_n788), .ZN(new_n809));
  INV_X1    g608(.A(G106gat), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n810), .B1(new_n781), .B2(new_n293), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n805), .B(new_n806), .C1(new_n809), .C2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n717), .A2(new_n293), .A3(new_n779), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(G106gat), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n789), .A2(new_n701), .A3(new_n807), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n814), .A2(new_n815), .A3(new_n804), .A4(KEYINPUT53), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n812), .A2(new_n816), .ZN(G1339gat));
  INV_X1    g616(.A(KEYINPUT119), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n818), .B1(new_n667), .B2(new_n570), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n758), .A2(KEYINPUT119), .A3(new_n571), .A4(new_n700), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n557), .A2(new_n558), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n547), .B1(new_n546), .B2(new_n548), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n565), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n569), .A2(new_n824), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n692), .A2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n660), .A2(new_n827), .A3(new_n643), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n663), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT54), .B1(new_n660), .B2(new_n643), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n830), .B(KEYINPUT55), .C1(new_n695), .C2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT55), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n831), .B1(new_n645), .B2(new_n647), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n833), .B1(new_n834), .B2(new_n829), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n826), .A2(new_n658), .A3(new_n832), .A4(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n698), .A2(new_n699), .A3(new_n825), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n835), .A2(new_n832), .A3(new_n570), .A4(new_n658), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n693), .B1(new_n839), .B2(KEYINPUT120), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT120), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n841), .B1(new_n837), .B2(new_n838), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n836), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n624), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n821), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n505), .A2(new_n509), .ZN(new_n846));
  NOR4_X1   g645(.A1(new_n845), .A2(new_n436), .A3(new_n672), .A4(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(G113gat), .B1(new_n847), .B2(new_n570), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n669), .A2(new_n387), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n680), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n843), .A2(new_n844), .ZN(new_n852));
  INV_X1    g651(.A(new_n821), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT121), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n854), .A2(new_n855), .A3(new_n292), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT121), .B1(new_n845), .B2(new_n293), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n851), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n571), .A2(new_n393), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n848), .B1(new_n858), .B2(new_n859), .ZN(G1340gat));
  AOI21_X1  g659(.A(G120gat), .B1(new_n847), .B2(new_n701), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n700), .A2(new_n394), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n861), .B1(new_n858), .B2(new_n862), .ZN(G1341gat));
  INV_X1    g662(.A(G127gat), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n847), .A2(new_n864), .A3(new_n624), .ZN(new_n865));
  AOI211_X1 g664(.A(new_n844), .B(new_n851), .C1(new_n856), .C2(new_n857), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n865), .B1(new_n866), .B2(new_n864), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(KEYINPUT122), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT122), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n865), .B(new_n869), .C1(new_n866), .C2(new_n864), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(G1342gat));
  INV_X1    g670(.A(G134gat), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n847), .A2(new_n872), .A3(new_n692), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n873), .A2(KEYINPUT56), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(KEYINPUT56), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n858), .A2(new_n692), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n874), .B(new_n875), .C1(new_n876), .C2(new_n872), .ZN(G1343gat));
  NAND2_X1  g676(.A1(new_n839), .A2(new_n693), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n624), .B1(new_n878), .B2(new_n836), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n293), .B1(new_n821), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(KEYINPUT57), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n770), .A2(new_n849), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT57), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n845), .A2(new_n292), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI22_X1  g685(.A1(new_n886), .A2(new_n570), .B1(new_n208), .B2(new_n210), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n477), .A2(new_n293), .A3(new_n387), .ZN(new_n888));
  AOI211_X1 g687(.A(new_n436), .B(new_n888), .C1(new_n852), .C2(new_n853), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(new_n207), .A3(new_n570), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(KEYINPUT58), .B1(new_n887), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n208), .A2(new_n210), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n885), .A2(new_n884), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n882), .A3(new_n881), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n893), .B1(new_n895), .B2(new_n571), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT58), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n896), .A2(new_n897), .A3(new_n890), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n892), .A2(new_n898), .ZN(G1344gat));
  NAND2_X1  g698(.A1(new_n213), .A2(new_n215), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n889), .A2(new_n901), .A3(new_n701), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT59), .ZN(new_n903));
  OAI21_X1  g702(.A(KEYINPUT57), .B1(new_n845), .B2(new_n292), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT123), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n667), .A2(new_n570), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n884), .B(new_n293), .C1(new_n879), .C2(new_n906), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n770), .A2(new_n700), .A3(new_n849), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n904), .A2(new_n905), .A3(new_n907), .A4(new_n908), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n909), .A2(G148gat), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n904), .A2(new_n907), .A3(new_n908), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(KEYINPUT123), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n903), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  AOI211_X1 g712(.A(KEYINPUT59), .B(new_n901), .C1(new_n886), .C2(new_n701), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n902), .B1(new_n913), .B2(new_n914), .ZN(G1345gat));
  OAI21_X1  g714(.A(G155gat), .B1(new_n895), .B2(new_n844), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n889), .A2(new_n221), .A3(new_n624), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1346gat));
  NAND3_X1  g717(.A1(new_n889), .A2(new_n222), .A3(new_n692), .ZN(new_n919));
  OAI21_X1  g718(.A(KEYINPUT124), .B1(new_n895), .B2(new_n693), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(G162gat), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n895), .A2(KEYINPUT124), .A3(new_n693), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n919), .B1(new_n921), .B2(new_n922), .ZN(G1347gat));
  NOR4_X1   g722(.A1(new_n845), .A2(new_n669), .A3(new_n387), .A4(new_n846), .ZN(new_n924));
  AOI21_X1  g723(.A(G169gat), .B1(new_n924), .B2(new_n570), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n669), .A2(new_n387), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n768), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n927), .B1(new_n856), .B2(new_n857), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n571), .A2(new_n327), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n925), .B1(new_n928), .B2(new_n929), .ZN(G1348gat));
  NOR2_X1   g729(.A1(new_n700), .A2(new_n328), .ZN(new_n931));
  AND3_X1   g730(.A1(new_n928), .A2(KEYINPUT125), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(KEYINPUT125), .B1(new_n928), .B2(new_n931), .ZN(new_n933));
  AOI21_X1  g732(.A(G176gat), .B1(new_n924), .B2(new_n701), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(G1349gat));
  NAND3_X1  g734(.A1(new_n924), .A2(new_n322), .A3(new_n624), .ZN(new_n936));
  AOI211_X1 g735(.A(new_n844), .B(new_n927), .C1(new_n856), .C2(new_n857), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n937), .B2(new_n309), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(KEYINPUT60), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT60), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n936), .B(new_n940), .C1(new_n937), .C2(new_n309), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(G1350gat));
  NAND3_X1  g741(.A1(new_n924), .A2(new_n313), .A3(new_n692), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT61), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n692), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n944), .B1(new_n945), .B2(G190gat), .ZN(new_n946));
  AOI211_X1 g745(.A(KEYINPUT61), .B(new_n313), .C1(new_n928), .C2(new_n692), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(G1351gat));
  NOR2_X1   g747(.A1(new_n845), .A2(new_n669), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n770), .A2(new_n292), .A3(new_n387), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(G197gat), .B1(new_n952), .B2(new_n570), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n477), .A2(new_n926), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n904), .A2(new_n907), .A3(new_n954), .ZN(new_n955));
  NOR3_X1   g754(.A1(new_n955), .A2(new_n250), .A3(new_n571), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n953), .A2(new_n956), .ZN(G1352gat));
  NAND2_X1  g756(.A1(new_n701), .A2(new_n251), .ZN(new_n958));
  OR3_X1    g757(.A1(new_n951), .A2(KEYINPUT62), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g758(.A(G204gat), .B1(new_n955), .B2(new_n700), .ZN(new_n960));
  OAI21_X1  g759(.A(KEYINPUT62), .B1(new_n951), .B2(new_n958), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(G1353gat));
  NAND3_X1  g761(.A1(new_n952), .A2(new_n244), .A3(new_n624), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n904), .A2(new_n624), .A3(new_n907), .A4(new_n954), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(G211gat), .ZN(new_n965));
  NOR2_X1   g764(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g766(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n965), .A2(new_n966), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n963), .B1(new_n969), .B2(new_n970), .ZN(G1354gat));
  OAI21_X1  g770(.A(G218gat), .B1(new_n955), .B2(new_n693), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n692), .A2(new_n245), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n972), .B1(new_n951), .B2(new_n973), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT127), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI211_X1 g775(.A(new_n972), .B(KEYINPUT127), .C1(new_n951), .C2(new_n973), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(G1355gat));
endmodule


