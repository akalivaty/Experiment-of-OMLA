

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743;

  AND2_X1 U366 ( .A1(n360), .A2(n634), .ZN(n345) );
  XNOR2_X2 U367 ( .A(n466), .B(G137), .ZN(n726) );
  XNOR2_X2 U368 ( .A(G131), .B(G134), .ZN(n466) );
  XNOR2_X1 U369 ( .A(n434), .B(n433), .ZN(n626) );
  NOR2_X2 U370 ( .A1(n740), .A2(n742), .ZN(n425) );
  XNOR2_X1 U371 ( .A(n557), .B(KEYINPUT32), .ZN(n739) );
  XNOR2_X1 U372 ( .A(n432), .B(n575), .ZN(n589) );
  AND2_X1 U373 ( .A1(n568), .A2(n569), .ZN(n352) );
  XNOR2_X1 U374 ( .A(n435), .B(KEYINPUT6), .ZN(n601) );
  XNOR2_X1 U375 ( .A(n556), .B(n351), .ZN(n362) );
  XNOR2_X1 U376 ( .A(n491), .B(G472), .ZN(n435) );
  XNOR2_X1 U377 ( .A(n702), .B(n701), .ZN(n703) );
  XNOR2_X1 U378 ( .A(n499), .B(n378), .ZN(n455) );
  XNOR2_X1 U379 ( .A(n381), .B(n531), .ZN(n720) );
  XNOR2_X1 U380 ( .A(n523), .B(n497), .ZN(n381) );
  XOR2_X1 U381 ( .A(G110), .B(KEYINPUT16), .Z(n497) );
  XNOR2_X1 U382 ( .A(n361), .B(n356), .ZN(n740) );
  NOR2_X2 U383 ( .A1(G902), .A2(n695), .ZN(n546) );
  XNOR2_X1 U384 ( .A(n429), .B(KEYINPUT4), .ZN(n428) );
  INV_X1 U385 ( .A(KEYINPUT67), .ZN(n429) );
  AND2_X1 U386 ( .A1(n364), .A2(n656), .ZN(n625) );
  NOR2_X1 U387 ( .A1(G953), .A2(G237), .ZN(n524) );
  XNOR2_X1 U388 ( .A(n726), .B(G146), .ZN(n541) );
  NAND2_X1 U389 ( .A1(n380), .A2(n379), .ZN(n499) );
  OR2_X1 U390 ( .A1(n408), .A2(n437), .ZN(n380) );
  XNOR2_X1 U391 ( .A(n561), .B(KEYINPUT33), .ZN(n687) );
  AND2_X1 U392 ( .A1(n571), .A2(n601), .ZN(n561) );
  XNOR2_X1 U393 ( .A(n369), .B(G478), .ZN(n567) );
  XNOR2_X1 U394 ( .A(n607), .B(KEYINPUT1), .ZN(n674) );
  NAND2_X1 U395 ( .A1(n414), .A2(n413), .ZN(n624) );
  AND2_X1 U396 ( .A1(n419), .A2(n418), .ZN(n414) );
  NOR2_X1 U397 ( .A1(n712), .A2(G902), .ZN(n556) );
  XNOR2_X1 U398 ( .A(n395), .B(KEYINPUT116), .ZN(n678) );
  NAND2_X1 U399 ( .A1(n396), .A2(n435), .ZN(n395) );
  XNOR2_X1 U400 ( .A(n398), .B(n397), .ZN(n396) );
  OR2_X1 U401 ( .A1(G902), .A2(G237), .ZN(n500) );
  INV_X1 U402 ( .A(KEYINPUT48), .ZN(n433) );
  NAND2_X1 U403 ( .A1(n495), .A2(n494), .ZN(n514) );
  INV_X1 U404 ( .A(KEYINPUT77), .ZN(n424) );
  XOR2_X1 U405 ( .A(KEYINPUT66), .B(G101), .Z(n484) );
  XNOR2_X1 U406 ( .A(KEYINPUT86), .B(KEYINPUT84), .ZN(n472) );
  XNOR2_X1 U407 ( .A(n514), .B(n474), .ZN(n473) );
  XNOR2_X1 U408 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n474) );
  AND2_X1 U409 ( .A1(n400), .A2(n399), .ZN(n681) );
  XNOR2_X1 U410 ( .A(n401), .B(KEYINPUT51), .ZN(n400) );
  NOR2_X1 U411 ( .A1(n402), .A2(n680), .ZN(n401) );
  NAND2_X1 U412 ( .A1(n601), .A2(n354), .ZN(n467) );
  XNOR2_X1 U413 ( .A(n541), .B(n431), .ZN(n490) );
  XNOR2_X1 U414 ( .A(n487), .B(n348), .ZN(n431) );
  XNOR2_X1 U415 ( .A(n371), .B(G107), .ZN(n531) );
  INV_X1 U416 ( .A(G122), .ZN(n371) );
  XNOR2_X1 U417 ( .A(n376), .B(n373), .ZN(n372) );
  XNOR2_X1 U418 ( .A(n535), .B(n377), .ZN(n376) );
  XNOR2_X1 U419 ( .A(n375), .B(n374), .ZN(n373) );
  INV_X1 U420 ( .A(G116), .ZN(n377) );
  INV_X1 U421 ( .A(KEYINPUT65), .ZN(n456) );
  NOR2_X1 U422 ( .A1(n577), .A2(KEYINPUT34), .ZN(n451) );
  NOR2_X1 U423 ( .A1(n347), .A2(n407), .ZN(n406) );
  INV_X1 U424 ( .A(n593), .ZN(n452) );
  XNOR2_X1 U425 ( .A(n470), .B(n388), .ZN(n469) );
  INV_X1 U426 ( .A(KEYINPUT22), .ZN(n388) );
  AND2_X1 U427 ( .A1(n611), .A2(n671), .ZN(n540) );
  NAND2_X1 U428 ( .A1(n591), .A2(n390), .ZN(n618) );
  XNOR2_X1 U429 ( .A(n590), .B(n391), .ZN(n390) );
  INV_X1 U430 ( .A(KEYINPUT30), .ZN(n391) );
  AND2_X1 U431 ( .A1(n605), .A2(n673), .ZN(n606) );
  INV_X1 U432 ( .A(KEYINPUT105), .ZN(n363) );
  NAND2_X1 U433 ( .A1(n710), .A2(G472), .ZN(n447) );
  XNOR2_X1 U434 ( .A(n482), .B(n481), .ZN(n712) );
  AND2_X1 U435 ( .A1(n551), .A2(G221), .ZN(n481) );
  XNOR2_X1 U436 ( .A(n483), .B(n550), .ZN(n482) );
  AND2_X1 U437 ( .A1(n440), .A2(n439), .ZN(n689) );
  XNOR2_X1 U438 ( .A(n393), .B(KEYINPUT119), .ZN(n439) );
  NAND2_X1 U439 ( .A1(n394), .A2(n357), .ZN(n393) );
  OR2_X1 U440 ( .A1(n623), .A2(n612), .ZN(n364) );
  OR2_X1 U441 ( .A1(n672), .A2(n671), .ZN(n398) );
  INV_X1 U442 ( .A(KEYINPUT49), .ZN(n397) );
  NOR2_X1 U443 ( .A1(KEYINPUT44), .A2(KEYINPUT83), .ZN(n559) );
  XNOR2_X1 U444 ( .A(n679), .B(n403), .ZN(n402) );
  INV_X1 U445 ( .A(KEYINPUT117), .ZN(n403) );
  NOR2_X1 U446 ( .A1(n441), .A2(n420), .ZN(n383) );
  XNOR2_X1 U447 ( .A(n612), .B(KEYINPUT38), .ZN(n616) );
  NAND2_X1 U448 ( .A1(G234), .A2(G237), .ZN(n504) );
  INV_X1 U449 ( .A(G113), .ZN(n485) );
  XOR2_X1 U450 ( .A(KEYINPUT73), .B(KEYINPUT5), .Z(n486) );
  XNOR2_X1 U451 ( .A(KEYINPUT7), .B(KEYINPUT102), .ZN(n374) );
  XNOR2_X1 U452 ( .A(KEYINPUT9), .B(KEYINPUT101), .ZN(n375) );
  XNOR2_X1 U453 ( .A(KEYINPUT100), .B(G134), .ZN(n535) );
  INV_X1 U454 ( .A(KEYINPUT2), .ZN(n460) );
  INV_X1 U455 ( .A(KEYINPUT74), .ZN(n438) );
  OR2_X1 U456 ( .A1(n616), .A2(n367), .ZN(n666) );
  INV_X1 U457 ( .A(n662), .ZN(n367) );
  INV_X1 U458 ( .A(KEYINPUT39), .ZN(n416) );
  NAND2_X1 U459 ( .A1(n617), .A2(KEYINPUT39), .ZN(n418) );
  XNOR2_X1 U460 ( .A(n368), .B(KEYINPUT104), .ZN(n611) );
  NOR2_X1 U461 ( .A1(n568), .A2(n567), .ZN(n368) );
  INV_X1 U462 ( .A(KEYINPUT107), .ZN(n588) );
  XNOR2_X1 U463 ( .A(n600), .B(n389), .ZN(n605) );
  INV_X1 U464 ( .A(KEYINPUT70), .ZN(n389) );
  XNOR2_X1 U465 ( .A(G116), .B(KEYINPUT3), .ZN(n488) );
  XOR2_X1 U466 ( .A(G119), .B(KEYINPUT72), .Z(n489) );
  XNOR2_X1 U467 ( .A(n582), .B(n454), .ZN(n453) );
  INV_X1 U468 ( .A(KEYINPUT45), .ZN(n454) );
  XNOR2_X1 U469 ( .A(G128), .B(G119), .ZN(n547) );
  XNOR2_X1 U470 ( .A(n392), .B(G110), .ZN(n548) );
  INV_X1 U471 ( .A(G137), .ZN(n392) );
  XNOR2_X1 U472 ( .A(G143), .B(KEYINPUT97), .ZN(n519) );
  XOR2_X1 U473 ( .A(KEYINPUT98), .B(KEYINPUT96), .Z(n520) );
  XNOR2_X1 U474 ( .A(G122), .B(G131), .ZN(n517) );
  XOR2_X1 U475 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n518) );
  XNOR2_X1 U476 ( .A(n525), .B(n427), .ZN(n426) );
  INV_X1 U477 ( .A(KEYINPUT99), .ZN(n427) );
  XNOR2_X1 U478 ( .A(n543), .B(n423), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n544), .B(n424), .ZN(n423) );
  XNOR2_X1 U480 ( .A(n720), .B(n498), .ZN(n378) );
  XNOR2_X1 U481 ( .A(n473), .B(n471), .ZN(n498) );
  XNOR2_X1 U482 ( .A(n496), .B(n472), .ZN(n471) );
  OR2_X1 U483 ( .A1(n684), .A2(n685), .ZN(n394) );
  INV_X1 U484 ( .A(n467), .ZN(n619) );
  XNOR2_X1 U485 ( .A(n366), .B(KEYINPUT41), .ZN(n686) );
  NOR2_X1 U486 ( .A1(n666), .A2(n665), .ZN(n366) );
  XNOR2_X1 U487 ( .A(n467), .B(n412), .ZN(n411) );
  INV_X1 U488 ( .A(KEYINPUT110), .ZN(n412) );
  INV_X1 U489 ( .A(KEYINPUT0), .ZN(n512) );
  INV_X1 U490 ( .A(KEYINPUT94), .ZN(n575) );
  AND2_X1 U491 ( .A1(n607), .A2(n671), .ZN(n475) );
  AND2_X1 U492 ( .A1(n469), .A2(n387), .ZN(n565) );
  XNOR2_X1 U493 ( .A(n442), .B(n536), .ZN(n708) );
  XNOR2_X1 U494 ( .A(n372), .B(n370), .ZN(n442) );
  NAND2_X1 U495 ( .A1(n624), .A2(n352), .ZN(n361) );
  NOR2_X1 U496 ( .A1(n603), .A2(n387), .ZN(n654) );
  XNOR2_X1 U497 ( .A(n409), .B(KEYINPUT36), .ZN(n603) );
  NAND2_X1 U498 ( .A1(n411), .A2(n410), .ZN(n409) );
  INV_X1 U499 ( .A(n602), .ZN(n410) );
  INV_X1 U500 ( .A(KEYINPUT35), .ZN(n404) );
  NAND2_X1 U501 ( .A1(n451), .A2(n450), .ZN(n449) );
  NAND2_X1 U502 ( .A1(n469), .A2(n468), .ZN(n557) );
  NOR2_X1 U503 ( .A1(n613), .A2(n609), .ZN(n647) );
  NAND2_X1 U504 ( .A1(n446), .A2(n634), .ZN(n445) );
  XNOR2_X1 U505 ( .A(n447), .B(n633), .ZN(n446) );
  NAND2_X1 U506 ( .A1(n479), .A2(n634), .ZN(n478) );
  XNOR2_X1 U507 ( .A(n480), .B(n358), .ZN(n479) );
  NOR2_X1 U508 ( .A1(G953), .A2(n690), .ZN(n691) );
  INV_X1 U509 ( .A(n364), .ZN(n657) );
  XNOR2_X1 U510 ( .A(n502), .B(n501), .ZN(n346) );
  AND2_X1 U511 ( .A1(n687), .A2(KEYINPUT34), .ZN(n347) );
  AND2_X1 U512 ( .A1(G210), .A2(n524), .ZN(n348) );
  INV_X1 U513 ( .A(n435), .ZN(n673) );
  INV_X1 U514 ( .A(n674), .ZN(n387) );
  XOR2_X1 U515 ( .A(KEYINPUT24), .B(KEYINPUT92), .Z(n349) );
  XOR2_X1 U516 ( .A(G110), .B(G107), .Z(n350) );
  XNOR2_X1 U517 ( .A(n555), .B(n554), .ZN(n351) );
  OR2_X1 U518 ( .A1(n387), .A2(n672), .ZN(n353) );
  AND2_X1 U519 ( .A1(n605), .A2(n352), .ZN(n354) );
  AND2_X1 U520 ( .A1(n625), .A2(KEYINPUT2), .ZN(n355) );
  XNOR2_X1 U521 ( .A(KEYINPUT40), .B(KEYINPUT109), .ZN(n356) );
  OR2_X1 U522 ( .A1(n687), .A2(n686), .ZN(n357) );
  XOR2_X1 U523 ( .A(n712), .B(n711), .Z(n358) );
  XNOR2_X1 U524 ( .A(G902), .B(KEYINPUT15), .ZN(n537) );
  XNOR2_X1 U525 ( .A(n693), .B(n692), .ZN(n359) );
  XNOR2_X1 U526 ( .A(n694), .B(n359), .ZN(n360) );
  XNOR2_X1 U527 ( .A(n541), .B(n422), .ZN(n421) );
  XNOR2_X1 U528 ( .A(n729), .B(n438), .ZN(n461) );
  INV_X1 U529 ( .A(n362), .ZN(n476) );
  NAND2_X1 U530 ( .A1(n362), .A2(n599), .ZN(n600) );
  AND2_X1 U531 ( .A1(n476), .A2(n671), .ZN(n675) );
  AND2_X1 U532 ( .A1(n435), .A2(n362), .ZN(n558) );
  XNOR2_X1 U533 ( .A(n476), .B(n363), .ZN(n672) );
  XNOR2_X2 U534 ( .A(n365), .B(n428), .ZN(n727) );
  XNOR2_X1 U535 ( .A(n365), .B(n531), .ZN(n370) );
  XNOR2_X2 U536 ( .A(n430), .B(G128), .ZN(n365) );
  INV_X1 U537 ( .A(n616), .ZN(n661) );
  OR2_X1 U538 ( .A1(n708), .A2(G902), .ZN(n369) );
  NAND2_X1 U539 ( .A1(n408), .A2(n437), .ZN(n379) );
  XNOR2_X2 U540 ( .A(n727), .B(n484), .ZN(n408) );
  NAND2_X1 U541 ( .A1(n384), .A2(n382), .ZN(n628) );
  NAND2_X1 U542 ( .A1(n383), .A2(n714), .ZN(n382) );
  NAND2_X1 U543 ( .A1(n385), .A2(n420), .ZN(n384) );
  NAND2_X1 U544 ( .A1(n386), .A2(n714), .ZN(n385) );
  XNOR2_X2 U545 ( .A(n583), .B(n453), .ZN(n714) );
  INV_X1 U546 ( .A(n441), .ZN(n386) );
  NAND2_X1 U547 ( .A1(n608), .A2(n607), .ZN(n613) );
  NOR2_X1 U548 ( .A1(n654), .A2(n464), .ZN(n463) );
  XNOR2_X1 U549 ( .A(n549), .B(n349), .ZN(n436) );
  XNOR2_X1 U550 ( .A(n552), .B(n436), .ZN(n483) );
  XOR2_X1 U551 ( .A(KEYINPUT47), .B(n610), .Z(n465) );
  NAND2_X1 U552 ( .A1(n612), .A2(n662), .ZN(n597) );
  XNOR2_X1 U553 ( .A(n499), .B(n490), .ZN(n630) );
  NAND2_X1 U554 ( .A1(n417), .A2(n415), .ZN(n413) );
  NAND2_X1 U555 ( .A1(n581), .A2(n580), .ZN(n583) );
  NAND2_X1 U556 ( .A1(n448), .A2(n452), .ZN(n407) );
  NAND2_X1 U557 ( .A1(n449), .A2(n406), .ZN(n405) );
  INV_X1 U558 ( .A(n686), .ZN(n399) );
  OR2_X2 U559 ( .A1(n738), .A2(KEYINPUT44), .ZN(n563) );
  XNOR2_X2 U560 ( .A(n405), .B(n404), .ZN(n738) );
  XNOR2_X1 U561 ( .A(n408), .B(n421), .ZN(n695) );
  AND2_X2 U562 ( .A1(n626), .A2(n625), .ZN(n729) );
  NAND2_X1 U563 ( .A1(n626), .A2(n355), .ZN(n441) );
  AND2_X1 U564 ( .A1(n477), .A2(n416), .ZN(n415) );
  INV_X1 U565 ( .A(n618), .ZN(n417) );
  NAND2_X1 U566 ( .A1(n618), .A2(KEYINPUT39), .ZN(n419) );
  INV_X1 U567 ( .A(KEYINPUT75), .ZN(n420) );
  XNOR2_X1 U568 ( .A(n425), .B(KEYINPUT46), .ZN(n462) );
  NAND2_X1 U569 ( .A1(n461), .A2(n460), .ZN(n459) );
  XOR2_X2 U570 ( .A(G113), .B(G104), .Z(n523) );
  NAND2_X1 U571 ( .A1(n462), .A2(n463), .ZN(n434) );
  INV_X1 U572 ( .A(n611), .ZN(n665) );
  XNOR2_X1 U573 ( .A(n426), .B(n523), .ZN(n526) );
  INV_X2 U574 ( .A(G143), .ZN(n430) );
  NAND2_X1 U575 ( .A1(n475), .A2(n476), .ZN(n432) );
  INV_X1 U576 ( .A(n719), .ZN(n437) );
  NAND2_X1 U577 ( .A1(n459), .A2(n629), .ZN(n458) );
  INV_X1 U578 ( .A(n617), .ZN(n477) );
  XNOR2_X1 U579 ( .A(n345), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U580 ( .A1(n739), .A2(n644), .ZN(n560) );
  XNOR2_X1 U581 ( .A(n660), .B(KEYINPUT81), .ZN(n440) );
  XNOR2_X1 U582 ( .A(n445), .B(KEYINPUT63), .ZN(G57) );
  INV_X1 U583 ( .A(n443), .ZN(n667) );
  NAND2_X1 U584 ( .A1(n647), .A2(n443), .ZN(n610) );
  OR2_X1 U585 ( .A1(n651), .A2(n352), .ZN(n443) );
  XNOR2_X1 U586 ( .A(n444), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X2 U587 ( .A1(n705), .A2(n713), .ZN(n444) );
  XNOR2_X1 U588 ( .A(n534), .B(KEYINPUT80), .ZN(n551) );
  NAND2_X1 U589 ( .A1(n465), .A2(n741), .ZN(n464) );
  NAND2_X1 U590 ( .A1(n577), .A2(KEYINPUT34), .ZN(n448) );
  INV_X1 U591 ( .A(n687), .ZN(n450) );
  XNOR2_X2 U592 ( .A(n573), .B(KEYINPUT91), .ZN(n577) );
  NOR2_X2 U593 ( .A1(n455), .A2(n629), .ZN(n503) );
  XNOR2_X1 U594 ( .A(n455), .B(KEYINPUT79), .ZN(n692) );
  XNOR2_X2 U595 ( .A(n457), .B(n456), .ZN(n710) );
  NOR2_X2 U596 ( .A1(n659), .A2(n458), .ZN(n457) );
  NAND2_X1 U597 ( .A1(n628), .A2(n627), .ZN(n659) );
  XNOR2_X2 U598 ( .A(n546), .B(n545), .ZN(n607) );
  INV_X1 U599 ( .A(n612), .ZN(n592) );
  XNOR2_X2 U600 ( .A(n597), .B(KEYINPUT19), .ZN(n604) );
  XNOR2_X2 U601 ( .A(n503), .B(n346), .ZN(n612) );
  NOR2_X1 U602 ( .A1(n601), .A2(n353), .ZN(n468) );
  NAND2_X1 U603 ( .A1(n573), .A2(n540), .ZN(n470) );
  XNOR2_X1 U604 ( .A(n589), .B(n588), .ZN(n591) );
  XNOR2_X1 U605 ( .A(n478), .B(KEYINPUT125), .ZN(G66) );
  NAND2_X1 U606 ( .A1(n710), .A2(G217), .ZN(n480) );
  XNOR2_X2 U607 ( .A(n516), .B(n515), .ZN(n550) );
  BUF_X1 U608 ( .A(n710), .Z(n706) );
  XNOR2_X1 U609 ( .A(n486), .B(n485), .ZN(n487) );
  INV_X1 U610 ( .A(n713), .ZN(n634) );
  XNOR2_X1 U611 ( .A(n704), .B(n703), .ZN(n705) );
  NOR2_X1 U612 ( .A1(G952), .A2(n730), .ZN(n713) );
  XNOR2_X1 U613 ( .A(n489), .B(n488), .ZN(n719) );
  NOR2_X1 U614 ( .A1(n630), .A2(G902), .ZN(n491) );
  NAND2_X1 U615 ( .A1(G214), .A2(n500), .ZN(n662) );
  INV_X1 U616 ( .A(n537), .ZN(n629) );
  INV_X1 U617 ( .A(G146), .ZN(n492) );
  NAND2_X1 U618 ( .A1(G125), .A2(n492), .ZN(n495) );
  INV_X1 U619 ( .A(G125), .ZN(n493) );
  NAND2_X1 U620 ( .A1(n493), .A2(G146), .ZN(n494) );
  INV_X2 U621 ( .A(G953), .ZN(n730) );
  NAND2_X1 U622 ( .A1(G224), .A2(n730), .ZN(n496) );
  XOR2_X1 U623 ( .A(KEYINPUT78), .B(KEYINPUT87), .Z(n502) );
  NAND2_X1 U624 ( .A1(G210), .A2(n500), .ZN(n501) );
  XNOR2_X1 U625 ( .A(n504), .B(KEYINPUT14), .ZN(n506) );
  NAND2_X1 U626 ( .A1(G952), .A2(n506), .ZN(n505) );
  XNOR2_X1 U627 ( .A(n505), .B(KEYINPUT88), .ZN(n685) );
  NOR2_X1 U628 ( .A1(G953), .A2(n685), .ZN(n587) );
  INV_X1 U629 ( .A(n587), .ZN(n509) );
  NAND2_X1 U630 ( .A1(n506), .A2(G902), .ZN(n507) );
  XNOR2_X1 U631 ( .A(n507), .B(KEYINPUT89), .ZN(n584) );
  NOR2_X1 U632 ( .A1(G898), .A2(n730), .ZN(n723) );
  NAND2_X1 U633 ( .A1(n584), .A2(n723), .ZN(n508) );
  NAND2_X1 U634 ( .A1(n509), .A2(n508), .ZN(n510) );
  XNOR2_X1 U635 ( .A(KEYINPUT90), .B(n510), .ZN(n511) );
  NAND2_X1 U636 ( .A1(n604), .A2(n511), .ZN(n513) );
  XNOR2_X2 U637 ( .A(n513), .B(n512), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n514), .B(G140), .ZN(n516) );
  XOR2_X1 U639 ( .A(KEYINPUT69), .B(KEYINPUT10), .Z(n515) );
  XNOR2_X1 U640 ( .A(n518), .B(n517), .ZN(n522) );
  XNOR2_X1 U641 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U642 ( .A(n522), .B(n521), .ZN(n527) );
  NAND2_X1 U643 ( .A1(n524), .A2(G214), .ZN(n525) );
  XNOR2_X1 U644 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U645 ( .A(n550), .B(n528), .ZN(n702) );
  NOR2_X1 U646 ( .A1(G902), .A2(n702), .ZN(n530) );
  XNOR2_X1 U647 ( .A(KEYINPUT13), .B(G475), .ZN(n529) );
  XNOR2_X1 U648 ( .A(n530), .B(n529), .ZN(n568) );
  XOR2_X1 U649 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n533) );
  NAND2_X1 U650 ( .A1(G234), .A2(n730), .ZN(n532) );
  XNOR2_X1 U651 ( .A(n533), .B(n532), .ZN(n534) );
  NAND2_X1 U652 ( .A1(n551), .A2(G217), .ZN(n536) );
  NAND2_X1 U653 ( .A1(G234), .A2(n537), .ZN(n538) );
  XNOR2_X1 U654 ( .A(KEYINPUT20), .B(n538), .ZN(n553) );
  NAND2_X1 U655 ( .A1(n553), .A2(G221), .ZN(n539) );
  XOR2_X1 U656 ( .A(n539), .B(KEYINPUT21), .Z(n671) );
  XNOR2_X1 U657 ( .A(G140), .B(G104), .ZN(n542) );
  XNOR2_X1 U658 ( .A(n350), .B(n542), .ZN(n543) );
  NAND2_X1 U659 ( .A1(G227), .A2(n730), .ZN(n544) );
  XNOR2_X1 U660 ( .A(KEYINPUT71), .B(G469), .ZN(n545) );
  XNOR2_X1 U661 ( .A(n548), .B(n547), .ZN(n552) );
  XOR2_X1 U662 ( .A(KEYINPUT93), .B(KEYINPUT23), .Z(n549) );
  XOR2_X1 U663 ( .A(KEYINPUT76), .B(KEYINPUT25), .Z(n555) );
  NAND2_X1 U664 ( .A1(n553), .A2(G217), .ZN(n554) );
  NAND2_X1 U665 ( .A1(n565), .A2(n558), .ZN(n644) );
  XNOR2_X1 U666 ( .A(n560), .B(n559), .ZN(n562) );
  NAND2_X1 U667 ( .A1(n568), .A2(n567), .ZN(n593) );
  INV_X1 U668 ( .A(n671), .ZN(n598) );
  AND2_X1 U669 ( .A1(n674), .A2(n675), .ZN(n571) );
  NAND2_X1 U670 ( .A1(n562), .A2(n738), .ZN(n564) );
  NAND2_X1 U671 ( .A1(n564), .A2(n563), .ZN(n581) );
  NAND2_X1 U672 ( .A1(n672), .A2(n565), .ZN(n566) );
  NOR2_X1 U673 ( .A1(n601), .A2(n566), .ZN(n635) );
  INV_X1 U674 ( .A(n567), .ZN(n569) );
  NOR2_X1 U675 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U676 ( .A(n570), .B(KEYINPUT103), .Z(n651) );
  NAND2_X1 U677 ( .A1(n571), .A2(n673), .ZN(n572) );
  XNOR2_X1 U678 ( .A(n572), .B(KEYINPUT95), .ZN(n680) );
  NAND2_X1 U679 ( .A1(n573), .A2(n680), .ZN(n574) );
  XNOR2_X1 U680 ( .A(n574), .B(KEYINPUT31), .ZN(n652) );
  NAND2_X1 U681 ( .A1(n435), .A2(n589), .ZN(n576) );
  NOR2_X1 U682 ( .A1(n577), .A2(n576), .ZN(n637) );
  NOR2_X1 U683 ( .A1(n652), .A2(n637), .ZN(n578) );
  NOR2_X1 U684 ( .A1(n667), .A2(n578), .ZN(n579) );
  NOR2_X1 U685 ( .A1(n635), .A2(n579), .ZN(n580) );
  XOR2_X1 U686 ( .A(KEYINPUT64), .B(KEYINPUT82), .Z(n582) );
  NAND2_X1 U687 ( .A1(G953), .A2(n584), .ZN(n585) );
  NOR2_X1 U688 ( .A1(G900), .A2(n585), .ZN(n586) );
  NOR2_X1 U689 ( .A1(n587), .A2(n586), .ZN(n615) );
  NAND2_X1 U690 ( .A1(n662), .A2(n673), .ZN(n590) );
  NOR2_X1 U691 ( .A1(n615), .A2(n618), .ZN(n595) );
  NOR2_X1 U692 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U693 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U694 ( .A(KEYINPUT108), .B(n596), .ZN(n741) );
  BUF_X1 U695 ( .A(n597), .Z(n602) );
  NOR2_X1 U696 ( .A1(n598), .A2(n615), .ZN(n599) );
  INV_X1 U697 ( .A(n604), .ZN(n609) );
  XNOR2_X1 U698 ( .A(KEYINPUT28), .B(n606), .ZN(n608) );
  NOR2_X1 U699 ( .A1(n613), .A2(n686), .ZN(n614) );
  XNOR2_X1 U700 ( .A(n614), .B(KEYINPUT42), .ZN(n742) );
  OR2_X1 U701 ( .A1(n616), .A2(n615), .ZN(n617) );
  NAND2_X1 U702 ( .A1(n619), .A2(n662), .ZN(n620) );
  XNOR2_X1 U703 ( .A(KEYINPUT106), .B(n620), .ZN(n621) );
  NOR2_X1 U704 ( .A1(n674), .A2(n621), .ZN(n622) );
  XNOR2_X1 U705 ( .A(n622), .B(KEYINPUT43), .ZN(n623) );
  NAND2_X1 U706 ( .A1(n651), .A2(n624), .ZN(n656) );
  OR2_X1 U707 ( .A1(n714), .A2(KEYINPUT2), .ZN(n627) );
  XOR2_X1 U708 ( .A(KEYINPUT111), .B(KEYINPUT62), .Z(n632) );
  XNOR2_X1 U709 ( .A(n630), .B(KEYINPUT85), .ZN(n631) );
  XNOR2_X1 U710 ( .A(n632), .B(n631), .ZN(n633) );
  XOR2_X1 U711 ( .A(G101), .B(n635), .Z(G3) );
  NAND2_X1 U712 ( .A1(n352), .A2(n637), .ZN(n636) );
  XNOR2_X1 U713 ( .A(G104), .B(n636), .ZN(G6) );
  NAND2_X1 U714 ( .A1(n637), .A2(n651), .ZN(n643) );
  XOR2_X1 U715 ( .A(KEYINPUT114), .B(KEYINPUT27), .Z(n639) );
  XNOR2_X1 U716 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n638) );
  XNOR2_X1 U717 ( .A(n639), .B(n638), .ZN(n641) );
  XOR2_X1 U718 ( .A(G107), .B(KEYINPUT26), .Z(n640) );
  XNOR2_X1 U719 ( .A(n641), .B(n640), .ZN(n642) );
  XNOR2_X1 U720 ( .A(n643), .B(n642), .ZN(G9) );
  XNOR2_X1 U721 ( .A(G110), .B(n644), .ZN(G12) );
  XOR2_X1 U722 ( .A(G128), .B(KEYINPUT29), .Z(n646) );
  NAND2_X1 U723 ( .A1(n647), .A2(n651), .ZN(n645) );
  XNOR2_X1 U724 ( .A(n646), .B(n645), .ZN(G30) );
  XOR2_X1 U725 ( .A(G146), .B(KEYINPUT115), .Z(n649) );
  NAND2_X1 U726 ( .A1(n647), .A2(n352), .ZN(n648) );
  XNOR2_X1 U727 ( .A(n649), .B(n648), .ZN(G48) );
  NAND2_X1 U728 ( .A1(n652), .A2(n352), .ZN(n650) );
  XNOR2_X1 U729 ( .A(n650), .B(G113), .ZN(G15) );
  NAND2_X1 U730 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U731 ( .A(n653), .B(G116), .ZN(G18) );
  XNOR2_X1 U732 ( .A(G125), .B(n654), .ZN(n655) );
  XNOR2_X1 U733 ( .A(n655), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U734 ( .A(G134), .B(n656), .ZN(G36) );
  XOR2_X1 U735 ( .A(G140), .B(n657), .Z(G42) );
  NOR2_X1 U736 ( .A1(KEYINPUT2), .A2(n729), .ZN(n658) );
  NOR2_X1 U737 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U738 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U739 ( .A(n663), .B(KEYINPUT118), .ZN(n664) );
  NOR2_X1 U740 ( .A1(n665), .A2(n664), .ZN(n669) );
  NOR2_X1 U741 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U742 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U743 ( .A1(n687), .A2(n670), .ZN(n682) );
  NOR2_X1 U744 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U745 ( .A(KEYINPUT50), .B(n676), .ZN(n677) );
  NOR2_X1 U746 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U747 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U748 ( .A(n683), .B(KEYINPUT52), .ZN(n684) );
  INV_X1 U749 ( .A(KEYINPUT120), .ZN(n688) );
  XNOR2_X1 U750 ( .A(n689), .B(n688), .ZN(n690) );
  XNOR2_X1 U751 ( .A(KEYINPUT53), .B(n691), .ZN(G75) );
  NAND2_X1 U752 ( .A1(n710), .A2(G210), .ZN(n694) );
  XOR2_X1 U753 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n693) );
  XNOR2_X1 U754 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n697) );
  XNOR2_X1 U755 ( .A(n695), .B(KEYINPUT57), .ZN(n696) );
  XNOR2_X1 U756 ( .A(n697), .B(n696), .ZN(n699) );
  NAND2_X1 U757 ( .A1(n706), .A2(G469), .ZN(n698) );
  XNOR2_X1 U758 ( .A(n699), .B(n698), .ZN(n700) );
  NOR2_X1 U759 ( .A1(n713), .A2(n700), .ZN(G54) );
  NAND2_X1 U760 ( .A1(n710), .A2(G475), .ZN(n704) );
  XOR2_X1 U761 ( .A(KEYINPUT59), .B(KEYINPUT122), .Z(n701) );
  NAND2_X1 U762 ( .A1(G478), .A2(n706), .ZN(n707) );
  XNOR2_X1 U763 ( .A(n708), .B(n707), .ZN(n709) );
  NOR2_X1 U764 ( .A1(n713), .A2(n709), .ZN(G63) );
  XOR2_X1 U765 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n711) );
  NAND2_X1 U766 ( .A1(n730), .A2(n714), .ZN(n718) );
  NAND2_X1 U767 ( .A1(G953), .A2(G224), .ZN(n715) );
  XNOR2_X1 U768 ( .A(KEYINPUT61), .B(n715), .ZN(n716) );
  NAND2_X1 U769 ( .A1(n716), .A2(G898), .ZN(n717) );
  NAND2_X1 U770 ( .A1(n718), .A2(n717), .ZN(n725) );
  XNOR2_X1 U771 ( .A(G101), .B(n719), .ZN(n721) );
  XNOR2_X1 U772 ( .A(n721), .B(n720), .ZN(n722) );
  NOR2_X1 U773 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U774 ( .A(n725), .B(n724), .ZN(G69) );
  XNOR2_X1 U775 ( .A(n726), .B(n550), .ZN(n728) );
  XOR2_X1 U776 ( .A(n727), .B(n728), .Z(n733) );
  XOR2_X1 U777 ( .A(n733), .B(n729), .Z(n731) );
  NAND2_X1 U778 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U779 ( .A(n732), .B(KEYINPUT126), .ZN(n737) );
  XNOR2_X1 U780 ( .A(G227), .B(n733), .ZN(n734) );
  NAND2_X1 U781 ( .A1(n734), .A2(G900), .ZN(n735) );
  NAND2_X1 U782 ( .A1(n735), .A2(G953), .ZN(n736) );
  NAND2_X1 U783 ( .A1(n737), .A2(n736), .ZN(G72) );
  XNOR2_X1 U784 ( .A(G122), .B(n738), .ZN(G24) );
  XNOR2_X1 U785 ( .A(n739), .B(G119), .ZN(G21) );
  XOR2_X1 U786 ( .A(n740), .B(G131), .Z(G33) );
  XNOR2_X1 U787 ( .A(G143), .B(n741), .ZN(G45) );
  XNOR2_X1 U788 ( .A(G137), .B(KEYINPUT127), .ZN(n743) );
  XNOR2_X1 U789 ( .A(n743), .B(n742), .ZN(G39) );
endmodule

