//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 1 1 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 0 0 1 1 1 1 0 0 0 0 1 0 1 0 0 1 0 1 0 1 0 0 1 0 1 1 1 1 1 1 1 0 1 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n575, new_n577, new_n578, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n587, new_n588, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n628, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT64), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT65), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT66), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n468));
  AND3_X1   g043(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n468), .B1(new_n465), .B2(new_n467), .ZN(new_n470));
  OAI21_X1  g045(.A(G125), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n463), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n465), .A2(new_n467), .ZN(new_n474));
  XNOR2_X1  g049(.A(KEYINPUT66), .B(G2105), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G137), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n464), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G101), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n473), .A2(new_n480), .ZN(G160));
  NOR2_X1   g056(.A1(new_n474), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT68), .ZN(new_n484));
  OAI221_X1 g059(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n463), .C2(G112), .ZN(new_n485));
  INV_X1    g060(.A(G124), .ZN(new_n486));
  XNOR2_X1  g061(.A(KEYINPUT3), .B(G2104), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(new_n475), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n485), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  OR2_X1    g064(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  NAND3_X1  g066(.A1(new_n463), .A2(new_n487), .A3(G138), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G138), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n495), .B1(new_n460), .B2(new_n462), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n496), .B1(new_n469), .B2(new_n470), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n459), .A2(G114), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AND2_X1   g076(.A1(G126), .A2(G2105), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n465), .A2(new_n467), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT69), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT69), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n487), .A2(new_n505), .A3(new_n502), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n501), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n498), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT72), .A2(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G62), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  XOR2_X1   g093(.A(new_n518), .B(KEYINPUT74), .Z(new_n519));
  AOI21_X1  g094(.A(new_n510), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT70), .A2(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT6), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT6), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n524), .A2(KEYINPUT70), .A3(G651), .ZN(new_n525));
  AND4_X1   g100(.A1(new_n512), .A2(new_n523), .A3(new_n514), .A4(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G88), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n523), .A2(new_n525), .A3(G50), .A4(G543), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n528), .A2(KEYINPUT71), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n528), .A2(KEYINPUT71), .ZN(new_n530));
  OAI211_X1 g105(.A(new_n527), .B(KEYINPUT73), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n528), .B(KEYINPUT71), .ZN(new_n533));
  AOI21_X1  g108(.A(KEYINPUT73), .B1(new_n533), .B2(new_n527), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n521), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(KEYINPUT75), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n527), .B1(new_n529), .B2(new_n530), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT73), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(new_n531), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n540), .A2(new_n541), .A3(new_n521), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n536), .A2(new_n542), .ZN(G166));
  NAND3_X1  g118(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT7), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n544), .B(new_n545), .ZN(new_n546));
  AND2_X1   g121(.A1(G63), .A2(G651), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n546), .B1(new_n516), .B2(new_n547), .ZN(new_n548));
  XOR2_X1   g123(.A(KEYINPUT76), .B(G51), .Z(new_n549));
  NAND2_X1  g124(.A1(new_n523), .A2(new_n525), .ZN(new_n550));
  OR3_X1    g125(.A1(new_n549), .A2(new_n550), .A3(new_n513), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n526), .A2(G89), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n548), .A2(new_n551), .A3(new_n552), .ZN(G286));
  INV_X1    g128(.A(G286), .ZN(G168));
  AND2_X1   g129(.A1(new_n523), .A2(new_n525), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  XOR2_X1   g132(.A(KEYINPUT77), .B(G52), .Z(new_n558));
  AOI22_X1  g133(.A1(new_n557), .A2(new_n558), .B1(G90), .B2(new_n526), .ZN(new_n559));
  NAND2_X1  g134(.A1(G77), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G64), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n515), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G651), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n559), .A2(new_n563), .ZN(G301));
  INV_X1    g139(.A(G301), .ZN(G171));
  NAND2_X1  g140(.A1(new_n516), .A2(new_n555), .ZN(new_n566));
  INV_X1    g141(.A(G81), .ZN(new_n567));
  INV_X1    g142(.A(G43), .ZN(new_n568));
  OAI22_X1  g143(.A1(new_n566), .A2(new_n567), .B1(new_n556), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n516), .A2(G56), .ZN(new_n570));
  NAND2_X1  g145(.A1(G68), .A2(G543), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n510), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G860), .ZN(G153));
  AND3_X1   g149(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G36), .ZN(G176));
  NAND2_X1  g151(.A1(G1), .A2(G3), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT8), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n575), .A2(new_n578), .ZN(G188));
  NAND2_X1  g154(.A1(G78), .A2(G543), .ZN(new_n580));
  XOR2_X1   g155(.A(KEYINPUT78), .B(G65), .Z(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n581), .B2(new_n515), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(G651), .B1(new_n526), .B2(G91), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n523), .A2(new_n525), .A3(G53), .A4(G543), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT9), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n583), .A2(new_n585), .ZN(G299));
  AOI21_X1  g161(.A(new_n541), .B1(new_n540), .B2(new_n521), .ZN(new_n587));
  AOI211_X1 g162(.A(KEYINPUT75), .B(new_n520), .C1(new_n539), .C2(new_n531), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n587), .A2(new_n588), .ZN(G303));
  OAI21_X1  g164(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n526), .A2(G87), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n555), .A2(G49), .A3(G543), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(G288));
  NAND4_X1  g168(.A1(new_n555), .A2(KEYINPUT80), .A3(G48), .A4(G543), .ZN(new_n594));
  NAND4_X1  g169(.A1(new_n523), .A2(new_n525), .A3(G48), .A4(G543), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT80), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n594), .A2(new_n597), .B1(G86), .B2(new_n526), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n512), .A2(new_n514), .A3(G61), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT79), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g176(.A1(new_n512), .A2(new_n514), .A3(KEYINPUT79), .A4(G61), .ZN(new_n602));
  NAND2_X1  g177(.A1(G73), .A2(G543), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G651), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n598), .A2(new_n605), .ZN(G305));
  NAND2_X1  g181(.A1(G72), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G60), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n515), .B2(new_n608), .ZN(new_n609));
  AND2_X1   g184(.A1(new_n609), .A2(KEYINPUT81), .ZN(new_n610));
  OAI21_X1  g185(.A(G651), .B1(new_n609), .B2(KEYINPUT81), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n557), .A2(G47), .B1(G85), .B2(new_n526), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(G290));
  NAND2_X1  g189(.A1(G301), .A2(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n526), .A2(G92), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT10), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(G79), .A2(G543), .ZN(new_n619));
  INV_X1    g194(.A(G66), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n515), .B2(new_n620), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n557), .A2(G54), .B1(new_n621), .B2(G651), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n615), .B1(new_n624), .B2(G868), .ZN(G284));
  OAI21_X1  g200(.A(new_n615), .B1(new_n624), .B2(G868), .ZN(G321));
  NAND2_X1  g201(.A1(G286), .A2(G868), .ZN(new_n627));
  INV_X1    g202(.A(G299), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(G868), .ZN(G297));
  OAI21_X1  g204(.A(new_n627), .B1(new_n628), .B2(G868), .ZN(G280));
  INV_X1    g205(.A(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n624), .B1(new_n631), .B2(G860), .ZN(G148));
  INV_X1    g207(.A(new_n573), .ZN(new_n633));
  INV_X1    g208(.A(G868), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n623), .A2(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n636), .B2(new_n634), .ZN(G323));
  XNOR2_X1  g212(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g213(.A1(new_n466), .A2(G2104), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n640));
  OAI21_X1  g215(.A(KEYINPUT67), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(new_n478), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n644), .B(new_n645), .Z(new_n646));
  XOR2_X1   g221(.A(KEYINPUT13), .B(G2100), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n463), .A2(G111), .ZN(new_n650));
  INV_X1    g225(.A(KEYINPUT83), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n652), .B1(new_n651), .B2(new_n650), .ZN(new_n653));
  INV_X1    g228(.A(new_n488), .ZN(new_n654));
  AOI22_X1  g229(.A1(new_n654), .A2(G123), .B1(new_n482), .B2(G135), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(G2096), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n648), .A2(new_n658), .ZN(G156));
  INV_X1    g234(.A(KEYINPUT14), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT15), .B(G2435), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT84), .B(G2438), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2427), .B(G2430), .Z(new_n664));
  AOI21_X1  g239(.A(new_n660), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n665), .B1(new_n664), .B2(new_n663), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2451), .B(G2454), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT16), .B(G1341), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2443), .B(G2446), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G1348), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n669), .B(new_n671), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n666), .A2(new_n672), .ZN(new_n674));
  AND3_X1   g249(.A1(new_n673), .A2(G14), .A3(new_n674), .ZN(G401));
  XOR2_X1   g250(.A(G2084), .B(G2090), .Z(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2067), .B(G2678), .Z(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n678), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n680), .A2(new_n681), .A3(KEYINPUT17), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT85), .B(KEYINPUT18), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(G2100), .Z(new_n685));
  XNOR2_X1  g260(.A(G2072), .B(G2078), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(new_n679), .B2(new_n683), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(new_n657), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n685), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(G227));
  XNOR2_X1  g265(.A(G1971), .B(G1976), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT19), .ZN(new_n692));
  XOR2_X1   g267(.A(G1956), .B(G2474), .Z(new_n693));
  XOR2_X1   g268(.A(G1961), .B(G1966), .Z(new_n694));
  OR2_X1    g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n693), .A2(new_n694), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n692), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n692), .A2(new_n696), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT20), .ZN(new_n699));
  OAI221_X1 g274(.A(new_n697), .B1(new_n692), .B2(new_n695), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(new_n699), .B2(new_n698), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT86), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT87), .B(KEYINPUT88), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n705));
  XNOR2_X1  g280(.A(G1981), .B(G1986), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(G1991), .B(G1996), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n704), .B(new_n709), .ZN(G229));
  INV_X1    g285(.A(G2090), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G35), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G162), .B2(new_n712), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n714), .A2(KEYINPUT29), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(KEYINPUT29), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n711), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G16), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G20), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT104), .Z(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT23), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G299), .B2(G16), .ZN(new_n722));
  INV_X1    g297(.A(G1956), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n717), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT25), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n482), .A2(G139), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT95), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n643), .A2(G127), .ZN(new_n732));
  INV_X1    g307(.A(G115), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(new_n733), .B2(new_n464), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(KEYINPUT96), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT96), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n732), .B(new_n736), .C1(new_n733), .C2(new_n464), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n735), .A2(new_n475), .A3(new_n737), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n731), .A2(G29), .A3(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G2072), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(KEYINPUT98), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n739), .B(new_n741), .C1(G29), .C2(G33), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n740), .A2(KEYINPUT98), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n742), .A2(new_n743), .ZN(new_n745));
  OAI22_X1  g320(.A1(new_n725), .A2(KEYINPUT105), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n715), .A2(new_n711), .A3(new_n716), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n747), .A2(KEYINPUT103), .ZN(new_n748));
  INV_X1    g323(.A(G34), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n749), .A2(KEYINPUT24), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n749), .A2(KEYINPUT24), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n712), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G160), .B2(new_n712), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT97), .ZN(new_n754));
  INV_X1    g329(.A(G2084), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n747), .A2(KEYINPUT103), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n748), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n718), .A2(G19), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n573), .B2(new_n718), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(G1341), .Z(new_n761));
  XOR2_X1   g336(.A(KEYINPUT27), .B(G1996), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n712), .A2(G32), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n654), .A2(G129), .ZN(new_n764));
  NAND3_X1  g339(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT26), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n767), .A2(new_n768), .B1(G105), .B2(new_n478), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n482), .A2(G141), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n764), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT99), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n763), .B1(new_n773), .B2(new_n712), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n761), .B1(new_n762), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n762), .B2(new_n774), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n718), .A2(G4), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n624), .B2(new_n718), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G1348), .ZN(new_n779));
  NOR2_X1   g354(.A1(G5), .A2(G16), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G171), .B2(G16), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n781), .A2(G1961), .ZN(new_n782));
  NOR2_X1   g357(.A1(G27), .A2(G29), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G164), .B2(G29), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G2078), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n779), .A2(new_n782), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(G168), .A2(G16), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G16), .B2(G21), .ZN(new_n788));
  INV_X1    g363(.A(G1966), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT100), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n653), .A2(G29), .A3(new_n655), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n792), .A2(KEYINPUT101), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT30), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n794), .A2(G28), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n712), .B1(new_n794), .B2(G28), .ZN(new_n796));
  AND2_X1   g371(.A1(KEYINPUT31), .A2(G11), .ZN(new_n797));
  NOR2_X1   g372(.A1(KEYINPUT31), .A2(G11), .ZN(new_n798));
  OAI22_X1  g373(.A1(new_n795), .A2(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(new_n792), .B2(KEYINPUT101), .ZN(new_n800));
  AOI22_X1  g375(.A1(G1961), .A2(new_n781), .B1(new_n788), .B2(new_n789), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n791), .A2(new_n793), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n776), .B(new_n786), .C1(new_n802), .C2(KEYINPUT102), .ZN(new_n803));
  NOR3_X1   g378(.A1(new_n746), .A2(new_n758), .A3(new_n803), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n654), .A2(G128), .B1(new_n482), .B2(G140), .ZN(new_n805));
  OAI221_X1 g380(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n463), .C2(G116), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT93), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(G29), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT94), .Z(new_n811));
  NAND2_X1  g386(.A1(new_n712), .A2(G26), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT28), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(G2067), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n802), .A2(KEYINPUT102), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n725), .A2(KEYINPUT105), .ZN(new_n818));
  AND3_X1   g393(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n804), .A2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT36), .ZN(new_n821));
  MUX2_X1   g396(.A(G6), .B(G305), .S(G16), .Z(new_n822));
  OR2_X1    g397(.A1(new_n822), .A2(KEYINPUT91), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(KEYINPUT91), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT32), .B(G1981), .Z(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n823), .A2(new_n824), .A3(new_n826), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n718), .A2(G23), .ZN(new_n830));
  INV_X1    g405(.A(G288), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n831), .B2(new_n718), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT33), .B(G1976), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT92), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n832), .B(new_n834), .ZN(new_n835));
  AND3_X1   g410(.A1(new_n828), .A2(new_n829), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(G16), .A2(G22), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(G166), .B2(G16), .ZN(new_n838));
  INV_X1    g413(.A(G1971), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n841), .A2(KEYINPUT34), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(G25), .A2(G29), .ZN(new_n844));
  AOI22_X1  g419(.A1(new_n654), .A2(G119), .B1(new_n482), .B2(G131), .ZN(new_n845));
  OAI221_X1 g420(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n463), .C2(G107), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT89), .Z(new_n848));
  AOI21_X1  g423(.A(new_n844), .B1(new_n848), .B2(G29), .ZN(new_n849));
  XNOR2_X1  g424(.A(KEYINPUT35), .B(G1991), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n849), .B(new_n850), .Z(new_n851));
  INV_X1    g426(.A(G290), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n852), .A2(new_n718), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(new_n718), .B2(G24), .ZN(new_n854));
  XOR2_X1   g429(.A(KEYINPUT90), .B(G1986), .Z(new_n855));
  OR2_X1    g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n855), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n851), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n858), .B1(new_n841), .B2(KEYINPUT34), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n821), .B1(new_n843), .B2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n843), .A2(new_n821), .A3(new_n859), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n820), .B1(new_n861), .B2(new_n862), .ZN(G311));
  INV_X1    g438(.A(new_n862), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n819), .B(new_n804), .C1(new_n864), .C2(new_n860), .ZN(G150));
  NOR2_X1   g440(.A1(new_n623), .A2(new_n631), .ZN(new_n866));
  XNOR2_X1  g441(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(G93), .ZN(new_n869));
  INV_X1    g444(.A(G55), .ZN(new_n870));
  OAI22_X1  g445(.A1(new_n566), .A2(new_n869), .B1(new_n556), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n516), .A2(G67), .ZN(new_n872));
  NAND2_X1  g447(.A1(G80), .A2(G543), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n510), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(new_n573), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n871), .A2(new_n874), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(new_n572), .B2(new_n569), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(G860), .B1(new_n868), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n881), .B1(new_n880), .B2(new_n868), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n875), .A2(G860), .ZN(new_n883));
  XOR2_X1   g458(.A(KEYINPUT106), .B(KEYINPUT37), .Z(new_n884));
  XNOR2_X1  g459(.A(new_n883), .B(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n882), .A2(new_n885), .ZN(G145));
  XNOR2_X1  g461(.A(new_n490), .B(G164), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n656), .B(G160), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n887), .B(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n731), .A2(new_n773), .A3(new_n738), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n771), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n893), .B1(new_n731), .B2(new_n738), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n646), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n894), .ZN(new_n896));
  INV_X1    g471(.A(new_n646), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n896), .A2(new_n897), .A3(new_n891), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n654), .A2(G130), .ZN(new_n899));
  OAI221_X1 g474(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n463), .C2(G118), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n482), .A2(G142), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n895), .A2(new_n898), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n902), .B1(new_n895), .B2(new_n898), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n890), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n895), .A2(new_n898), .ZN(new_n907));
  INV_X1    g482(.A(new_n902), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n909), .A2(new_n889), .A3(new_n903), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n809), .B(new_n847), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n906), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(G37), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n911), .B1(new_n906), .B2(new_n910), .ZN(new_n915));
  OR3_X1    g490(.A1(new_n914), .A2(KEYINPUT40), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(KEYINPUT40), .B1(new_n914), .B2(new_n915), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(G395));
  INV_X1    g493(.A(KEYINPUT107), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT42), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n831), .B1(new_n587), .B2(new_n588), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n536), .A2(new_n542), .A3(G288), .ZN(new_n922));
  XNOR2_X1  g497(.A(G290), .B(G305), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n923), .B1(new_n921), .B2(new_n922), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n920), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n923), .ZN(new_n927));
  NOR3_X1   g502(.A1(new_n587), .A2(new_n588), .A3(new_n831), .ZN(new_n928));
  AOI21_X1  g503(.A(G288), .B1(new_n536), .B2(new_n542), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n931));
  XNOR2_X1  g506(.A(KEYINPUT107), .B(KEYINPUT42), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n926), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n880), .A2(new_n636), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n879), .B1(G559), .B2(new_n623), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n623), .A2(new_n628), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n618), .A2(G299), .A3(new_n622), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n937), .A2(new_n938), .A3(new_n941), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n939), .A2(KEYINPUT41), .A3(new_n940), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT41), .B1(new_n939), .B2(new_n940), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n937), .A2(new_n938), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n942), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n935), .A2(new_n936), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n945), .B1(new_n937), .B2(new_n938), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n926), .B(new_n934), .C1(new_n950), .C2(new_n942), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n936), .B1(new_n935), .B2(new_n948), .ZN(new_n953));
  OAI21_X1  g528(.A(G868), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n875), .A2(new_n634), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(G331));
  NAND2_X1  g531(.A1(G331), .A2(KEYINPUT109), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT109), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n954), .A2(new_n958), .A3(new_n955), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n959), .ZN(G295));
  NAND2_X1  g535(.A1(G301), .A2(G168), .ZN(new_n961));
  NAND3_X1  g536(.A1(G286), .A2(new_n559), .A3(new_n563), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AOI22_X1  g538(.A1(new_n879), .A2(new_n963), .B1(new_n939), .B2(new_n940), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n876), .A2(new_n878), .A3(new_n961), .A4(new_n962), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT110), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n965), .A2(new_n966), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n964), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n879), .A2(new_n963), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n965), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n971), .B1(new_n943), .B2(new_n944), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n969), .A2(new_n972), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n973), .A2(new_n924), .A3(new_n925), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n973), .B1(new_n924), .B2(new_n925), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n913), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n974), .B1(new_n976), .B2(KEYINPUT111), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT111), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n975), .A2(new_n978), .A3(new_n913), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT43), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n974), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n964), .A2(new_n965), .ZN(new_n982));
  INV_X1    g557(.A(new_n968), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n965), .A2(new_n966), .ZN(new_n984));
  AOI22_X1  g559(.A1(new_n983), .A2(new_n984), .B1(new_n879), .B2(new_n963), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n982), .B1(new_n985), .B2(new_n945), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n986), .B1(new_n924), .B2(new_n925), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n981), .A2(new_n987), .A3(new_n913), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT43), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT44), .B1(new_n980), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT44), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n989), .B1(new_n977), .B2(new_n979), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n988), .A2(KEYINPUT43), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n991), .A2(new_n995), .ZN(G397));
  INV_X1    g571(.A(G1384), .ZN(new_n997));
  AOI22_X1  g572(.A1(new_n643), .A2(new_n496), .B1(new_n492), .B2(KEYINPUT4), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n505), .B1(new_n487), .B2(new_n502), .ZN(new_n999));
  AND4_X1   g574(.A1(new_n505), .A2(new_n465), .A3(new_n467), .A4(new_n502), .ZN(new_n1000));
  OAI22_X1  g575(.A1(new_n999), .A2(new_n1000), .B1(new_n499), .B2(new_n500), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n997), .B1(new_n998), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI22_X1  g579(.A1(new_n476), .A2(G137), .B1(G101), .B2(new_n478), .ZN(new_n1005));
  XOR2_X1   g580(.A(KEYINPUT112), .B(G40), .Z(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  AOI22_X1  g582(.A1(new_n643), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1005), .B(new_n1007), .C1(new_n1008), .C2(new_n463), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1004), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n809), .B(G2067), .ZN(new_n1011));
  INV_X1    g586(.A(G1996), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n893), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1010), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  NOR3_X1   g589(.A1(new_n1004), .A2(G1996), .A3(new_n1009), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1015), .A2(KEYINPUT114), .A3(new_n773), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1015), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1017), .B1(new_n1018), .B2(new_n772), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n1014), .A2(new_n1016), .A3(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n847), .B(new_n850), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1010), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G1986), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n852), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n852), .A2(new_n1024), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1010), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  XOR2_X1   g603(.A(new_n1028), .B(KEYINPUT113), .Z(new_n1029));
  NOR2_X1   g604(.A1(new_n1023), .A2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n1030), .B(KEYINPUT115), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n590), .A2(new_n591), .A3(G1976), .A4(new_n592), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n1032), .B(KEYINPUT116), .ZN(new_n1033));
  NAND4_X1  g608(.A1(G160), .A2(new_n997), .A3(new_n508), .A4(new_n1007), .ZN(new_n1034));
  XOR2_X1   g609(.A(KEYINPUT117), .B(G1976), .Z(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT52), .B1(G288), .B2(new_n1035), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1033), .A2(new_n1034), .A3(G8), .A4(new_n1036), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1033), .A2(new_n1034), .A3(G8), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT52), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1037), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G1981), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n598), .A2(new_n605), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n598), .A2(new_n605), .A3(KEYINPUT118), .A4(new_n1041), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT119), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n605), .B1(new_n598), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n594), .A2(new_n597), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n526), .A2(G86), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(new_n1047), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(G1981), .B1(new_n1048), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1046), .A2(new_n1053), .A3(KEYINPUT49), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT120), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1046), .A2(new_n1053), .A3(KEYINPUT120), .A4(KEYINPUT49), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT49), .B1(new_n1046), .B2(new_n1053), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1009), .A2(new_n1002), .ZN(new_n1060));
  INV_X1    g635(.A(G8), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1059), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1040), .B1(new_n1058), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1002), .A2(KEYINPUT50), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n473), .A2(new_n480), .A3(new_n1006), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT50), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n508), .A2(new_n1068), .A3(new_n997), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1066), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n711), .ZN(new_n1071));
  OAI211_X1 g646(.A(KEYINPUT45), .B(new_n997), .C1(new_n998), .C2(new_n1001), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1004), .A2(new_n1067), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n839), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1061), .B1(new_n1071), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n536), .A2(G8), .A3(new_n542), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT55), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1075), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n1070), .A2(new_n711), .B1(new_n1073), .B2(new_n839), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1081), .B(new_n1082), .C1(new_n1061), .C2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n1085));
  INV_X1    g660(.A(G2078), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1004), .A2(new_n1086), .A3(new_n1067), .A4(new_n1072), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1066), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1088));
  INV_X1    g663(.A(G1961), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1085), .A2(new_n1087), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT45), .B1(new_n508), .B2(new_n997), .ZN(new_n1091));
  AOI211_X1 g666(.A(new_n1003), .B(G1384), .C1(new_n498), .C2(new_n507), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1093), .A2(KEYINPUT53), .A3(new_n1086), .A4(new_n1067), .ZN(new_n1094));
  AOI21_X1  g669(.A(G301), .B1(new_n1090), .B2(new_n1094), .ZN(new_n1095));
  AND4_X1   g670(.A1(new_n1065), .A2(new_n1080), .A3(new_n1084), .A4(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1073), .A2(new_n789), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1066), .A2(new_n1069), .A3(new_n755), .A4(new_n1067), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1061), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT51), .B1(new_n1099), .B2(KEYINPUT124), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1070), .A2(new_n755), .B1(new_n1073), .B2(new_n789), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1061), .B1(new_n1101), .B2(G168), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1099), .ZN(new_n1104));
  NAND2_X1  g679(.A1(G286), .A2(G8), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1104), .A2(KEYINPUT124), .A3(KEYINPUT51), .A4(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT62), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1103), .A2(new_n1106), .A3(new_n1107), .A4(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1096), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1108), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1107), .B1(new_n1112), .B2(new_n1106), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT126), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1113), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT126), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1115), .A2(new_n1116), .A3(new_n1110), .A4(new_n1096), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(G299), .A2(KEYINPUT121), .A3(KEYINPUT57), .ZN(new_n1119));
  OR2_X1    g694(.A1(KEYINPUT121), .A2(KEYINPUT57), .ZN(new_n1120));
  NAND2_X1  g695(.A1(KEYINPUT121), .A2(KEYINPUT57), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n583), .A2(new_n585), .A3(new_n1120), .A4(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1009), .B1(KEYINPUT50), .B2(new_n1002), .ZN(new_n1124));
  AOI21_X1  g699(.A(G1956), .B1(new_n1124), .B2(new_n1069), .ZN(new_n1125));
  XNOR2_X1  g700(.A(KEYINPUT56), .B(G2072), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1004), .A2(new_n1067), .A3(new_n1072), .A4(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1123), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(G1348), .B1(new_n1124), .B2(new_n1069), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1060), .A2(new_n815), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1129), .B1(new_n1133), .B2(new_n623), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1088), .A2(new_n723), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1123), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1135), .A2(new_n1136), .A3(new_n1127), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1135), .A2(new_n1136), .A3(new_n1127), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1136), .B1(new_n1135), .B2(new_n1127), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1139), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT60), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1143), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1144));
  OAI211_X1 g719(.A(KEYINPUT60), .B(new_n1131), .C1(new_n1070), .C2(G1348), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1144), .A2(new_n624), .A3(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1129), .A2(KEYINPUT61), .A3(new_n1137), .ZN(new_n1147));
  XOR2_X1   g722(.A(KEYINPUT58), .B(G1341), .Z(new_n1148));
  NAND2_X1  g723(.A1(new_n1034), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1034), .A2(KEYINPUT122), .A3(new_n1148), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1004), .A2(new_n1012), .A3(new_n1067), .A4(new_n1072), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(KEYINPUT123), .A2(KEYINPUT59), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n633), .B1(KEYINPUT123), .B2(KEYINPUT59), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1154), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1142), .A2(new_n1146), .A3(new_n1147), .A4(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1133), .A2(KEYINPUT60), .A3(new_n623), .ZN(new_n1160));
  AND2_X1   g735(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1160), .B1(new_n1161), .B2(new_n1156), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1138), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT54), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1087), .A2(new_n1085), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1166));
  AND3_X1   g741(.A1(new_n1086), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1004), .A2(G160), .A3(new_n1072), .A4(new_n1167), .ZN(new_n1168));
  AND4_X1   g743(.A1(G301), .A2(new_n1165), .A3(new_n1166), .A4(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1164), .B1(new_n1095), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT125), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  OAI211_X1 g747(.A(KEYINPUT125), .B(new_n1164), .C1(new_n1095), .C2(new_n1169), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  AND3_X1   g749(.A1(new_n1065), .A2(new_n1080), .A3(new_n1084), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1094), .A2(new_n1165), .A3(G301), .A4(new_n1166), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(KEYINPUT54), .ZN(new_n1177));
  AOI21_X1  g752(.A(G301), .B1(new_n1090), .B2(new_n1168), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1179), .B1(new_n1112), .B2(new_n1106), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1163), .A2(new_n1174), .A3(new_n1175), .A4(new_n1180), .ZN(new_n1181));
  AND2_X1   g756(.A1(new_n1080), .A2(new_n1084), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1104), .A2(G286), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1182), .A2(KEYINPUT63), .A3(new_n1065), .A4(new_n1183), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1065), .A2(new_n1080), .A3(new_n1183), .A4(new_n1084), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT63), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1184), .A2(new_n1187), .ZN(new_n1188));
  AND2_X1   g763(.A1(new_n1058), .A2(new_n1064), .ZN(new_n1189));
  NOR3_X1   g764(.A1(new_n1189), .A2(new_n1080), .A3(new_n1040), .ZN(new_n1190));
  OR2_X1    g765(.A1(G288), .A2(G1976), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1046), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1190), .B1(new_n1062), .B2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1181), .A2(new_n1188), .A3(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1031), .B1(new_n1118), .B2(new_n1194), .ZN(new_n1195));
  OR2_X1    g770(.A1(new_n1023), .A2(KEYINPUT127), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1023), .A2(KEYINPUT127), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1026), .A2(new_n1010), .ZN(new_n1198));
  XNOR2_X1  g773(.A(new_n1198), .B(KEYINPUT48), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1196), .A2(new_n1197), .A3(new_n1199), .ZN(new_n1200));
  INV_X1    g775(.A(new_n848), .ZN(new_n1201));
  NOR2_X1   g776(.A1(new_n1201), .A2(new_n850), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1020), .A2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1203), .B1(G2067), .B2(new_n809), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1204), .A2(new_n1010), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1010), .B1(new_n1011), .B2(new_n771), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1015), .A2(KEYINPUT46), .ZN(new_n1207));
  OR2_X1    g782(.A1(new_n1015), .A2(KEYINPUT46), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  XNOR2_X1  g784(.A(new_n1209), .B(KEYINPUT47), .ZN(new_n1210));
  AND3_X1   g785(.A1(new_n1200), .A2(new_n1205), .A3(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1195), .A2(new_n1211), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g787(.A(G401), .ZN(new_n1214));
  NAND3_X1  g788(.A1(new_n689), .A2(G319), .A3(new_n1214), .ZN(new_n1215));
  NOR2_X1   g789(.A1(G229), .A2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g790(.A(new_n1216), .B1(new_n914), .B2(new_n915), .ZN(new_n1217));
  NOR2_X1   g791(.A1(new_n993), .A2(new_n994), .ZN(new_n1218));
  NOR2_X1   g792(.A1(new_n1217), .A2(new_n1218), .ZN(G308));
  OAI221_X1 g793(.A(new_n1216), .B1(new_n914), .B2(new_n915), .C1(new_n993), .C2(new_n994), .ZN(G225));
endmodule


