//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 1 1 0 1 1 0 0 1 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 1 1 0 0 1 0 1 0 1 0 0 0 1 0 0 0 0 0 0 1 0 1 0 0 1 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n447, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n566, new_n567, new_n569, new_n570, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n612, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n840, new_n841, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1166,
    new_n1167, new_n1168, new_n1169;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT67), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XOR2_X1   g013(.A(KEYINPUT68), .B(G69), .Z(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  AND2_X1   g017(.A1(G2072), .A2(G2078), .ZN(new_n443));
  NAND3_X1  g018(.A1(new_n443), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  NAND2_X1  g021(.A1(G94), .A2(G452), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT69), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  XOR2_X1   g029(.A(KEYINPUT70), .B(KEYINPUT71), .Z(new_n455));
  XNOR2_X1  g030(.A(new_n454), .B(new_n455), .ZN(new_n456));
  OR4_X1    g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n456), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT73), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n461), .B1(new_n462), .B2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n461), .A2(new_n462), .A3(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT74), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n469), .A2(new_n470), .A3(G137), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  OAI21_X1  g047(.A(KEYINPUT74), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n471), .A2(new_n473), .B1(G101), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n474), .A2(KEYINPUT3), .ZN(new_n478));
  AOI21_X1  g053(.A(KEYINPUT72), .B1(new_n464), .B2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n464), .A2(new_n478), .A3(KEYINPUT72), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n477), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AND2_X1   g057(.A1(G113), .A2(G2104), .ZN(new_n483));
  OAI21_X1  g058(.A(G2105), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n476), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G160));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT75), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n474), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI221_X1 g064(.A(new_n489), .B1(new_n488), .B2(new_n487), .C1(G112), .C2(new_n466), .ZN(new_n490));
  INV_X1    g065(.A(G136), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(new_n468), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n465), .A2(G2105), .A3(new_n467), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n492), .B1(G124), .B2(new_n494), .ZN(G162));
  OR3_X1    g070(.A1(new_n466), .A2(KEYINPUT76), .A3(G114), .ZN(new_n496));
  OR2_X1    g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(KEYINPUT76), .B1(new_n466), .B2(G114), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n496), .A2(G2104), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G126), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n499), .B1(new_n493), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G138), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n502), .A2(G2105), .ZN(new_n503));
  AOI21_X1  g078(.A(KEYINPUT73), .B1(new_n474), .B2(KEYINPUT3), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n474), .A2(KEYINPUT3), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n467), .B(new_n503), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT77), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT77), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n465), .A2(new_n508), .A3(new_n467), .A4(new_n503), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n507), .A2(KEYINPUT4), .A3(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT4), .ZN(new_n511));
  INV_X1    g086(.A(new_n481), .ZN(new_n512));
  OAI211_X1 g087(.A(new_n511), .B(new_n503), .C1(new_n512), .C2(new_n479), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n501), .B1(new_n510), .B2(new_n513), .ZN(G164));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  XOR2_X1   g090(.A(new_n515), .B(KEYINPUT79), .Z(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT5), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT5), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G543), .ZN(new_n520));
  AND3_X1   g095(.A1(new_n518), .A2(new_n520), .A3(G62), .ZN(new_n521));
  OAI21_X1  g096(.A(G651), .B1(new_n516), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT80), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n518), .A2(new_n520), .ZN(new_n524));
  AND2_X1   g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  NOR2_X1   g100(.A1(KEYINPUT6), .A2(G651), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OR3_X1    g102(.A1(new_n524), .A2(new_n527), .A3(KEYINPUT78), .ZN(new_n528));
  OAI21_X1  g103(.A(KEYINPUT78), .B1(new_n524), .B2(new_n527), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G88), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n527), .A2(new_n517), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G50), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n523), .A2(new_n531), .A3(new_n533), .ZN(G303));
  INV_X1    g109(.A(G303), .ZN(G166));
  AND2_X1   g110(.A1(new_n518), .A2(new_n520), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n536), .A2(G63), .A3(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n532), .A2(G51), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n528), .A2(G89), .A3(new_n529), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT7), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n539), .A2(KEYINPUT81), .A3(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(KEYINPUT81), .B1(new_n539), .B2(new_n541), .ZN(new_n544));
  OAI211_X1 g119(.A(new_n537), .B(new_n538), .C1(new_n543), .C2(new_n544), .ZN(G286));
  INV_X1    g120(.A(G286), .ZN(G168));
  NAND2_X1  g121(.A1(G77), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G64), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n524), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G651), .ZN(new_n550));
  INV_X1    g125(.A(G52), .ZN(new_n551));
  INV_X1    g126(.A(new_n532), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n553), .B1(new_n530), .B2(G90), .ZN(G171));
  NAND3_X1  g129(.A1(new_n528), .A2(G81), .A3(new_n529), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n532), .A2(G43), .ZN(new_n556));
  NAND2_X1  g131(.A1(G68), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G56), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n524), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G651), .ZN(new_n560));
  AND2_X1   g135(.A1(new_n560), .A2(KEYINPUT82), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n560), .A2(KEYINPUT82), .ZN(new_n562));
  OAI211_X1 g137(.A(new_n555), .B(new_n556), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  AND3_X1   g140(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G36), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT83), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n566), .A2(new_n570), .ZN(G188));
  NAND2_X1  g146(.A1(new_n530), .A2(G91), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n532), .A2(G53), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT9), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n536), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G651), .ZN(new_n576));
  OR2_X1    g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n572), .A2(new_n574), .A3(new_n577), .ZN(G299));
  INV_X1    g153(.A(G171), .ZN(G301));
  NAND2_X1  g154(.A1(new_n532), .A2(G49), .ZN(new_n580));
  XOR2_X1   g155(.A(new_n580), .B(KEYINPUT84), .Z(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n536), .B2(G74), .ZN(new_n582));
  XOR2_X1   g157(.A(new_n582), .B(KEYINPUT85), .Z(new_n583));
  NAND2_X1  g158(.A1(new_n530), .A2(G87), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n581), .A2(new_n583), .A3(new_n584), .ZN(G288));
  NAND2_X1  g160(.A1(new_n530), .A2(G86), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G61), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n524), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(G651), .B1(new_n532), .B2(G48), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n586), .A2(new_n590), .ZN(G305));
  NAND2_X1  g166(.A1(new_n530), .A2(G85), .ZN(new_n592));
  NAND2_X1  g167(.A1(G72), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G60), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n524), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n595), .A2(G651), .B1(new_n532), .B2(G47), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n592), .A2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n530), .A2(G92), .ZN(new_n599));
  XOR2_X1   g174(.A(new_n599), .B(KEYINPUT10), .Z(new_n600));
  NAND2_X1  g175(.A1(new_n532), .A2(G54), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n536), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n602), .A2(new_n576), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n598), .B1(new_n605), .B2(G868), .ZN(G284));
  OAI21_X1  g181(.A(new_n598), .B1(new_n605), .B2(G868), .ZN(G321));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(G299), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G168), .B2(new_n608), .ZN(G297));
  OAI21_X1  g185(.A(new_n609), .B1(G168), .B2(new_n608), .ZN(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n605), .B1(new_n612), .B2(G860), .ZN(G148));
  NAND2_X1  g188(.A1(new_n605), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G868), .B2(new_n564), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n480), .A2(new_n481), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(new_n475), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n619), .B(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT13), .Z(new_n623));
  NAND2_X1  g198(.A1(KEYINPUT87), .A2(G2100), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n494), .A2(G123), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n469), .A2(G135), .ZN(new_n627));
  NOR2_X1   g202(.A1(G99), .A2(G2105), .ZN(new_n628));
  OAI21_X1  g203(.A(G2104), .B1(new_n466), .B2(G111), .ZN(new_n629));
  OAI211_X1 g204(.A(new_n626), .B(new_n627), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT88), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2096), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n625), .B(new_n632), .C1(KEYINPUT87), .C2(G2100), .ZN(G156));
  XNOR2_X1  g208(.A(G2427), .B(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2430), .ZN(new_n635));
  XOR2_X1   g210(.A(KEYINPUT15), .B(G2435), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(KEYINPUT14), .ZN(new_n638));
  XOR2_X1   g213(.A(G2451), .B(G2454), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT16), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n640), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G1341), .B(G1348), .Z(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n646), .A2(KEYINPUT89), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n643), .A2(new_n645), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(KEYINPUT89), .ZN(new_n649));
  NAND4_X1  g224(.A1(new_n647), .A2(G14), .A3(new_n648), .A4(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(G401));
  NOR2_X1   g226(.A1(G2072), .A2(G2078), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n443), .A2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(KEYINPUT90), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2067), .B(G2678), .Z(new_n656));
  OAI21_X1  g231(.A(KEYINPUT90), .B1(new_n443), .B2(new_n652), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT91), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n653), .B(KEYINPUT17), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n662), .B1(new_n656), .B2(new_n663), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n660), .A2(new_n653), .A3(new_n656), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT18), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n663), .A2(new_n659), .A3(new_n656), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n664), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2100), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT92), .B(G2096), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(G227));
  XNOR2_X1  g247(.A(G1971), .B(G1976), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  XOR2_X1   g249(.A(G1956), .B(G2474), .Z(new_n675));
  XOR2_X1   g250(.A(G1961), .B(G1966), .Z(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n674), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n675), .A2(new_n676), .ZN(new_n680));
  AOI22_X1  g255(.A1(new_n678), .A2(KEYINPUT20), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n680), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n682), .A2(new_n674), .A3(new_n677), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n681), .B(new_n683), .C1(KEYINPUT20), .C2(new_n678), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1986), .B(G1996), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G1981), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G1991), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n686), .B(new_n689), .ZN(G229));
  INV_X1    g265(.A(G16), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n691), .A2(G23), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(G288), .B2(G16), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT94), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI211_X1 g270(.A(KEYINPUT94), .B(new_n692), .C1(G288), .C2(G16), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT33), .B(G1976), .Z(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  OR3_X1    g273(.A1(new_n695), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(G303), .A2(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n691), .A2(G22), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G1971), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n699), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT34), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n691), .A2(G6), .ZN(new_n707));
  INV_X1    g282(.A(G305), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(new_n691), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT32), .B(G1981), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n698), .B1(new_n695), .B2(new_n696), .ZN(new_n712));
  NAND4_X1  g287(.A1(new_n705), .A2(new_n706), .A3(new_n711), .A4(new_n712), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n691), .A2(G24), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(G290), .B2(G16), .ZN(new_n715));
  INV_X1    g290(.A(G1986), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G25), .ZN(new_n719));
  INV_X1    g294(.A(G119), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n493), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT93), .ZN(new_n722));
  OR2_X1    g297(.A1(G95), .A2(G2105), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n723), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n469), .A2(G131), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n722), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n719), .B1(new_n727), .B2(new_n718), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT35), .B(G1991), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n717), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n729), .B2(new_n728), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n699), .A2(new_n704), .A3(new_n711), .A4(new_n712), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(KEYINPUT34), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n715), .A2(new_n716), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n713), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(KEYINPUT95), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT95), .ZN(new_n737));
  NAND4_X1  g312(.A1(new_n713), .A2(new_n733), .A3(new_n737), .A4(new_n734), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT36), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n718), .A2(G35), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G162), .B2(new_n718), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT29), .B(G2090), .Z(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n736), .A2(KEYINPUT36), .A3(new_n738), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n718), .A2(G32), .ZN(new_n747));
  INV_X1    g322(.A(G129), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n493), .A2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT101), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND3_X1  g326(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT26), .Z(new_n753));
  AOI22_X1  g328(.A1(new_n469), .A2(G141), .B1(G105), .B2(new_n475), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n751), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT102), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n755), .A2(new_n756), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n747), .B1(new_n760), .B2(new_n718), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT27), .B(G1996), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n691), .A2(G20), .ZN(new_n764));
  INV_X1    g339(.A(G299), .ZN(new_n765));
  OAI211_X1 g340(.A(KEYINPUT23), .B(new_n764), .C1(new_n765), .C2(new_n691), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(KEYINPUT23), .B2(new_n764), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G1956), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n763), .A2(new_n768), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n691), .A2(G4), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n604), .B2(G16), .ZN(new_n771));
  INV_X1    g346(.A(G1348), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n691), .A2(G5), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G171), .B2(new_n691), .ZN(new_n776));
  AND2_X1   g351(.A1(new_n776), .A2(G1961), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n776), .A2(G1961), .ZN(new_n778));
  INV_X1    g353(.A(G28), .ZN(new_n779));
  NOR3_X1   g354(.A1(new_n779), .A2(KEYINPUT104), .A3(KEYINPUT30), .ZN(new_n780));
  OAI21_X1  g355(.A(KEYINPUT104), .B1(new_n779), .B2(KEYINPUT30), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(new_n718), .ZN(new_n782));
  AOI211_X1 g357(.A(new_n780), .B(new_n782), .C1(KEYINPUT30), .C2(new_n779), .ZN(new_n783));
  NOR3_X1   g358(.A1(new_n777), .A2(new_n778), .A3(new_n783), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT96), .B(KEYINPUT28), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT97), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n718), .A2(G26), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n786), .B(new_n787), .Z(new_n788));
  INV_X1    g363(.A(G140), .ZN(new_n789));
  NOR2_X1   g364(.A1(G104), .A2(G2105), .ZN(new_n790));
  OAI21_X1  g365(.A(G2104), .B1(new_n466), .B2(G116), .ZN(new_n791));
  OAI22_X1  g366(.A1(new_n468), .A2(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G128), .B2(new_n494), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n788), .B1(new_n793), .B2(new_n718), .ZN(new_n794));
  INV_X1    g369(.A(G2067), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT103), .B(KEYINPUT31), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G11), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n631), .A2(G29), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n784), .A2(new_n796), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  AND2_X1   g375(.A1(KEYINPUT24), .A2(G34), .ZN(new_n801));
  NOR2_X1   g376(.A1(KEYINPUT24), .A2(G34), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n801), .A2(new_n802), .A3(G29), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(new_n485), .B2(G29), .ZN(new_n804));
  INV_X1    g379(.A(G2084), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NOR4_X1   g381(.A1(new_n773), .A2(new_n774), .A3(new_n800), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n691), .A2(G19), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(new_n564), .B2(new_n691), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(G1341), .Z(new_n810));
  NAND2_X1  g385(.A1(new_n691), .A2(G21), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G168), .B2(new_n691), .ZN(new_n812));
  INV_X1    g387(.A(G1966), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n769), .A2(new_n807), .A3(new_n810), .A4(new_n814), .ZN(new_n815));
  AOI22_X1  g390(.A1(new_n618), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT98), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(G2105), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n469), .A2(G139), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n475), .A2(G103), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT25), .Z(new_n821));
  NAND3_X1  g396(.A1(new_n818), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(G29), .ZN(new_n824));
  OR2_X1    g399(.A1(G29), .A2(G33), .ZN(new_n825));
  AOI21_X1  g400(.A(G2072), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT99), .Z(new_n827));
  NAND3_X1  g402(.A1(new_n824), .A2(G2072), .A3(new_n825), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT100), .Z(new_n829));
  INV_X1    g404(.A(G27), .ZN(new_n830));
  OAI21_X1  g405(.A(KEYINPUT105), .B1(new_n830), .B2(G29), .ZN(new_n831));
  OR3_X1    g406(.A1(new_n830), .A2(KEYINPUT105), .A3(G29), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n831), .B(new_n832), .C1(G164), .C2(new_n718), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT106), .Z(new_n834));
  OR2_X1    g409(.A1(new_n834), .A2(G2078), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(G2078), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n827), .A2(new_n829), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n815), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n741), .A2(new_n745), .A3(new_n746), .A4(new_n838), .ZN(G150));
  INV_X1    g414(.A(KEYINPUT107), .ZN(new_n840));
  NAND2_X1  g415(.A1(G150), .A2(new_n840), .ZN(new_n841));
  AND2_X1   g416(.A1(new_n746), .A2(new_n838), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n842), .A2(KEYINPUT107), .A3(new_n745), .A4(new_n741), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(G311));
  AOI22_X1  g419(.A1(new_n536), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n845), .A2(new_n576), .ZN(new_n846));
  XOR2_X1   g421(.A(KEYINPUT108), .B(G93), .Z(new_n847));
  NAND3_X1  g422(.A1(new_n528), .A2(new_n529), .A3(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(G55), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n846), .B(new_n848), .C1(new_n849), .C2(new_n552), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(G860), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT37), .Z(new_n852));
  NAND2_X1  g427(.A1(new_n605), .A2(G559), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT38), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n563), .B(new_n850), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(KEYINPUT39), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n854), .B(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n852), .B1(new_n857), .B2(G860), .ZN(G145));
  INV_X1    g433(.A(G162), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n510), .A2(new_n513), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT109), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n510), .A2(KEYINPUT109), .A3(new_n513), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n501), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n793), .B1(new_n758), .B2(new_n759), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n755), .A2(new_n756), .ZN(new_n866));
  INV_X1    g441(.A(new_n793), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n866), .A2(new_n867), .A3(new_n757), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n865), .A2(new_n868), .A3(new_n822), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n822), .B1(new_n865), .B2(new_n868), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n864), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n865), .A2(new_n868), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(new_n823), .ZN(new_n874));
  INV_X1    g449(.A(new_n501), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n510), .A2(KEYINPUT109), .A3(new_n513), .ZN(new_n876));
  AOI21_X1  g451(.A(KEYINPUT109), .B1(new_n510), .B2(new_n513), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n874), .A2(new_n878), .A3(new_n869), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n494), .A2(G130), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n469), .A2(G142), .ZN(new_n881));
  NOR2_X1   g456(.A1(G106), .A2(G2105), .ZN(new_n882));
  OAI21_X1  g457(.A(G2104), .B1(new_n466), .B2(G118), .ZN(new_n883));
  OAI211_X1 g458(.A(new_n880), .B(new_n881), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n622), .B(new_n884), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n885), .A2(new_n727), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n727), .ZN(new_n887));
  AOI21_X1  g462(.A(KEYINPUT110), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n872), .A2(new_n879), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n886), .A2(KEYINPUT110), .A3(new_n887), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n892), .A2(new_n888), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n893), .B1(new_n872), .B2(new_n879), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n631), .B(G160), .ZN(new_n895));
  NOR3_X1   g470(.A1(new_n891), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n895), .ZN(new_n897));
  NOR3_X1   g472(.A1(new_n870), .A2(new_n871), .A3(new_n864), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n878), .B1(new_n874), .B2(new_n869), .ZN(new_n899));
  OAI22_X1  g474(.A1(new_n898), .A2(new_n899), .B1(new_n888), .B2(new_n892), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n897), .B1(new_n900), .B2(new_n890), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n859), .B1(new_n896), .B2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(KEYINPUT111), .B(G37), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n895), .B1(new_n891), .B2(new_n894), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n900), .A2(new_n897), .A3(new_n890), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n904), .A2(new_n905), .A3(G162), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n902), .A2(new_n903), .A3(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g483(.A1(new_n850), .A2(new_n608), .ZN(new_n909));
  INV_X1    g484(.A(G288), .ZN(new_n910));
  NAND2_X1  g485(.A1(G166), .A2(G305), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n708), .A2(G303), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(G290), .B(KEYINPUT113), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n914), .A2(new_n912), .A3(new_n911), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n910), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n916), .A2(new_n910), .A3(new_n917), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n921), .A2(KEYINPUT42), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT114), .ZN(new_n923));
  INV_X1    g498(.A(new_n920), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n923), .B1(new_n924), .B2(new_n918), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n919), .A2(new_n920), .A3(KEYINPUT114), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n922), .B1(new_n928), .B2(KEYINPUT42), .ZN(new_n929));
  XOR2_X1   g504(.A(new_n855), .B(KEYINPUT112), .Z(new_n930));
  XNOR2_X1  g505(.A(new_n930), .B(new_n614), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n604), .A2(G299), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n600), .A2(new_n765), .A3(new_n601), .A4(new_n603), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n932), .A2(KEYINPUT41), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(KEYINPUT41), .B1(new_n932), .B2(new_n933), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n931), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n932), .A2(new_n933), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n937), .B1(new_n938), .B2(new_n931), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n929), .B(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n909), .B1(new_n940), .B2(new_n608), .ZN(G295));
  OAI21_X1  g516(.A(new_n909), .B1(new_n940), .B2(new_n608), .ZN(G331));
  INV_X1    g517(.A(KEYINPUT116), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT115), .ZN(new_n944));
  INV_X1    g519(.A(new_n544), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n542), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n946), .A2(new_n537), .A3(new_n538), .A4(G301), .ZN(new_n947));
  NAND2_X1  g522(.A1(G286), .A2(G171), .ZN(new_n948));
  AOI211_X1 g523(.A(new_n944), .B(new_n855), .C1(new_n947), .C2(new_n948), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n948), .A2(new_n947), .A3(new_n855), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n855), .B1(new_n948), .B2(new_n947), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n949), .B1(new_n952), .B2(new_n944), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n943), .B1(new_n953), .B2(new_n938), .ZN(new_n954));
  OR3_X1    g529(.A1(new_n934), .A2(new_n935), .A3(new_n952), .ZN(new_n955));
  INV_X1    g530(.A(new_n938), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n950), .A2(new_n951), .A3(KEYINPUT115), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n956), .B(KEYINPUT116), .C1(new_n957), .C2(new_n949), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n954), .A2(new_n955), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n928), .ZN(new_n960));
  INV_X1    g535(.A(G37), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n927), .A2(new_n954), .A3(new_n955), .A4(new_n958), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT43), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AOI22_X1  g540(.A1(new_n936), .A2(new_n953), .B1(new_n956), .B2(new_n952), .ZN(new_n966));
  OR2_X1    g541(.A1(new_n966), .A2(new_n927), .ZN(new_n967));
  AND4_X1   g542(.A1(KEYINPUT43), .A2(new_n967), .A3(new_n903), .A4(new_n962), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT44), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n967), .A2(new_n962), .A3(new_n964), .A4(new_n903), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT44), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n969), .A2(new_n974), .ZN(G397));
  INV_X1    g550(.A(G1384), .ZN(new_n976));
  AOI21_X1  g551(.A(KEYINPUT45), .B1(new_n878), .B2(new_n976), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n476), .A2(G40), .A3(new_n484), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n979), .A2(G1996), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT117), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n980), .B(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT46), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n982), .B(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n793), .B(new_n795), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n758), .A2(new_n759), .A3(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n984), .B1(new_n979), .B2(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n987), .B(KEYINPUT47), .ZN(new_n988));
  INV_X1    g563(.A(G1996), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n760), .A2(new_n989), .ZN(new_n990));
  OR2_X1    g565(.A1(new_n990), .A2(new_n985), .ZN(new_n991));
  INV_X1    g566(.A(new_n979), .ZN(new_n992));
  AOI22_X1  g567(.A1(new_n982), .A2(new_n760), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n726), .A2(new_n729), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n995), .B1(G2067), .B2(new_n867), .ZN(new_n996));
  AND2_X1   g571(.A1(new_n726), .A2(new_n729), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n992), .B1(new_n997), .B2(new_n994), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n993), .A2(new_n998), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n979), .A2(G1986), .A3(G290), .ZN(new_n1000));
  XOR2_X1   g575(.A(new_n1000), .B(KEYINPUT48), .Z(new_n1001));
  AOI22_X1  g576(.A1(new_n996), .A2(new_n992), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n988), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT54), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT50), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n878), .A2(new_n1005), .A3(new_n976), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n860), .A2(new_n875), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n976), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT50), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1006), .A2(new_n978), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT122), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1961), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1006), .A2(KEYINPUT122), .A3(new_n978), .A4(new_n1009), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(G164), .A2(G1384), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT119), .B1(new_n1016), .B2(KEYINPUT45), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n476), .A2(G40), .A3(new_n484), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT119), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT45), .ZN(new_n1020));
  NOR4_X1   g595(.A1(G164), .A2(new_n1019), .A3(new_n1020), .A4(G1384), .ZN(new_n1021));
  NOR4_X1   g596(.A1(new_n977), .A2(new_n1017), .A3(new_n1018), .A4(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1023), .A2(G2078), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n878), .A2(KEYINPUT45), .A3(new_n976), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1008), .A2(new_n1020), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1026), .A2(new_n1027), .A3(new_n978), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1023), .B1(new_n1028), .B2(G2078), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1015), .A2(new_n1025), .A3(new_n1029), .ZN(new_n1030));
  AND2_X1   g605(.A1(new_n1030), .A2(G171), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1020), .B1(new_n864), .B2(G1384), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1032), .A2(new_n1026), .A3(new_n978), .A4(new_n1024), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1015), .A2(new_n1029), .A3(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1034), .A2(G171), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1004), .B1(new_n1031), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(G305), .A2(G1981), .ZN(new_n1037));
  XNOR2_X1  g612(.A(KEYINPUT118), .B(G1981), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n586), .A2(new_n590), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  XNOR2_X1  g615(.A(new_n1040), .B(KEYINPUT49), .ZN(new_n1041));
  INV_X1    g616(.A(G8), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n864), .A2(G1384), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1042), .B1(new_n1043), .B2(new_n978), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1041), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n910), .A2(G1976), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(KEYINPUT52), .ZN(new_n1048));
  INV_X1    g623(.A(G1976), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT52), .B1(G288), .B2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1044), .A2(new_n1046), .A3(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1045), .A2(new_n1048), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1006), .A2(new_n978), .A3(new_n1009), .ZN(new_n1054));
  INV_X1    g629(.A(G2090), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1028), .A2(new_n703), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1042), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(G303), .A2(G8), .ZN(new_n1059));
  XOR2_X1   g634(.A(new_n1059), .B(KEYINPUT55), .Z(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1060), .ZN(new_n1062));
  OAI21_X1  g637(.A(KEYINPUT50), .B1(new_n864), .B2(G1384), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1007), .A2(new_n1005), .A3(new_n976), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1063), .A2(new_n978), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1066), .A2(new_n1055), .B1(new_n1028), .B2(new_n703), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1062), .B1(new_n1067), .B2(new_n1042), .ZN(new_n1068));
  AND3_X1   g643(.A1(new_n1053), .A2(new_n1061), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT51), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1006), .A2(new_n805), .A3(new_n978), .A4(new_n1009), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(new_n1022), .B2(G1966), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1070), .B(G8), .C1(new_n1072), .C2(G286), .ZN(new_n1073));
  NAND2_X1  g648(.A1(G286), .A2(G8), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1019), .B1(new_n1008), .B2(new_n1020), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1021), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1032), .A2(new_n978), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n813), .A2(new_n1077), .B1(new_n1054), .B2(new_n805), .ZN(new_n1078));
  OAI211_X1 g653(.A(KEYINPUT51), .B(new_n1074), .C1(new_n1078), .C2(new_n1042), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1074), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT126), .B1(new_n1072), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT126), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1077), .A2(new_n813), .ZN(new_n1083));
  AOI211_X1 g658(.A(new_n1082), .B(new_n1074), .C1(new_n1083), .C2(new_n1071), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1073), .B(new_n1079), .C1(new_n1081), .C2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1034), .A2(G171), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1086), .B(KEYINPUT54), .C1(G171), .C2(new_n1030), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1036), .A2(new_n1069), .A3(new_n1085), .A4(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1012), .A2(new_n772), .A3(new_n1014), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1043), .A2(new_n795), .A3(new_n978), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT60), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1089), .A2(KEYINPUT60), .A3(new_n1090), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT125), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1094), .A2(new_n1095), .A3(new_n604), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1089), .A2(KEYINPUT125), .A3(KEYINPUT60), .A4(new_n1090), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(new_n605), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1093), .B(new_n1096), .C1(new_n1097), .C2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1043), .A2(new_n978), .ZN(new_n1101));
  XOR2_X1   g676(.A(KEYINPUT58), .B(G1341), .Z(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1026), .A2(new_n989), .A3(new_n1027), .A4(new_n978), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n563), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g680(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1105), .B(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g682(.A(KEYINPUT56), .B(G2072), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1026), .A2(new_n1027), .A3(new_n978), .A4(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(G1956), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT121), .B1(new_n1065), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1005), .B1(new_n878), .B2(new_n976), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n978), .A2(new_n1064), .ZN(new_n1113));
  OAI211_X1 g688(.A(KEYINPUT121), .B(new_n1110), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1109), .B1(new_n1111), .B2(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g691(.A(G299), .B(KEYINPUT57), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1110), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT121), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n1114), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1117), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1122), .A2(new_n1123), .A3(new_n1109), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1118), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT61), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1107), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1123), .B1(new_n1122), .B2(new_n1109), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1109), .ZN(new_n1129));
  AOI211_X1 g704(.A(new_n1117), .B(new_n1129), .C1(new_n1121), .C2(new_n1114), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT124), .B1(new_n1131), .B2(KEYINPUT61), .ZN(new_n1132));
  AND4_X1   g707(.A1(KEYINPUT124), .A2(new_n1118), .A3(KEYINPUT61), .A4(new_n1124), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1100), .B(new_n1127), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n604), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1124), .B1(new_n1128), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1088), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1069), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1085), .A2(KEYINPUT62), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1082), .B1(new_n1078), .B2(new_n1074), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1072), .A2(KEYINPUT126), .A3(new_n1080), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT62), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1142), .A2(new_n1143), .A3(new_n1073), .A4(new_n1079), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1139), .A2(new_n1031), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT63), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1078), .A2(new_n1042), .ZN(new_n1147));
  AOI21_X1  g722(.A(KEYINPUT120), .B1(new_n1147), .B2(G168), .ZN(new_n1148));
  AND4_X1   g723(.A1(KEYINPUT120), .A2(new_n1072), .A3(G8), .A4(G168), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1146), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1138), .B1(new_n1145), .B2(new_n1150), .ZN(new_n1151));
  OR2_X1    g726(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1152), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1053), .A2(new_n1061), .ZN(new_n1154));
  OAI21_X1  g729(.A(KEYINPUT63), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  OR2_X1    g730(.A1(new_n1061), .A2(new_n1052), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1045), .A2(new_n1049), .A3(new_n910), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(new_n1039), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(new_n1044), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1155), .A2(new_n1156), .A3(new_n1159), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n1137), .A2(new_n1151), .A3(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g736(.A(G290), .B(new_n716), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n999), .B1(new_n979), .B2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1003), .B1(new_n1161), .B2(new_n1163), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g739(.A(G229), .ZN(new_n1166));
  NAND3_X1  g740(.A1(new_n650), .A2(G319), .A3(new_n671), .ZN(new_n1167));
  OAI21_X1  g741(.A(new_n1166), .B1(new_n1167), .B2(KEYINPUT127), .ZN(new_n1168));
  AOI21_X1  g742(.A(new_n1168), .B1(KEYINPUT127), .B2(new_n1167), .ZN(new_n1169));
  NAND3_X1  g743(.A1(new_n972), .A2(new_n907), .A3(new_n1169), .ZN(G225));
  INV_X1    g744(.A(G225), .ZN(G308));
endmodule


