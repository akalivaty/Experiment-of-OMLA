

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U550 ( .A(KEYINPUT1), .B(n543), .Z(n653) );
  AND2_X1 U551 ( .A1(G1348), .A2(n983), .ZN(n692) );
  NAND2_X1 U552 ( .A1(n718), .A2(n514), .ZN(n720) );
  XOR2_X1 U553 ( .A(n717), .B(KEYINPUT28), .Z(n514) );
  OR2_X1 U554 ( .A1(n739), .A2(n707), .ZN(n708) );
  NOR2_X1 U555 ( .A1(n694), .A2(n721), .ZN(n695) );
  INV_X1 U556 ( .A(KEYINPUT29), .ZN(n719) );
  INV_X1 U557 ( .A(KEYINPUT99), .ZN(n767) );
  INV_X1 U558 ( .A(KEYINPUT101), .ZN(n817) );
  NOR2_X1 U559 ( .A1(G651), .A2(n637), .ZN(n545) );
  NAND2_X1 U560 ( .A1(n585), .A2(n584), .ZN(n587) );
  AND2_X1 U561 ( .A1(n527), .A2(n526), .ZN(G160) );
  INV_X1 U562 ( .A(KEYINPUT66), .ZN(n519) );
  NOR2_X1 U563 ( .A1(G2104), .A2(G2105), .ZN(n515) );
  XOR2_X2 U564 ( .A(KEYINPUT17), .B(n515), .Z(n893) );
  NAND2_X1 U565 ( .A1(G137), .A2(n893), .ZN(n517) );
  AND2_X1 U566 ( .A1(G2104), .A2(G2105), .ZN(n885) );
  NAND2_X1 U567 ( .A1(G113), .A2(n885), .ZN(n516) );
  NAND2_X1 U568 ( .A1(n517), .A2(n516), .ZN(n518) );
  OR2_X1 U569 ( .A1(n519), .A2(n518), .ZN(n521) );
  NAND2_X1 U570 ( .A1(n519), .A2(n518), .ZN(n520) );
  NAND2_X1 U571 ( .A1(n521), .A2(n520), .ZN(n527) );
  INV_X1 U572 ( .A(G2105), .ZN(n523) );
  AND2_X1 U573 ( .A1(n523), .A2(G2104), .ZN(n890) );
  NAND2_X1 U574 ( .A1(G101), .A2(n890), .ZN(n522) );
  XOR2_X1 U575 ( .A(KEYINPUT23), .B(n522), .Z(n525) );
  NOR2_X1 U576 ( .A1(G2104), .A2(n523), .ZN(n886) );
  NAND2_X1 U577 ( .A1(n886), .A2(G125), .ZN(n524) );
  AND2_X1 U578 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U579 ( .A(G2443), .B(G2446), .Z(n529) );
  XNOR2_X1 U580 ( .A(G2427), .B(G2451), .ZN(n528) );
  XNOR2_X1 U581 ( .A(n529), .B(n528), .ZN(n535) );
  XOR2_X1 U582 ( .A(G2430), .B(G2454), .Z(n531) );
  XNOR2_X1 U583 ( .A(G1348), .B(G1341), .ZN(n530) );
  XNOR2_X1 U584 ( .A(n531), .B(n530), .ZN(n533) );
  XOR2_X1 U585 ( .A(G2435), .B(G2438), .Z(n532) );
  XNOR2_X1 U586 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U587 ( .A(n535), .B(n534), .Z(n536) );
  AND2_X1 U588 ( .A1(G14), .A2(n536), .ZN(G401) );
  XNOR2_X1 U589 ( .A(KEYINPUT9), .B(KEYINPUT70), .ZN(n541) );
  XOR2_X1 U590 ( .A(G543), .B(KEYINPUT0), .Z(n637) );
  INV_X1 U591 ( .A(G651), .ZN(n542) );
  NOR2_X1 U592 ( .A1(n637), .A2(n542), .ZN(n658) );
  NAND2_X1 U593 ( .A1(n658), .A2(G77), .ZN(n539) );
  NOR2_X1 U594 ( .A1(G651), .A2(G543), .ZN(n654) );
  NAND2_X1 U595 ( .A1(n654), .A2(G90), .ZN(n537) );
  XOR2_X1 U596 ( .A(KEYINPUT69), .B(n537), .Z(n538) );
  NAND2_X1 U597 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U598 ( .A(n541), .B(n540), .Z(n550) );
  NOR2_X1 U599 ( .A1(G543), .A2(n542), .ZN(n543) );
  NAND2_X1 U600 ( .A1(n653), .A2(G64), .ZN(n544) );
  XOR2_X1 U601 ( .A(KEYINPUT67), .B(n544), .Z(n547) );
  XOR2_X1 U602 ( .A(KEYINPUT65), .B(n545), .Z(n652) );
  NAND2_X1 U603 ( .A1(n652), .A2(G52), .ZN(n546) );
  NAND2_X1 U604 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U605 ( .A(KEYINPUT68), .B(n548), .ZN(n549) );
  NOR2_X1 U606 ( .A1(n550), .A2(n549), .ZN(G171) );
  NAND2_X1 U607 ( .A1(G65), .A2(n653), .ZN(n552) );
  NAND2_X1 U608 ( .A1(G53), .A2(n652), .ZN(n551) );
  NAND2_X1 U609 ( .A1(n552), .A2(n551), .ZN(n556) );
  NAND2_X1 U610 ( .A1(G91), .A2(n654), .ZN(n554) );
  NAND2_X1 U611 ( .A1(G78), .A2(n658), .ZN(n553) );
  NAND2_X1 U612 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U613 ( .A1(n556), .A2(n555), .ZN(n715) );
  INV_X1 U614 ( .A(n715), .ZN(G299) );
  INV_X1 U615 ( .A(G57), .ZN(G237) );
  INV_X1 U616 ( .A(G132), .ZN(G219) );
  INV_X1 U617 ( .A(G82), .ZN(G220) );
  NAND2_X1 U618 ( .A1(G102), .A2(n890), .ZN(n558) );
  NAND2_X1 U619 ( .A1(G138), .A2(n893), .ZN(n557) );
  NAND2_X1 U620 ( .A1(n558), .A2(n557), .ZN(n562) );
  NAND2_X1 U621 ( .A1(G114), .A2(n885), .ZN(n560) );
  NAND2_X1 U622 ( .A1(G126), .A2(n886), .ZN(n559) );
  NAND2_X1 U623 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U624 ( .A1(n562), .A2(n561), .ZN(G164) );
  NAND2_X1 U625 ( .A1(G94), .A2(G452), .ZN(n563) );
  XNOR2_X1 U626 ( .A(n563), .B(KEYINPUT71), .ZN(G173) );
  NAND2_X1 U627 ( .A1(G7), .A2(G661), .ZN(n564) );
  XNOR2_X1 U628 ( .A(n564), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U629 ( .A(G223), .ZN(n837) );
  NAND2_X1 U630 ( .A1(n837), .A2(G567), .ZN(n565) );
  XOR2_X1 U631 ( .A(KEYINPUT11), .B(n565), .Z(G234) );
  NAND2_X1 U632 ( .A1(n653), .A2(G56), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n566), .B(KEYINPUT14), .ZN(n568) );
  NAND2_X1 U634 ( .A1(G43), .A2(n652), .ZN(n567) );
  NAND2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n575) );
  NAND2_X1 U636 ( .A1(n654), .A2(G81), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n569), .B(KEYINPUT12), .ZN(n571) );
  NAND2_X1 U638 ( .A1(G68), .A2(n658), .ZN(n570) );
  NAND2_X1 U639 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U640 ( .A(KEYINPUT72), .B(n572), .Z(n573) );
  XNOR2_X1 U641 ( .A(KEYINPUT13), .B(n573), .ZN(n574) );
  NOR2_X1 U642 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U643 ( .A(KEYINPUT73), .B(n576), .ZN(n989) );
  INV_X1 U644 ( .A(G860), .ZN(n622) );
  OR2_X1 U645 ( .A1(n989), .A2(n622), .ZN(G153) );
  XOR2_X1 U646 ( .A(G171), .B(KEYINPUT74), .Z(G301) );
  NAND2_X1 U647 ( .A1(G868), .A2(G301), .ZN(n589) );
  NAND2_X1 U648 ( .A1(G79), .A2(n658), .ZN(n577) );
  XNOR2_X1 U649 ( .A(n577), .B(KEYINPUT76), .ZN(n585) );
  NAND2_X1 U650 ( .A1(n652), .A2(G54), .ZN(n579) );
  NAND2_X1 U651 ( .A1(G92), .A2(n654), .ZN(n578) );
  NAND2_X1 U652 ( .A1(n579), .A2(n578), .ZN(n583) );
  INV_X1 U653 ( .A(KEYINPUT75), .ZN(n581) );
  AND2_X1 U654 ( .A1(G66), .A2(n653), .ZN(n580) );
  XNOR2_X1 U655 ( .A(n581), .B(n580), .ZN(n582) );
  NOR2_X1 U656 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U657 ( .A(KEYINPUT77), .B(KEYINPUT15), .ZN(n586) );
  XNOR2_X2 U658 ( .A(n587), .B(n586), .ZN(n983) );
  INV_X1 U659 ( .A(G868), .ZN(n672) );
  NAND2_X1 U660 ( .A1(n983), .A2(n672), .ZN(n588) );
  NAND2_X1 U661 ( .A1(n589), .A2(n588), .ZN(G284) );
  NAND2_X1 U662 ( .A1(G89), .A2(n654), .ZN(n590) );
  XNOR2_X1 U663 ( .A(n590), .B(KEYINPUT78), .ZN(n591) );
  XNOR2_X1 U664 ( .A(n591), .B(KEYINPUT4), .ZN(n593) );
  NAND2_X1 U665 ( .A1(G76), .A2(n658), .ZN(n592) );
  NAND2_X1 U666 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U667 ( .A(n594), .B(KEYINPUT5), .ZN(n599) );
  NAND2_X1 U668 ( .A1(G63), .A2(n653), .ZN(n596) );
  NAND2_X1 U669 ( .A1(G51), .A2(n652), .ZN(n595) );
  NAND2_X1 U670 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U671 ( .A(KEYINPUT6), .B(n597), .Z(n598) );
  NAND2_X1 U672 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U673 ( .A(n600), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U674 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U675 ( .A1(G286), .A2(n672), .ZN(n602) );
  NOR2_X1 U676 ( .A1(G868), .A2(G299), .ZN(n601) );
  NOR2_X1 U677 ( .A1(n602), .A2(n601), .ZN(G297) );
  NAND2_X1 U678 ( .A1(n622), .A2(G559), .ZN(n603) );
  INV_X1 U679 ( .A(n983), .ZN(n620) );
  NAND2_X1 U680 ( .A1(n603), .A2(n620), .ZN(n604) );
  XNOR2_X1 U681 ( .A(n604), .B(KEYINPUT79), .ZN(n605) );
  XOR2_X1 U682 ( .A(KEYINPUT16), .B(n605), .Z(G148) );
  OR2_X1 U683 ( .A1(G559), .A2(n983), .ZN(n606) );
  NAND2_X1 U684 ( .A1(n606), .A2(G868), .ZN(n608) );
  NAND2_X1 U685 ( .A1(n989), .A2(n672), .ZN(n607) );
  NAND2_X1 U686 ( .A1(n608), .A2(n607), .ZN(G282) );
  NAND2_X1 U687 ( .A1(G99), .A2(n890), .ZN(n610) );
  NAND2_X1 U688 ( .A1(G111), .A2(n885), .ZN(n609) );
  NAND2_X1 U689 ( .A1(n610), .A2(n609), .ZN(n617) );
  NAND2_X1 U690 ( .A1(G123), .A2(n886), .ZN(n611) );
  XNOR2_X1 U691 ( .A(n611), .B(KEYINPUT18), .ZN(n612) );
  XNOR2_X1 U692 ( .A(n612), .B(KEYINPUT80), .ZN(n614) );
  NAND2_X1 U693 ( .A1(G135), .A2(n893), .ZN(n613) );
  NAND2_X1 U694 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U695 ( .A(KEYINPUT81), .B(n615), .Z(n616) );
  NOR2_X1 U696 ( .A1(n617), .A2(n616), .ZN(n925) );
  XNOR2_X1 U697 ( .A(G2096), .B(n925), .ZN(n619) );
  INV_X1 U698 ( .A(G2100), .ZN(n618) );
  NAND2_X1 U699 ( .A1(n619), .A2(n618), .ZN(G156) );
  XOR2_X1 U700 ( .A(KEYINPUT82), .B(KEYINPUT85), .Z(n624) );
  NAND2_X1 U701 ( .A1(G559), .A2(n620), .ZN(n621) );
  XOR2_X1 U702 ( .A(n989), .B(n621), .Z(n670) );
  NAND2_X1 U703 ( .A1(n670), .A2(n622), .ZN(n623) );
  XNOR2_X1 U704 ( .A(n624), .B(n623), .ZN(n633) );
  NAND2_X1 U705 ( .A1(G55), .A2(n652), .ZN(n625) );
  XNOR2_X1 U706 ( .A(n625), .B(KEYINPUT84), .ZN(n632) );
  NAND2_X1 U707 ( .A1(G67), .A2(n653), .ZN(n627) );
  NAND2_X1 U708 ( .A1(G93), .A2(n654), .ZN(n626) );
  NAND2_X1 U709 ( .A1(n627), .A2(n626), .ZN(n630) );
  NAND2_X1 U710 ( .A1(G80), .A2(n658), .ZN(n628) );
  XNOR2_X1 U711 ( .A(KEYINPUT83), .B(n628), .ZN(n629) );
  NOR2_X1 U712 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U713 ( .A1(n632), .A2(n631), .ZN(n673) );
  XNOR2_X1 U714 ( .A(n633), .B(n673), .ZN(G145) );
  NAND2_X1 U715 ( .A1(G49), .A2(n652), .ZN(n635) );
  NAND2_X1 U716 ( .A1(G74), .A2(G651), .ZN(n634) );
  NAND2_X1 U717 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U718 ( .A1(n653), .A2(n636), .ZN(n639) );
  NAND2_X1 U719 ( .A1(n637), .A2(G87), .ZN(n638) );
  NAND2_X1 U720 ( .A1(n639), .A2(n638), .ZN(G288) );
  NAND2_X1 U721 ( .A1(G88), .A2(n654), .ZN(n641) );
  NAND2_X1 U722 ( .A1(G75), .A2(n658), .ZN(n640) );
  NAND2_X1 U723 ( .A1(n641), .A2(n640), .ZN(n645) );
  NAND2_X1 U724 ( .A1(G62), .A2(n653), .ZN(n643) );
  NAND2_X1 U725 ( .A1(G50), .A2(n652), .ZN(n642) );
  NAND2_X1 U726 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U727 ( .A1(n645), .A2(n644), .ZN(G166) );
  AND2_X1 U728 ( .A1(n653), .A2(G60), .ZN(n649) );
  NAND2_X1 U729 ( .A1(G47), .A2(n652), .ZN(n647) );
  NAND2_X1 U730 ( .A1(G85), .A2(n654), .ZN(n646) );
  NAND2_X1 U731 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U732 ( .A1(n649), .A2(n648), .ZN(n651) );
  NAND2_X1 U733 ( .A1(n658), .A2(G72), .ZN(n650) );
  NAND2_X1 U734 ( .A1(n651), .A2(n650), .ZN(G290) );
  NAND2_X1 U735 ( .A1(n652), .A2(G48), .ZN(n663) );
  NAND2_X1 U736 ( .A1(G61), .A2(n653), .ZN(n656) );
  NAND2_X1 U737 ( .A1(G86), .A2(n654), .ZN(n655) );
  NAND2_X1 U738 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U739 ( .A(KEYINPUT86), .B(n657), .ZN(n661) );
  NAND2_X1 U740 ( .A1(n658), .A2(G73), .ZN(n659) );
  XOR2_X1 U741 ( .A(KEYINPUT2), .B(n659), .Z(n660) );
  NOR2_X1 U742 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U743 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U744 ( .A(KEYINPUT87), .B(n664), .Z(G305) );
  XNOR2_X1 U745 ( .A(G288), .B(KEYINPUT19), .ZN(n666) );
  XNOR2_X1 U746 ( .A(n715), .B(G166), .ZN(n665) );
  XNOR2_X1 U747 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U748 ( .A(n667), .B(G290), .ZN(n668) );
  XNOR2_X1 U749 ( .A(n668), .B(n673), .ZN(n669) );
  XNOR2_X1 U750 ( .A(n669), .B(G305), .ZN(n910) );
  XNOR2_X1 U751 ( .A(n670), .B(n910), .ZN(n671) );
  NAND2_X1 U752 ( .A1(n671), .A2(G868), .ZN(n675) );
  NAND2_X1 U753 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U754 ( .A1(n675), .A2(n674), .ZN(G295) );
  XOR2_X1 U755 ( .A(KEYINPUT20), .B(KEYINPUT88), .Z(n677) );
  NAND2_X1 U756 ( .A1(G2084), .A2(G2078), .ZN(n676) );
  XNOR2_X1 U757 ( .A(n677), .B(n676), .ZN(n678) );
  NAND2_X1 U758 ( .A1(G2090), .A2(n678), .ZN(n679) );
  XNOR2_X1 U759 ( .A(KEYINPUT21), .B(n679), .ZN(n680) );
  NAND2_X1 U760 ( .A1(n680), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U761 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U762 ( .A1(G220), .A2(G219), .ZN(n681) );
  XOR2_X1 U763 ( .A(KEYINPUT22), .B(n681), .Z(n682) );
  NOR2_X1 U764 ( .A1(G218), .A2(n682), .ZN(n683) );
  NAND2_X1 U765 ( .A1(G96), .A2(n683), .ZN(n842) );
  NAND2_X1 U766 ( .A1(G2106), .A2(n842), .ZN(n687) );
  NAND2_X1 U767 ( .A1(G108), .A2(G120), .ZN(n684) );
  NOR2_X1 U768 ( .A1(G237), .A2(n684), .ZN(n685) );
  NAND2_X1 U769 ( .A1(G69), .A2(n685), .ZN(n843) );
  NAND2_X1 U770 ( .A1(G567), .A2(n843), .ZN(n686) );
  NAND2_X1 U771 ( .A1(n687), .A2(n686), .ZN(n864) );
  NAND2_X1 U772 ( .A1(G661), .A2(G483), .ZN(n688) );
  XOR2_X1 U773 ( .A(KEYINPUT89), .B(n688), .Z(n689) );
  NOR2_X1 U774 ( .A1(n864), .A2(n689), .ZN(n841) );
  NAND2_X1 U775 ( .A1(n841), .A2(G36), .ZN(G176) );
  INV_X1 U776 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U777 ( .A(KEYINPUT64), .B(KEYINPUT26), .ZN(n696) );
  INV_X1 U778 ( .A(G1341), .ZN(n690) );
  NAND2_X1 U779 ( .A1(n696), .A2(n690), .ZN(n691) );
  NOR2_X1 U780 ( .A1(n692), .A2(n691), .ZN(n694) );
  NOR2_X1 U781 ( .A1(G164), .A2(G1384), .ZN(n785) );
  AND2_X1 U782 ( .A1(n785), .A2(G40), .ZN(n693) );
  NAND2_X1 U783 ( .A1(G160), .A2(n693), .ZN(n739) );
  INV_X1 U784 ( .A(n739), .ZN(n721) );
  NOR2_X1 U785 ( .A1(n695), .A2(n989), .ZN(n703) );
  OR2_X1 U786 ( .A1(G1996), .A2(n696), .ZN(n701) );
  NAND2_X1 U787 ( .A1(G2067), .A2(n983), .ZN(n698) );
  NAND2_X1 U788 ( .A1(G1996), .A2(n696), .ZN(n697) );
  NAND2_X1 U789 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U790 ( .A1(n699), .A2(n721), .ZN(n700) );
  AND2_X1 U791 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U792 ( .A1(n703), .A2(n702), .ZN(n714) );
  NAND2_X1 U793 ( .A1(G1348), .A2(n739), .ZN(n705) );
  NAND2_X1 U794 ( .A1(G2067), .A2(n721), .ZN(n704) );
  NAND2_X1 U795 ( .A1(n705), .A2(n704), .ZN(n706) );
  OR2_X1 U796 ( .A1(n706), .A2(n983), .ZN(n712) );
  INV_X1 U797 ( .A(G2072), .ZN(n707) );
  XNOR2_X1 U798 ( .A(n708), .B(KEYINPUT27), .ZN(n710) );
  AND2_X1 U799 ( .A1(G1956), .A2(n739), .ZN(n709) );
  NOR2_X1 U800 ( .A1(n710), .A2(n709), .ZN(n716) );
  NAND2_X1 U801 ( .A1(n716), .A2(n715), .ZN(n711) );
  AND2_X1 U802 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U803 ( .A1(n714), .A2(n713), .ZN(n718) );
  NOR2_X1 U804 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U805 ( .A(n720), .B(n719), .ZN(n726) );
  INV_X1 U806 ( .A(G1961), .ZN(n996) );
  NAND2_X1 U807 ( .A1(n739), .A2(n996), .ZN(n723) );
  XNOR2_X1 U808 ( .A(G2078), .B(KEYINPUT25), .ZN(n952) );
  NAND2_X1 U809 ( .A1(n721), .A2(n952), .ZN(n722) );
  NAND2_X1 U810 ( .A1(n723), .A2(n722), .ZN(n727) );
  NAND2_X1 U811 ( .A1(G171), .A2(n727), .ZN(n724) );
  XOR2_X1 U812 ( .A(KEYINPUT95), .B(n724), .Z(n725) );
  NAND2_X1 U813 ( .A1(n726), .A2(n725), .ZN(n737) );
  XNOR2_X1 U814 ( .A(KEYINPUT31), .B(KEYINPUT97), .ZN(n735) );
  NOR2_X1 U815 ( .A1(G171), .A2(n727), .ZN(n728) );
  XNOR2_X1 U816 ( .A(n728), .B(KEYINPUT96), .ZN(n733) );
  NAND2_X1 U817 ( .A1(G8), .A2(n739), .ZN(n779) );
  NOR2_X1 U818 ( .A1(G1966), .A2(n779), .ZN(n750) );
  NOR2_X1 U819 ( .A1(G2084), .A2(n739), .ZN(n747) );
  NOR2_X1 U820 ( .A1(n750), .A2(n747), .ZN(n729) );
  NAND2_X1 U821 ( .A1(G8), .A2(n729), .ZN(n730) );
  XNOR2_X1 U822 ( .A(KEYINPUT30), .B(n730), .ZN(n731) );
  NOR2_X1 U823 ( .A1(n731), .A2(G168), .ZN(n732) );
  NOR2_X1 U824 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U825 ( .A(n735), .B(n734), .ZN(n736) );
  NAND2_X1 U826 ( .A1(n737), .A2(n736), .ZN(n748) );
  NAND2_X1 U827 ( .A1(n748), .A2(G286), .ZN(n738) );
  XNOR2_X1 U828 ( .A(n738), .B(KEYINPUT98), .ZN(n744) );
  NOR2_X1 U829 ( .A1(G1971), .A2(n779), .ZN(n741) );
  NOR2_X1 U830 ( .A1(G2090), .A2(n739), .ZN(n740) );
  NOR2_X1 U831 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U832 ( .A1(n742), .A2(G303), .ZN(n743) );
  NAND2_X1 U833 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U834 ( .A1(n745), .A2(G8), .ZN(n746) );
  XNOR2_X1 U835 ( .A(n746), .B(KEYINPUT32), .ZN(n771) );
  NAND2_X1 U836 ( .A1(G8), .A2(n747), .ZN(n752) );
  INV_X1 U837 ( .A(n748), .ZN(n749) );
  NOR2_X1 U838 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U839 ( .A1(n752), .A2(n751), .ZN(n772) );
  NAND2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n976) );
  AND2_X1 U841 ( .A1(n772), .A2(n976), .ZN(n754) );
  OR2_X1 U842 ( .A1(n779), .A2(KEYINPUT33), .ZN(n762) );
  INV_X1 U843 ( .A(n762), .ZN(n753) );
  AND2_X1 U844 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U845 ( .A1(n771), .A2(n755), .ZN(n766) );
  NOR2_X1 U846 ( .A1(G1976), .A2(G288), .ZN(n759) );
  INV_X1 U847 ( .A(n779), .ZN(n756) );
  NAND2_X1 U848 ( .A1(n759), .A2(n756), .ZN(n757) );
  NAND2_X1 U849 ( .A1(n757), .A2(KEYINPUT33), .ZN(n764) );
  INV_X1 U850 ( .A(n976), .ZN(n760) );
  NOR2_X1 U851 ( .A1(G1971), .A2(G303), .ZN(n758) );
  NOR2_X1 U852 ( .A1(n759), .A2(n758), .ZN(n980) );
  OR2_X1 U853 ( .A1(n760), .A2(n980), .ZN(n761) );
  OR2_X1 U854 ( .A1(n762), .A2(n761), .ZN(n763) );
  AND2_X1 U855 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U856 ( .A1(n766), .A2(n765), .ZN(n768) );
  XNOR2_X1 U857 ( .A(n768), .B(n767), .ZN(n769) );
  XOR2_X1 U858 ( .A(G1981), .B(G305), .Z(n972) );
  NAND2_X1 U859 ( .A1(n769), .A2(n972), .ZN(n770) );
  XNOR2_X1 U860 ( .A(n770), .B(KEYINPUT100), .ZN(n783) );
  NAND2_X1 U861 ( .A1(n772), .A2(n771), .ZN(n775) );
  NOR2_X1 U862 ( .A1(G2090), .A2(G303), .ZN(n773) );
  NAND2_X1 U863 ( .A1(G8), .A2(n773), .ZN(n774) );
  NAND2_X1 U864 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U865 ( .A1(n776), .A2(n779), .ZN(n781) );
  NOR2_X1 U866 ( .A1(G1981), .A2(G305), .ZN(n777) );
  XOR2_X1 U867 ( .A(n777), .B(KEYINPUT24), .Z(n778) );
  NOR2_X1 U868 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X1 U869 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n816) );
  NAND2_X1 U871 ( .A1(G160), .A2(G40), .ZN(n784) );
  NOR2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n832) );
  NAND2_X1 U873 ( .A1(n893), .A2(G140), .ZN(n786) );
  XNOR2_X1 U874 ( .A(n786), .B(KEYINPUT90), .ZN(n788) );
  NAND2_X1 U875 ( .A1(G104), .A2(n890), .ZN(n787) );
  NAND2_X1 U876 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U877 ( .A(KEYINPUT34), .B(n789), .ZN(n795) );
  NAND2_X1 U878 ( .A1(n886), .A2(G128), .ZN(n790) );
  XOR2_X1 U879 ( .A(KEYINPUT91), .B(n790), .Z(n792) );
  NAND2_X1 U880 ( .A1(n885), .A2(G116), .ZN(n791) );
  NAND2_X1 U881 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U882 ( .A(n793), .B(KEYINPUT35), .Z(n794) );
  NOR2_X1 U883 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U884 ( .A(KEYINPUT36), .B(n796), .Z(n797) );
  XOR2_X1 U885 ( .A(KEYINPUT92), .B(n797), .Z(n908) );
  XNOR2_X1 U886 ( .A(G2067), .B(KEYINPUT37), .ZN(n821) );
  NOR2_X1 U887 ( .A1(n908), .A2(n821), .ZN(n946) );
  NAND2_X1 U888 ( .A1(n832), .A2(n946), .ZN(n829) );
  NAND2_X1 U889 ( .A1(G141), .A2(n893), .ZN(n798) );
  XNOR2_X1 U890 ( .A(n798), .B(KEYINPUT94), .ZN(n805) );
  NAND2_X1 U891 ( .A1(G117), .A2(n885), .ZN(n800) );
  NAND2_X1 U892 ( .A1(G129), .A2(n886), .ZN(n799) );
  NAND2_X1 U893 ( .A1(n800), .A2(n799), .ZN(n803) );
  NAND2_X1 U894 ( .A1(n890), .A2(G105), .ZN(n801) );
  XOR2_X1 U895 ( .A(KEYINPUT38), .B(n801), .Z(n802) );
  NOR2_X1 U896 ( .A1(n803), .A2(n802), .ZN(n804) );
  NAND2_X1 U897 ( .A1(n805), .A2(n804), .ZN(n897) );
  NAND2_X1 U898 ( .A1(G1996), .A2(n897), .ZN(n814) );
  NAND2_X1 U899 ( .A1(G95), .A2(n890), .ZN(n807) );
  NAND2_X1 U900 ( .A1(G107), .A2(n885), .ZN(n806) );
  NAND2_X1 U901 ( .A1(n807), .A2(n806), .ZN(n810) );
  NAND2_X1 U902 ( .A1(G119), .A2(n886), .ZN(n808) );
  XNOR2_X1 U903 ( .A(KEYINPUT93), .B(n808), .ZN(n809) );
  NOR2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n812) );
  NAND2_X1 U905 ( .A1(n893), .A2(G131), .ZN(n811) );
  NAND2_X1 U906 ( .A1(n812), .A2(n811), .ZN(n898) );
  NAND2_X1 U907 ( .A1(G1991), .A2(n898), .ZN(n813) );
  NAND2_X1 U908 ( .A1(n814), .A2(n813), .ZN(n924) );
  NAND2_X1 U909 ( .A1(n832), .A2(n924), .ZN(n825) );
  AND2_X1 U910 ( .A1(n829), .A2(n825), .ZN(n815) );
  AND2_X1 U911 ( .A1(n816), .A2(n815), .ZN(n818) );
  XNOR2_X1 U912 ( .A(n818), .B(n817), .ZN(n820) );
  XNOR2_X1 U913 ( .A(G1986), .B(G290), .ZN(n982) );
  NAND2_X1 U914 ( .A1(n982), .A2(n832), .ZN(n819) );
  NAND2_X1 U915 ( .A1(n820), .A2(n819), .ZN(n835) );
  NAND2_X1 U916 ( .A1(n908), .A2(n821), .ZN(n943) );
  NOR2_X1 U917 ( .A1(G1986), .A2(G290), .ZN(n823) );
  NOR2_X1 U918 ( .A1(n898), .A2(G1991), .ZN(n822) );
  XNOR2_X1 U919 ( .A(n822), .B(KEYINPUT102), .ZN(n934) );
  NOR2_X1 U920 ( .A1(n823), .A2(n934), .ZN(n824) );
  XNOR2_X1 U921 ( .A(n824), .B(KEYINPUT103), .ZN(n826) );
  NAND2_X1 U922 ( .A1(n826), .A2(n825), .ZN(n827) );
  OR2_X1 U923 ( .A1(n897), .A2(G1996), .ZN(n937) );
  NAND2_X1 U924 ( .A1(n827), .A2(n937), .ZN(n828) );
  XOR2_X1 U925 ( .A(KEYINPUT39), .B(n828), .Z(n830) );
  NAND2_X1 U926 ( .A1(n830), .A2(n829), .ZN(n831) );
  NAND2_X1 U927 ( .A1(n943), .A2(n831), .ZN(n833) );
  NAND2_X1 U928 ( .A1(n833), .A2(n832), .ZN(n834) );
  NAND2_X1 U929 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U930 ( .A(KEYINPUT40), .B(n836), .ZN(G329) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n837), .ZN(G217) );
  NAND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n838) );
  XOR2_X1 U933 ( .A(KEYINPUT104), .B(n838), .Z(n839) );
  NAND2_X1 U934 ( .A1(G661), .A2(n839), .ZN(G259) );
  NAND2_X1 U935 ( .A1(G3), .A2(G1), .ZN(n840) );
  NAND2_X1 U936 ( .A1(n841), .A2(n840), .ZN(G188) );
  XNOR2_X1 U937 ( .A(G120), .B(KEYINPUT105), .ZN(G236) );
  INV_X1 U939 ( .A(G108), .ZN(G238) );
  INV_X1 U940 ( .A(G96), .ZN(G221) );
  NOR2_X1 U941 ( .A1(n843), .A2(n842), .ZN(G325) );
  INV_X1 U942 ( .A(G325), .ZN(G261) );
  XOR2_X1 U943 ( .A(KEYINPUT107), .B(G2084), .Z(n845) );
  XNOR2_X1 U944 ( .A(G2078), .B(G2072), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U946 ( .A(n846), .B(G2096), .Z(n848) );
  XNOR2_X1 U947 ( .A(G2067), .B(G2090), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U949 ( .A(KEYINPUT43), .B(G2678), .Z(n850) );
  XNOR2_X1 U950 ( .A(KEYINPUT42), .B(G2100), .ZN(n849) );
  XNOR2_X1 U951 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U952 ( .A(n852), .B(n851), .Z(G227) );
  XOR2_X1 U953 ( .A(KEYINPUT109), .B(G1981), .Z(n854) );
  XNOR2_X1 U954 ( .A(G1986), .B(G1966), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U956 ( .A(n855), .B(KEYINPUT41), .Z(n857) );
  XNOR2_X1 U957 ( .A(G1996), .B(G1991), .ZN(n856) );
  XNOR2_X1 U958 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U959 ( .A(G1976), .B(G1971), .Z(n859) );
  XNOR2_X1 U960 ( .A(G1961), .B(G1956), .ZN(n858) );
  XNOR2_X1 U961 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U962 ( .A(n861), .B(n860), .Z(n863) );
  XNOR2_X1 U963 ( .A(KEYINPUT108), .B(G2474), .ZN(n862) );
  XNOR2_X1 U964 ( .A(n863), .B(n862), .ZN(G229) );
  XOR2_X1 U965 ( .A(KEYINPUT106), .B(n864), .Z(G319) );
  NAND2_X1 U966 ( .A1(n890), .A2(G100), .ZN(n865) );
  XOR2_X1 U967 ( .A(KEYINPUT111), .B(n865), .Z(n867) );
  NAND2_X1 U968 ( .A1(n885), .A2(G112), .ZN(n866) );
  NAND2_X1 U969 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U970 ( .A(KEYINPUT112), .B(n868), .ZN(n874) );
  NAND2_X1 U971 ( .A1(G124), .A2(n886), .ZN(n869) );
  XNOR2_X1 U972 ( .A(n869), .B(KEYINPUT110), .ZN(n870) );
  XNOR2_X1 U973 ( .A(n870), .B(KEYINPUT44), .ZN(n872) );
  NAND2_X1 U974 ( .A1(G136), .A2(n893), .ZN(n871) );
  NAND2_X1 U975 ( .A1(n872), .A2(n871), .ZN(n873) );
  NOR2_X1 U976 ( .A1(n874), .A2(n873), .ZN(G162) );
  NAND2_X1 U977 ( .A1(G118), .A2(n885), .ZN(n876) );
  NAND2_X1 U978 ( .A1(G130), .A2(n886), .ZN(n875) );
  NAND2_X1 U979 ( .A1(n876), .A2(n875), .ZN(n881) );
  NAND2_X1 U980 ( .A1(G106), .A2(n890), .ZN(n878) );
  NAND2_X1 U981 ( .A1(G142), .A2(n893), .ZN(n877) );
  NAND2_X1 U982 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U983 ( .A(KEYINPUT45), .B(n879), .Z(n880) );
  NOR2_X1 U984 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U985 ( .A(n882), .B(n925), .Z(n884) );
  XNOR2_X1 U986 ( .A(G160), .B(G162), .ZN(n883) );
  XNOR2_X1 U987 ( .A(n884), .B(n883), .ZN(n901) );
  NAND2_X1 U988 ( .A1(G115), .A2(n885), .ZN(n888) );
  NAND2_X1 U989 ( .A1(G127), .A2(n886), .ZN(n887) );
  NAND2_X1 U990 ( .A1(n888), .A2(n887), .ZN(n889) );
  XNOR2_X1 U991 ( .A(n889), .B(KEYINPUT47), .ZN(n892) );
  NAND2_X1 U992 ( .A1(G103), .A2(n890), .ZN(n891) );
  NAND2_X1 U993 ( .A1(n892), .A2(n891), .ZN(n896) );
  NAND2_X1 U994 ( .A1(n893), .A2(G139), .ZN(n894) );
  XOR2_X1 U995 ( .A(KEYINPUT114), .B(n894), .Z(n895) );
  NOR2_X1 U996 ( .A1(n896), .A2(n895), .ZN(n927) );
  XNOR2_X1 U997 ( .A(n927), .B(n897), .ZN(n899) );
  XNOR2_X1 U998 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U999 ( .A(n901), .B(n900), .Z(n906) );
  XOR2_X1 U1000 ( .A(KEYINPUT113), .B(KEYINPUT46), .Z(n903) );
  XNOR2_X1 U1001 ( .A(KEYINPUT48), .B(KEYINPUT115), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(G164), .B(n904), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1005 ( .A(n908), .B(n907), .Z(n909) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n909), .ZN(G395) );
  XNOR2_X1 U1007 ( .A(KEYINPUT117), .B(KEYINPUT116), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(n983), .B(n910), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1010 ( .A(G171), .B(n913), .Z(n914) );
  XNOR2_X1 U1011 ( .A(n989), .B(n914), .ZN(n915) );
  XOR2_X1 U1012 ( .A(G286), .B(n915), .Z(n916) );
  NOR2_X1 U1013 ( .A1(G37), .A2(n916), .ZN(G397) );
  NOR2_X1 U1014 ( .A1(G227), .A2(G229), .ZN(n917) );
  XOR2_X1 U1015 ( .A(KEYINPUT49), .B(n917), .Z(n918) );
  NAND2_X1 U1016 ( .A1(n918), .A2(G319), .ZN(n919) );
  NOR2_X1 U1017 ( .A1(G401), .A2(n919), .ZN(n920) );
  XNOR2_X1 U1018 ( .A(KEYINPUT118), .B(n920), .ZN(n922) );
  NOR2_X1 U1019 ( .A1(G395), .A2(G397), .ZN(n921) );
  NAND2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n923) );
  XOR2_X1 U1021 ( .A(KEYINPUT119), .B(n923), .Z(G225) );
  INV_X1 U1022 ( .A(G225), .ZN(G308) );
  INV_X1 U1023 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n936) );
  XNOR2_X1 U1025 ( .A(G164), .B(G2078), .ZN(n926) );
  XNOR2_X1 U1026 ( .A(n926), .B(KEYINPUT121), .ZN(n929) );
  XOR2_X1 U1027 ( .A(G2072), .B(n927), .Z(n928) );
  NOR2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1029 ( .A(KEYINPUT50), .B(n930), .ZN(n932) );
  XNOR2_X1 U1030 ( .A(G160), .B(G2084), .ZN(n931) );
  NAND2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n942) );
  XNOR2_X1 U1034 ( .A(G162), .B(G2090), .ZN(n938) );
  NAND2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1036 ( .A(KEYINPUT120), .B(n939), .Z(n940) );
  XNOR2_X1 U1037 ( .A(KEYINPUT51), .B(n940), .ZN(n941) );
  NOR2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n944) );
  NAND2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1040 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1041 ( .A(KEYINPUT52), .B(n947), .ZN(n948) );
  XOR2_X1 U1042 ( .A(KEYINPUT55), .B(KEYINPUT122), .Z(n968) );
  NAND2_X1 U1043 ( .A1(n948), .A2(n968), .ZN(n949) );
  NAND2_X1 U1044 ( .A1(n949), .A2(G29), .ZN(n1026) );
  XNOR2_X1 U1045 ( .A(G2090), .B(G35), .ZN(n963) );
  XNOR2_X1 U1046 ( .A(G2067), .B(G26), .ZN(n951) );
  XNOR2_X1 U1047 ( .A(G1996), .B(G32), .ZN(n950) );
  NOR2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n956) );
  XOR2_X1 U1049 ( .A(n952), .B(G27), .Z(n954) );
  XNOR2_X1 U1050 ( .A(G33), .B(G2072), .ZN(n953) );
  NOR2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1053 ( .A(KEYINPUT123), .B(n957), .ZN(n958) );
  NAND2_X1 U1054 ( .A1(n958), .A2(G28), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(G25), .B(G1991), .ZN(n959) );
  NOR2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1057 ( .A(KEYINPUT53), .B(n961), .ZN(n962) );
  NOR2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n966) );
  XOR2_X1 U1059 ( .A(G2084), .B(G34), .Z(n964) );
  XNOR2_X1 U1060 ( .A(KEYINPUT54), .B(n964), .ZN(n965) );
  NAND2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1062 ( .A(n968), .B(n967), .ZN(n970) );
  INV_X1 U1063 ( .A(G29), .ZN(n969) );
  NAND2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1065 ( .A1(G11), .A2(n971), .ZN(n1024) );
  XNOR2_X1 U1066 ( .A(G16), .B(KEYINPUT56), .ZN(n995) );
  XNOR2_X1 U1067 ( .A(G1966), .B(G168), .ZN(n973) );
  NAND2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(n974), .B(KEYINPUT57), .ZN(n993) );
  NAND2_X1 U1070 ( .A1(G1971), .A2(G303), .ZN(n975) );
  NAND2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n978) );
  XNOR2_X1 U1072 ( .A(G1956), .B(G299), .ZN(n977) );
  NOR2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n987) );
  XOR2_X1 U1076 ( .A(G171), .B(G1961), .Z(n985) );
  XNOR2_X1 U1077 ( .A(n983), .B(G1348), .ZN(n984) );
  NOR2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1080 ( .A(KEYINPUT124), .B(n988), .ZN(n991) );
  XNOR2_X1 U1081 ( .A(G1341), .B(n989), .ZN(n990) );
  NOR2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n1022) );
  INV_X1 U1085 ( .A(G16), .ZN(n1020) );
  XNOR2_X1 U1086 ( .A(G5), .B(n996), .ZN(n1010) );
  XNOR2_X1 U1087 ( .A(G1956), .B(G20), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(KEYINPUT59), .B(KEYINPUT125), .ZN(n997) );
  XNOR2_X1 U1089 ( .A(n997), .B(G4), .ZN(n998) );
  XNOR2_X1 U1090 ( .A(n998), .B(G1348), .ZN(n999) );
  NOR2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1004) );
  XNOR2_X1 U1092 ( .A(G1341), .B(G19), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(G1981), .B(G6), .ZN(n1001) );
  NOR2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1096 ( .A(n1005), .B(KEYINPUT60), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(KEYINPUT126), .B(G1966), .ZN(n1006) );
  XNOR2_X1 U1098 ( .A(G21), .B(n1006), .ZN(n1007) );
  NOR2_X1 U1099 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1017) );
  XNOR2_X1 U1101 ( .A(G1971), .B(G22), .ZN(n1012) );
  XNOR2_X1 U1102 ( .A(G23), .B(G1976), .ZN(n1011) );
  NOR2_X1 U1103 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  XOR2_X1 U1104 ( .A(G1986), .B(G24), .Z(n1013) );
  NAND2_X1 U1105 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1106 ( .A(KEYINPUT58), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1108 ( .A(KEYINPUT61), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1109 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1113 ( .A(n1027), .B(KEYINPUT62), .ZN(n1028) );
  XNOR2_X1 U1114 ( .A(KEYINPUT127), .B(n1028), .ZN(G311) );
  INV_X1 U1115 ( .A(G311), .ZN(G150) );
endmodule

