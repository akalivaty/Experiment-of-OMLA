//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 1 0 1 1 1 0 1 0 0 0 0 0 0 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1275, new_n1276, new_n1277, new_n1279,
    new_n1280, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G77), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(G355));
  NOR2_X1   g0006(.A1(G58), .A2(G68), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G50), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(G13), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT0), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT65), .Z(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n215), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n214), .B(new_n218), .C1(new_n225), .C2(KEYINPUT1), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G250), .B(G257), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT66), .ZN(new_n229));
  XOR2_X1   g0029(.A(G264), .B(G270), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n231), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT67), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  NAND3_X1  g0045(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(new_n211), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n202), .A2(G20), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT8), .B(G58), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(G20), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  AOI22_X1  g0054(.A1(new_n251), .A2(new_n253), .B1(G150), .B2(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n248), .B1(new_n249), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G13), .A3(G20), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(new_n247), .ZN(new_n260));
  OR3_X1    g0060(.A1(new_n212), .A2(KEYINPUT69), .A3(G1), .ZN(new_n261));
  OAI21_X1  g0061(.A(KEYINPUT69), .B1(new_n212), .B2(G1), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n260), .A2(new_n263), .A3(G50), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n264), .B1(G50), .B2(new_n258), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n256), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT3), .B(G33), .ZN(new_n267));
  INV_X1    g0067(.A(G1698), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(G222), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G77), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n267), .A2(G1698), .ZN(new_n271));
  INV_X1    g0071(.A(G223), .ZN(new_n272));
  OAI221_X1 g0072(.A(new_n269), .B1(new_n270), .B2(new_n267), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G33), .A2(G41), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(G1), .A3(G13), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  AND2_X1   g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  OAI21_X1  g0078(.A(G274), .B1(new_n278), .B2(new_n211), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n257), .B1(G41), .B2(G45), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT68), .ZN(new_n281));
  INV_X1    g0081(.A(G41), .ZN(new_n282));
  INV_X1    g0082(.A(G45), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT68), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n284), .A2(new_n285), .A3(new_n257), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n279), .B1(new_n281), .B2(new_n286), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n275), .A2(new_n280), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n287), .B1(G226), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n277), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G169), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n266), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n290), .ZN(new_n293));
  INV_X1    g0093(.A(G179), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n266), .A2(KEYINPUT9), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT70), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n297), .B(new_n298), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n293), .A2(G190), .B1(new_n266), .B2(KEYINPUT9), .ZN(new_n300));
  INV_X1    g0100(.A(G200), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n301), .B1(new_n277), .B2(new_n289), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT71), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n303), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n300), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NOR3_X1   g0106(.A1(new_n299), .A2(new_n306), .A3(KEYINPUT10), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT10), .ZN(new_n308));
  AND3_X1   g0108(.A1(new_n300), .A2(new_n304), .A3(new_n305), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n297), .B(KEYINPUT70), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n296), .B1(new_n307), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G68), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n259), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n314), .B(KEYINPUT12), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n254), .A2(G50), .B1(G20), .B2(new_n313), .ZN(new_n316));
  INV_X1    g0116(.A(new_n253), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n316), .B1(new_n317), .B2(new_n270), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n318), .A2(KEYINPUT11), .A3(new_n247), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n260), .A2(new_n263), .A3(G68), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n315), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT11), .B1(new_n318), .B2(new_n247), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(G33), .A2(G97), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n267), .A2(new_n268), .ZN(new_n326));
  INV_X1    g0126(.A(G226), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT3), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G33), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NOR3_X1   g0132(.A1(new_n332), .A2(new_n233), .A3(new_n268), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n276), .B1(new_n328), .B2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n287), .B1(G238), .B2(new_n288), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT13), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT13), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n334), .A2(new_n335), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT72), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT14), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n340), .A2(G169), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n337), .A2(G179), .A3(new_n339), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n342), .B1(new_n340), .B2(G169), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n324), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n340), .A2(G200), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n337), .A2(G190), .A3(new_n339), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(new_n323), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n270), .B1(new_n261), .B2(new_n262), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n352), .A2(new_n260), .B1(new_n270), .B2(new_n259), .ZN(new_n353));
  INV_X1    g0153(.A(new_n254), .ZN(new_n354));
  OAI22_X1  g0154(.A1(new_n250), .A2(new_n354), .B1(new_n212), .B2(new_n270), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT15), .B(G87), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n356), .A2(new_n317), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n247), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(G238), .ZN(new_n361));
  INV_X1    g0161(.A(G107), .ZN(new_n362));
  OAI22_X1  g0162(.A1(new_n271), .A2(new_n361), .B1(new_n362), .B2(new_n267), .ZN(new_n363));
  NOR3_X1   g0163(.A1(new_n332), .A2(new_n233), .A3(G1698), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n276), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n287), .B1(G244), .B2(new_n288), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n360), .B1(new_n291), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(G179), .B2(new_n367), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n359), .B1(new_n367), .B2(G200), .ZN(new_n370));
  INV_X1    g0170(.A(G190), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n370), .B1(new_n371), .B2(new_n367), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  NOR3_X1   g0173(.A1(new_n312), .A2(new_n351), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT16), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT7), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n376), .B1(new_n267), .B2(G20), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n332), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n313), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G58), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n380), .A2(new_n313), .ZN(new_n381));
  OAI21_X1  g0181(.A(G20), .B1(new_n381), .B2(new_n207), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n254), .A2(G159), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n375), .B1(new_n379), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT74), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n384), .ZN(new_n388));
  NOR3_X1   g0188(.A1(new_n267), .A2(new_n376), .A3(G20), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT73), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n330), .A2(G33), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n329), .A2(new_n331), .A3(KEYINPUT73), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n393), .A2(new_n212), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n389), .B1(new_n395), .B2(new_n376), .ZN(new_n396));
  OAI211_X1 g0196(.A(KEYINPUT16), .B(new_n388), .C1(new_n396), .C2(new_n313), .ZN(new_n397));
  OAI211_X1 g0197(.A(KEYINPUT74), .B(new_n375), .C1(new_n379), .C2(new_n384), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n387), .A2(new_n397), .A3(new_n247), .A4(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n275), .A2(G232), .A3(new_n280), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT75), .B1(new_n287), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(G274), .ZN(new_n403));
  AND2_X1   g0203(.A1(G1), .A2(G13), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n403), .B1(new_n404), .B2(new_n274), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n285), .B1(new_n284), .B2(new_n257), .ZN(new_n406));
  NOR2_X1   g0206(.A1(G41), .A2(G45), .ZN(new_n407));
  NOR3_X1   g0207(.A1(new_n407), .A2(KEYINPUT68), .A3(G1), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n405), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT75), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n409), .A2(new_n410), .A3(new_n400), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n329), .A2(new_n331), .A3(G226), .A4(G1698), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n329), .A2(new_n331), .A3(G223), .A4(new_n268), .ZN(new_n413));
  INV_X1    g0213(.A(G87), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n412), .B(new_n413), .C1(new_n252), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n276), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n402), .A2(new_n411), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n301), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n402), .A2(new_n411), .A3(new_n416), .A4(new_n371), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n263), .A2(new_n251), .ZN(new_n421));
  INV_X1    g0221(.A(new_n260), .ZN(new_n422));
  OAI22_X1  g0222(.A1(new_n421), .A2(new_n422), .B1(new_n258), .B2(new_n251), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n399), .A2(new_n420), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT17), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n399), .A2(new_n420), .A3(KEYINPUT17), .A4(new_n424), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n399), .A2(new_n424), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n417), .A2(G169), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n402), .A2(new_n411), .A3(new_n416), .A4(G179), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT76), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT76), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n431), .A2(new_n435), .A3(new_n432), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n430), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT18), .ZN(new_n438));
  AND3_X1   g0238(.A1(new_n431), .A2(new_n435), .A3(new_n432), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n435), .B1(new_n431), .B2(new_n432), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT18), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n441), .A2(new_n442), .A3(new_n430), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n429), .A2(new_n438), .A3(new_n443), .ZN(new_n444));
  OR2_X1    g0244(.A1(new_n444), .A2(KEYINPUT77), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(KEYINPUT77), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n374), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT78), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n448), .B1(new_n282), .B2(KEYINPUT5), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT5), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n449), .B1(new_n450), .B2(G41), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n257), .A2(G45), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n450), .A2(G41), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n452), .B1(new_n453), .B2(new_n448), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n276), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n455), .A2(KEYINPUT84), .A3(G264), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n283), .A2(G1), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n448), .A2(new_n282), .A3(KEYINPUT5), .ZN(new_n458));
  AOI21_X1  g0258(.A(KEYINPUT78), .B1(new_n450), .B2(G41), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n457), .B(new_n458), .C1(new_n459), .C2(new_n453), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n460), .A2(G264), .A3(new_n275), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT84), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n267), .A2(G257), .A3(G1698), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G294), .ZN(new_n465));
  INV_X1    g0265(.A(G250), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n464), .B(new_n465), .C1(new_n326), .C2(new_n466), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n456), .A2(new_n463), .B1(new_n276), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n451), .A2(new_n454), .A3(new_n405), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n468), .A2(new_n294), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n467), .A2(new_n276), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT84), .B1(new_n455), .B2(G264), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n461), .A2(new_n462), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n469), .B(new_n471), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n291), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n267), .A2(new_n212), .A3(G87), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT22), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT22), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n267), .A2(new_n478), .A3(new_n212), .A4(G87), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT23), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n481), .A2(new_n362), .A3(G20), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT83), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n484), .B1(new_n481), .B2(new_n362), .ZN(new_n485));
  AOI21_X1  g0285(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n486));
  OAI22_X1  g0286(.A1(new_n482), .A2(new_n483), .B1(new_n486), .B2(G20), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n480), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT24), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT24), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n480), .A2(new_n491), .A3(new_n488), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n248), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(KEYINPUT25), .B1(new_n259), .B2(new_n362), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n259), .A2(KEYINPUT25), .A3(new_n362), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n257), .A2(G33), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n258), .A2(new_n497), .A3(new_n211), .A4(new_n246), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n495), .A2(new_n496), .B1(G107), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n470), .B(new_n475), .C1(new_n493), .C2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n474), .A2(G200), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n480), .A2(new_n491), .A3(new_n488), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n491), .B1(new_n480), .B2(new_n488), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n247), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n468), .A2(G190), .A3(new_n469), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n503), .A2(new_n506), .A3(new_n507), .A4(new_n500), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n502), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n460), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n455), .A2(G257), .B1(new_n510), .B2(new_n405), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G33), .A2(G283), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n329), .A2(new_n331), .A3(G250), .A4(G1698), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n329), .A2(new_n331), .A3(G244), .A4(new_n268), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT4), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n512), .B(new_n513), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n514), .A2(new_n515), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n276), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n511), .A2(new_n518), .A3(G179), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n291), .B1(new_n511), .B2(new_n518), .ZN(new_n520));
  AOI21_X1  g0320(.A(KEYINPUT7), .B1(new_n332), .B2(new_n212), .ZN(new_n521));
  OAI21_X1  g0321(.A(G107), .B1(new_n389), .B2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT6), .ZN(new_n523));
  AND2_X1   g0323(.A1(G97), .A2(G107), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n523), .B1(new_n524), .B2(new_n204), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n362), .A2(KEYINPUT6), .A3(G97), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n527), .A2(G20), .B1(G77), .B2(new_n254), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n248), .B1(new_n522), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n258), .A2(G97), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n530), .B1(new_n499), .B2(G97), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  OAI22_X1  g0332(.A1(new_n519), .A2(new_n520), .B1(new_n529), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n511), .A2(new_n518), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G200), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n522), .A2(new_n528), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n532), .B1(new_n536), .B2(new_n247), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n535), .B(new_n537), .C1(new_n371), .C2(new_n534), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n361), .A2(new_n268), .ZN(new_n539));
  INV_X1    g0339(.A(G244), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(G1698), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n329), .A2(new_n539), .A3(new_n331), .A4(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(G116), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n252), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n275), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n466), .B1(new_n257), .B2(G45), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n275), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n279), .B2(new_n452), .ZN(new_n549));
  OAI21_X1  g0349(.A(KEYINPUT79), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n405), .A2(new_n457), .B1(new_n275), .B2(new_n547), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT79), .ZN(new_n552));
  NOR2_X1   g0352(.A1(G238), .A2(G1698), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n553), .B1(new_n540), .B2(G1698), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n544), .B1(new_n554), .B2(new_n267), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n551), .B(new_n552), .C1(new_n555), .C2(new_n275), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n550), .A2(new_n556), .A3(new_n294), .ZN(new_n557));
  INV_X1    g0357(.A(new_n356), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n558), .A2(new_n258), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n267), .A2(new_n212), .A3(G68), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT19), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n212), .B1(new_n325), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(G87), .B2(new_n205), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n212), .A2(G33), .A3(G97), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT80), .ZN(new_n565));
  AND3_X1   g0365(.A1(new_n564), .A2(new_n565), .A3(new_n561), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n565), .B1(new_n564), .B2(new_n561), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n560), .B(new_n563), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n559), .B1(new_n568), .B2(new_n247), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n499), .A2(new_n558), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n550), .A2(new_n556), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n557), .B(new_n571), .C1(new_n572), .C2(G169), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n550), .A2(new_n556), .A3(G190), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n498), .A2(new_n414), .ZN(new_n575));
  AOI211_X1 g0375(.A(new_n559), .B(new_n575), .C1(new_n568), .C2(new_n247), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n574), .B(new_n576), .C1(new_n572), .C2(new_n301), .ZN(new_n577));
  AND4_X1   g0377(.A1(new_n533), .A2(new_n538), .A3(new_n573), .A4(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(G97), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n512), .B(new_n212), .C1(G33), .C2(new_n579), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n580), .B(new_n247), .C1(new_n212), .C2(G116), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT20), .ZN(new_n582));
  XNOR2_X1  g0382(.A(new_n581), .B(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n258), .A2(G116), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n584), .B1(new_n499), .B2(G116), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n291), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT81), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n460), .A2(G270), .A3(new_n275), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n588), .B1(new_n589), .B2(new_n469), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n588), .A3(new_n469), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n329), .A2(new_n331), .A3(G264), .A4(G1698), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n329), .A2(new_n331), .A3(G257), .A4(new_n268), .ZN(new_n594));
  INV_X1    g0394(.A(G303), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n593), .B(new_n594), .C1(new_n595), .C2(new_n267), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n276), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(KEYINPUT82), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT82), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n596), .A2(new_n599), .A3(new_n276), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n591), .A2(new_n592), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(KEYINPUT21), .B1(new_n587), .B2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n592), .ZN(new_n603));
  INV_X1    g0403(.A(new_n600), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n599), .B1(new_n596), .B2(new_n276), .ZN(new_n605));
  OAI22_X1  g0405(.A1(new_n603), .A2(new_n590), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT21), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n606), .A2(new_n607), .A3(new_n586), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n583), .A2(new_n585), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n610), .A2(new_n294), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n602), .A2(new_n608), .B1(new_n601), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n606), .A2(G200), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n613), .B(new_n610), .C1(new_n371), .C2(new_n606), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n509), .A2(new_n578), .A3(new_n612), .A4(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n447), .A2(new_n615), .ZN(G372));
  INV_X1    g0416(.A(new_n296), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n430), .A2(new_n433), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(KEYINPUT18), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n399), .A2(new_n424), .B1(new_n431), .B2(new_n432), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n442), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g0422(.A(new_n369), .B(KEYINPUT88), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n346), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n625), .A2(new_n344), .A3(new_n343), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n624), .A2(new_n350), .B1(new_n324), .B2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n429), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n622), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT89), .ZN(new_n630));
  OR2_X1    g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(KEYINPUT10), .B1(new_n299), .B2(new_n306), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n309), .A2(new_n310), .A3(new_n308), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n629), .A2(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n617), .B1(new_n631), .B2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT85), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n546), .A2(new_n549), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n636), .B1(new_n637), .B2(new_n301), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n551), .B1(new_n555), .B2(new_n275), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n639), .A2(KEYINPUT85), .A3(G200), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n576), .A2(new_n574), .A3(new_n638), .A4(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n639), .A2(new_n291), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n571), .A2(new_n557), .A3(new_n642), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n644), .A2(new_n508), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n538), .A2(new_n533), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(KEYINPUT86), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT86), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n645), .A2(new_n649), .A3(new_n646), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n611), .A2(new_n601), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n607), .B1(new_n606), .B2(new_n586), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n606), .A2(new_n586), .A3(new_n607), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n502), .B(new_n651), .C1(new_n652), .C2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n648), .A2(new_n650), .A3(new_n654), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n573), .A2(new_n577), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n534), .A2(G169), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n511), .A2(new_n518), .A3(G179), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n537), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n656), .A2(KEYINPUT26), .A3(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT26), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n641), .A2(new_n643), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n661), .B1(new_n662), .B2(new_n533), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n660), .A2(KEYINPUT87), .A3(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n643), .B1(new_n660), .B2(KEYINPUT87), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n655), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n635), .B1(new_n447), .B2(new_n667), .ZN(G369));
  NAND2_X1  g0468(.A1(new_n602), .A2(new_n608), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n651), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n257), .A2(new_n212), .A3(G13), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(G213), .A3(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(G343), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n610), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n670), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n669), .A2(new_n614), .A3(new_n651), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n679), .B1(new_n680), .B2(new_n678), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(G330), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n676), .B1(new_n493), .B2(new_n501), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n509), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n502), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n676), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n683), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n612), .A2(new_n676), .ZN(new_n690));
  XOR2_X1   g0490(.A(new_n676), .B(KEYINPUT90), .Z(new_n691));
  AOI22_X1  g0491(.A1(new_n690), .A2(new_n509), .B1(new_n686), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n689), .A2(new_n692), .ZN(G399));
  NOR3_X1   g0493(.A1(new_n205), .A2(G87), .A3(G116), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n216), .A2(new_n282), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(new_n695), .A3(G1), .ZN(new_n696));
  OAI22_X1  g0496(.A1(new_n696), .A2(KEYINPUT91), .B1(new_n209), .B2(new_n695), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n697), .B1(KEYINPUT91), .B2(new_n696), .ZN(new_n698));
  XOR2_X1   g0498(.A(new_n698), .B(KEYINPUT28), .Z(new_n699));
  INV_X1    g0499(.A(KEYINPUT94), .ZN(new_n700));
  INV_X1    g0500(.A(G330), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n656), .A2(new_n533), .A3(new_n538), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n502), .A2(new_n508), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n680), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT93), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(new_n705), .A3(new_n691), .ZN(new_n706));
  INV_X1    g0506(.A(new_n691), .ZN(new_n707));
  OAI21_X1  g0507(.A(KEYINPUT93), .B1(new_n615), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n707), .A2(KEYINPUT31), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n550), .A2(new_n556), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n713), .A2(KEYINPUT30), .A3(new_n601), .A4(new_n519), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n637), .A2(G179), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n606), .A2(new_n474), .A3(new_n534), .A4(new_n715), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT30), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n519), .A2(new_n468), .A3(new_n572), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n718), .B1(new_n719), .B2(new_n606), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n710), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT92), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  OAI211_X1 g0523(.A(KEYINPUT92), .B(new_n718), .C1(new_n719), .C2(new_n606), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n717), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n676), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT31), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n721), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  AOI211_X1 g0528(.A(new_n700), .B(new_n701), .C1(new_n709), .C2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n705), .B1(new_n704), .B2(new_n691), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n615), .A2(KEYINPUT93), .A3(new_n707), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n728), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(KEYINPUT94), .B1(new_n732), .B2(G330), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(KEYINPUT26), .B1(new_n662), .B2(new_n533), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n659), .A2(new_n661), .A3(new_n573), .A4(new_n577), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n735), .A2(new_n643), .A3(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT95), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n654), .A2(new_n645), .A3(new_n646), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n735), .A2(new_n736), .A3(KEYINPUT95), .A4(new_n643), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n739), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n742), .A2(KEYINPUT96), .A3(new_n677), .ZN(new_n743));
  AOI21_X1  g0543(.A(KEYINPUT96), .B1(new_n742), .B2(new_n677), .ZN(new_n744));
  OAI21_X1  g0544(.A(KEYINPUT29), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n707), .B1(new_n655), .B2(new_n666), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n745), .B1(KEYINPUT29), .B2(new_n746), .ZN(new_n747));
  AND2_X1   g0547(.A1(new_n734), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n699), .B1(new_n748), .B2(G1), .ZN(G364));
  AND2_X1   g0549(.A1(new_n212), .A2(G13), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n257), .B1(new_n750), .B2(G45), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n695), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n683), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(G330), .B2(new_n681), .ZN(new_n756));
  INV_X1    g0556(.A(G355), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n267), .A2(new_n216), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n757), .A2(new_n758), .B1(G116), .B2(new_n216), .ZN(new_n759));
  AND2_X1   g0559(.A1(new_n393), .A2(new_n394), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(new_n216), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n761), .B1(new_n283), .B2(new_n210), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n244), .A2(G45), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n759), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G13), .A2(G33), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n211), .B1(G20), .B2(new_n291), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n754), .B1(new_n764), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n212), .A2(G179), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n772), .A2(new_n371), .A3(G200), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n773), .B(KEYINPUT99), .Z(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G107), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n371), .A2(new_n301), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(new_n772), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n267), .B1(new_n777), .B2(new_n414), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(KEYINPUT98), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n778), .A2(KEYINPUT98), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n775), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT100), .Z(new_n782));
  NOR2_X1   g0582(.A1(new_n212), .A2(new_n294), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n784), .A2(new_n371), .A3(G200), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n776), .A2(new_n783), .ZN(new_n787));
  INV_X1    g0587(.A(G50), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n786), .A2(new_n380), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NOR3_X1   g0589(.A1(new_n784), .A2(new_n301), .A3(G190), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G190), .A2(G200), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n783), .A2(new_n792), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n791), .A2(new_n313), .B1(new_n793), .B2(new_n270), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n789), .A2(new_n794), .ZN(new_n795));
  NOR3_X1   g0595(.A1(new_n371), .A2(G179), .A3(G200), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n212), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G97), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n772), .A2(new_n792), .ZN(new_n800));
  XNOR2_X1  g0600(.A(KEYINPUT97), .B(G159), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT32), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n795), .A2(new_n799), .A3(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n332), .B1(new_n777), .B2(new_n595), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT101), .ZN(new_n806));
  INV_X1    g0606(.A(new_n793), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G311), .ZN(new_n808));
  INV_X1    g0608(.A(G322), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n808), .B1(new_n786), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(G294), .B2(new_n798), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n774), .A2(G283), .ZN(new_n812));
  XNOR2_X1  g0612(.A(KEYINPUT33), .B(G317), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n790), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n787), .ZN(new_n815));
  INV_X1    g0615(.A(new_n800), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n815), .A2(G326), .B1(new_n816), .B2(G329), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n811), .A2(new_n812), .A3(new_n814), .A4(new_n817), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n782), .A2(new_n804), .B1(new_n806), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n771), .B1(new_n819), .B2(new_n768), .ZN(new_n820));
  INV_X1    g0620(.A(new_n767), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n820), .B1(new_n681), .B2(new_n821), .ZN(new_n822));
  AND2_X1   g0622(.A1(new_n756), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(G396));
  INV_X1    g0624(.A(new_n734), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n360), .A2(new_n677), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n369), .A2(new_n372), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n623), .B2(new_n827), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n746), .B(new_n830), .ZN(new_n831));
  OR2_X1    g0631(.A1(new_n825), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n754), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n825), .A2(new_n831), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n768), .A2(new_n765), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n754), .B1(G77), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(G294), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n786), .A2(new_n839), .B1(new_n793), .B2(new_n543), .ZN(new_n840));
  INV_X1    g0640(.A(new_n777), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n267), .B(new_n840), .C1(G107), .C2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n774), .A2(G87), .ZN(new_n843));
  INV_X1    g0643(.A(G283), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n791), .A2(new_n844), .B1(new_n787), .B2(new_n595), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(G311), .B2(new_n816), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n842), .A2(new_n799), .A3(new_n843), .A4(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(G137), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n787), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(G143), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n786), .A2(new_n850), .B1(new_n793), .B2(new_n801), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n849), .B(new_n851), .C1(G150), .C2(new_n790), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n852), .A2(KEYINPUT34), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT102), .ZN(new_n854));
  INV_X1    g0654(.A(new_n760), .ZN(new_n855));
  INV_X1    g0655(.A(G132), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n855), .B1(new_n856), .B2(new_n800), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n853), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n854), .B2(new_n857), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n852), .A2(KEYINPUT34), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n774), .A2(G68), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n798), .A2(G58), .B1(new_n841), .B2(G50), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n847), .B1(new_n859), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n838), .B1(new_n864), .B2(new_n768), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n829), .B2(new_n766), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n835), .A2(new_n866), .ZN(G384));
  OR2_X1    g0667(.A1(new_n527), .A2(KEYINPUT35), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n527), .A2(KEYINPUT35), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n868), .A2(G116), .A3(new_n213), .A4(new_n869), .ZN(new_n870));
  XOR2_X1   g0670(.A(new_n870), .B(KEYINPUT36), .Z(new_n871));
  OR3_X1    g0671(.A1(new_n209), .A2(new_n270), .A3(new_n381), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n788), .A2(G68), .ZN(new_n873));
  AOI211_X1 g0673(.A(new_n257), .B(G13), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n397), .A2(new_n247), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n388), .B1(new_n396), .B2(new_n313), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n375), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n423), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n879), .A2(new_n674), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n444), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n433), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n425), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT37), .B1(new_n883), .B2(new_n880), .ZN(new_n884));
  INV_X1    g0684(.A(new_n674), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n430), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT37), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n437), .A2(new_n886), .A3(new_n887), .A4(new_n425), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n881), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT38), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n881), .A2(new_n889), .A3(KEYINPUT38), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n350), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n324), .B(new_n676), .C1(new_n626), .C2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n324), .A2(new_n676), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n347), .A2(new_n350), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n829), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n726), .B(KEYINPUT31), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n900), .B1(new_n901), .B2(new_n709), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT40), .B1(new_n894), .B2(new_n902), .ZN(new_n903));
  AND3_X1   g0703(.A1(new_n399), .A2(new_n424), .A3(new_n420), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n674), .B1(new_n399), .B2(new_n424), .ZN(new_n905));
  NOR3_X1   g0705(.A1(new_n904), .A2(new_n620), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n888), .B1(new_n906), .B2(new_n887), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT103), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n619), .A2(new_n427), .A3(new_n428), .A4(new_n621), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n907), .A2(new_n908), .B1(new_n905), .B2(new_n909), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n888), .B(KEYINPUT103), .C1(new_n906), .C2(new_n887), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n891), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT104), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n881), .A2(new_n889), .A3(KEYINPUT38), .ZN(new_n916));
  AOI21_X1  g0716(.A(KEYINPUT38), .B1(new_n910), .B2(new_n911), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n916), .B1(new_n917), .B2(KEYINPUT104), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n901), .A2(new_n709), .ZN(new_n920));
  INV_X1    g0720(.A(new_n900), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT40), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n903), .B1(new_n919), .B2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n447), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n925), .A2(new_n926), .A3(new_n920), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n925), .B1(new_n926), .B2(new_n920), .ZN(new_n928));
  OR3_X1    g0728(.A1(new_n927), .A2(new_n928), .A3(new_n701), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n892), .A2(new_n893), .ZN(new_n930));
  INV_X1    g0730(.A(new_n899), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n369), .A2(new_n676), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n746), .B2(new_n829), .ZN(new_n933));
  NOR3_X1   g0733(.A1(new_n930), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n622), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n934), .B1(new_n935), .B2(new_n674), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT39), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n909), .A2(new_n905), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n618), .A2(new_n886), .A3(new_n425), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n905), .B1(new_n441), .B2(new_n430), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n904), .A2(KEYINPUT37), .ZN(new_n941));
  AOI22_X1  g0741(.A1(KEYINPUT37), .A2(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n938), .B1(new_n942), .B2(KEYINPUT103), .ZN(new_n943));
  INV_X1    g0743(.A(new_n911), .ZN(new_n944));
  OAI211_X1 g0744(.A(KEYINPUT104), .B(new_n891), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n893), .ZN(new_n946));
  AOI21_X1  g0746(.A(KEYINPUT104), .B1(new_n912), .B2(new_n891), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n937), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n626), .A2(new_n324), .A3(new_n677), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n930), .A2(KEYINPUT39), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n948), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n936), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n635), .B1(new_n747), .B2(new_n447), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n953), .B(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n929), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n257), .B2(new_n750), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n929), .A2(new_n955), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n875), .B1(new_n957), .B2(new_n958), .ZN(G367));
  AND3_X1   g0759(.A1(new_n231), .A2(new_n216), .A3(new_n760), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n769), .B1(new_n216), .B2(new_n356), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n754), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(G150), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n786), .A2(new_n963), .B1(new_n800), .B2(new_n848), .ZN(new_n964));
  INV_X1    g0764(.A(new_n773), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n332), .B(new_n964), .C1(G77), .C2(new_n965), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n791), .A2(new_n801), .B1(new_n793), .B2(new_n788), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n787), .A2(new_n850), .B1(new_n777), .B2(new_n380), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n966), .B(new_n969), .C1(new_n313), .C2(new_n797), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n785), .A2(G303), .B1(G283), .B2(new_n807), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n971), .B(new_n760), .C1(new_n362), .C2(new_n797), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n841), .A2(G116), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT46), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n790), .A2(G294), .B1(G97), .B2(new_n965), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n815), .A2(G311), .B1(new_n816), .B2(G317), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n974), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n970), .B1(new_n972), .B2(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT47), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n962), .B1(new_n979), .B2(new_n768), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n576), .A2(new_n677), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n981), .A2(new_n557), .A3(new_n571), .A4(new_n642), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n662), .B2(new_n981), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n983), .A2(new_n821), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n980), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n670), .A2(new_n509), .A3(new_n677), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n538), .B(new_n533), .C1(new_n537), .C2(new_n691), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n659), .A2(new_n707), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n686), .A2(new_n691), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n986), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT45), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n991), .B(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT44), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n692), .B2(new_n989), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n986), .A2(new_n990), .ZN(new_n996));
  INV_X1    g0796(.A(new_n989), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n996), .A2(KEYINPUT44), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n993), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n689), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n993), .A2(new_n689), .A3(new_n999), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n986), .B1(new_n688), .B2(new_n690), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(new_n682), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n747), .B(new_n734), .C1(new_n1004), .C2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n695), .B(KEYINPUT41), .Z(new_n1008));
  AND3_X1   g0808(.A1(new_n1007), .A2(KEYINPUT106), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(KEYINPUT106), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1010));
  NOR3_X1   g0810(.A1(new_n1009), .A2(new_n1010), .A3(new_n752), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT107), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n986), .A2(new_n997), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT42), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n533), .B1(new_n987), .B2(new_n502), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n691), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  OR3_X1    g0817(.A1(new_n1017), .A2(KEYINPUT43), .A3(new_n983), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n983), .B(KEYINPUT43), .Z(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(KEYINPUT105), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT105), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1017), .A2(new_n1022), .A3(new_n1019), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1018), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n689), .B2(new_n997), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n689), .A2(new_n997), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1018), .A2(new_n1021), .A3(new_n1026), .A4(new_n1023), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  NOR3_X1   g0828(.A1(new_n1011), .A2(new_n1012), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT106), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n752), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1007), .A2(KEYINPUT106), .A3(new_n1008), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1028), .ZN(new_n1035));
  AOI21_X1  g0835(.A(KEYINPUT107), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n985), .B1(new_n1029), .B2(new_n1036), .ZN(G387));
  INV_X1    g0837(.A(new_n1006), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n685), .A2(new_n687), .A3(new_n767), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n694), .A2(new_n758), .B1(G107), .B2(new_n216), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n694), .ZN(new_n1041));
  AOI211_X1 g0841(.A(G45), .B(new_n1041), .C1(G68), .C2(G77), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n250), .A2(G50), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT50), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n761), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n236), .A2(G45), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1040), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n754), .B1(new_n1047), .B2(new_n770), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(G68), .A2(new_n807), .B1(new_n816), .B2(G150), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n841), .A2(G77), .ZN(new_n1050));
  INV_X1    g0850(.A(G159), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1049), .B(new_n1050), .C1(new_n1051), .C2(new_n787), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(G97), .B2(new_n774), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n788), .A2(new_n786), .B1(new_n791), .B2(new_n250), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n797), .A2(new_n356), .ZN(new_n1055));
  NOR3_X1   g0855(.A1(new_n1054), .A2(new_n760), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1053), .A2(new_n1056), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n965), .A2(G116), .B1(new_n816), .B2(G326), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n797), .A2(new_n844), .B1(new_n777), .B2(new_n839), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n790), .A2(G311), .B1(new_n815), .B2(G322), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n785), .A2(G317), .B1(G303), .B2(new_n807), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT48), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1059), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n1063), .B2(new_n1062), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT49), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n760), .B(new_n1058), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1057), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1048), .B1(new_n1069), .B2(new_n768), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n1038), .A2(new_n752), .B1(new_n1039), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n748), .A2(new_n1038), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n753), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n748), .A2(new_n1038), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1071), .B1(new_n1073), .B2(new_n1074), .ZN(G393));
  NOR2_X1   g0875(.A1(new_n241), .A2(new_n761), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n769), .B1(new_n579), .B2(new_n216), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n754), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n791), .A2(new_n595), .B1(new_n800), .B2(new_n809), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(G283), .B2(new_n841), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n332), .B1(new_n793), .B2(new_n839), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(G116), .B2(new_n798), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1080), .A2(new_n775), .A3(new_n1082), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n785), .A2(G311), .B1(new_n815), .B2(G317), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT52), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n786), .A2(new_n1051), .B1(new_n787), .B2(new_n963), .ZN(new_n1086));
  XOR2_X1   g0886(.A(KEYINPUT109), .B(KEYINPUT51), .Z(new_n1087));
  OR2_X1    g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1088), .A2(new_n843), .A3(new_n1089), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n790), .A2(G50), .B1(new_n251), .B2(new_n807), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(G68), .A2(new_n841), .B1(new_n816), .B2(G143), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n798), .A2(G77), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1091), .A2(new_n855), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n1083), .A2(new_n1085), .B1(new_n1090), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1078), .B1(new_n1095), .B2(new_n768), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n989), .B2(new_n821), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1003), .A2(KEYINPUT108), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(new_n1002), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1097), .B1(new_n1099), .B2(new_n751), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1072), .A2(new_n1004), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1101), .A2(new_n695), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1072), .A2(new_n1099), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1100), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(G390));
  AOI21_X1  g0905(.A(new_n701), .B1(new_n901), .B2(new_n709), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n899), .B1(new_n1106), .B2(new_n829), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n829), .B1(new_n743), .B2(new_n744), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n932), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n829), .B(new_n899), .C1(new_n729), .C2(new_n733), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1106), .A2(new_n921), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n829), .B1(new_n729), .B2(new_n733), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1115), .B1(new_n1116), .B2(new_n931), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1113), .B1(new_n1117), .B2(new_n933), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n926), .A2(new_n1106), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n635), .B(new_n1119), .C1(new_n747), .C2(new_n447), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT111), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n948), .A2(new_n951), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n949), .B1(new_n933), .B2(new_n931), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT110), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n950), .B1(new_n915), .B2(new_n918), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n742), .A2(new_n677), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT96), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n742), .A2(KEYINPUT96), .A3(new_n677), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n830), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n899), .B1(new_n1134), .B2(new_n932), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1128), .B1(new_n1129), .B2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n949), .B1(new_n946), .B2(new_n947), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n931), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1138));
  NOR3_X1   g0938(.A1(new_n1137), .A2(KEYINPUT110), .A3(new_n1138), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1127), .B(new_n1112), .C1(new_n1136), .C2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1127), .B1(new_n1136), .B2(new_n1139), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n1115), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1124), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(KEYINPUT111), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1140), .ZN(new_n1145));
  OAI21_X1  g0945(.A(KEYINPUT110), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n919), .A2(new_n1135), .A3(new_n1128), .A4(new_n949), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n1146), .A2(new_n1147), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1148), .A2(new_n1114), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1144), .B1(new_n1145), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1143), .A2(new_n1150), .A3(new_n753), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1145), .A2(new_n1149), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1125), .A2(new_n765), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n754), .B1(new_n251), .B2(new_n837), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n790), .A2(G107), .B1(new_n815), .B2(G283), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n579), .B2(new_n793), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n1156), .B(KEYINPUT113), .Z(new_n1157));
  AOI21_X1  g0957(.A(new_n267), .B1(new_n841), .B2(G87), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n785), .A2(G116), .B1(G294), .B2(new_n816), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n861), .A2(new_n1093), .A3(new_n1158), .A4(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(G125), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n791), .A2(new_n848), .B1(new_n800), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(G159), .B2(new_n798), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n777), .A2(new_n963), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT53), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n785), .A2(G132), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(KEYINPUT54), .B(G143), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(G128), .A2(new_n815), .B1(new_n807), .B2(new_n1168), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1163), .A2(new_n1165), .A3(new_n1166), .A4(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n267), .B1(new_n773), .B2(new_n788), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT112), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n1157), .A2(new_n1160), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1154), .B1(new_n1173), .B2(new_n768), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n1152), .A2(new_n752), .B1(new_n1153), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1151), .A2(new_n1175), .ZN(G378));
  INV_X1    g0976(.A(KEYINPUT57), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1140), .B(new_n1118), .C1(new_n1148), .C2(new_n1114), .ZN(new_n1178));
  AND2_X1   g0978(.A1(new_n1178), .A2(new_n1121), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT116), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n632), .A2(new_n633), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1182), .B1(new_n1183), .B2(new_n296), .ZN(new_n1184));
  AOI211_X1 g0984(.A(KEYINPUT116), .B(new_n617), .C1(new_n632), .C2(new_n633), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n885), .B1(new_n256), .B2(new_n265), .ZN(new_n1186));
  XOR2_X1   g0986(.A(new_n1186), .B(KEYINPUT55), .Z(new_n1187));
  NOR3_X1   g0987(.A1(new_n1184), .A2(new_n1185), .A3(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1187), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n312), .A2(KEYINPUT116), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1183), .A2(new_n1182), .A3(new_n296), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1189), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1181), .B1(new_n1188), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT118), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1187), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1190), .A2(new_n1189), .A3(new_n1191), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1195), .A2(new_n1196), .A3(new_n1180), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1193), .A2(new_n1194), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(new_n925), .B2(G330), .ZN(new_n1199));
  OAI211_X1 g0999(.A(KEYINPUT40), .B(new_n902), .C1(new_n946), .C2(new_n947), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n923), .B1(new_n930), .B2(new_n922), .ZN(new_n1201));
  AND4_X1   g1001(.A1(G330), .A2(new_n1200), .A3(new_n1198), .A4(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n953), .B1(new_n1199), .B2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1200), .A2(new_n1201), .A3(G330), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1198), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1200), .A2(new_n1198), .A3(new_n1201), .A4(G330), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1206), .A2(new_n952), .A3(new_n936), .A4(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1203), .A2(KEYINPUT119), .A3(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT119), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n953), .B(new_n1210), .C1(new_n1199), .C2(new_n1202), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1209), .A2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1177), .B1(new_n1179), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1178), .A2(new_n1121), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1177), .B1(new_n1203), .B2(new_n1208), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n695), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1213), .A2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1209), .A2(new_n752), .A3(new_n1211), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n754), .B1(G50), .B2(new_n837), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1193), .A2(new_n765), .A3(new_n1197), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(G33), .A2(G41), .ZN(new_n1221));
  INV_X1    g1021(.A(G124), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1221), .B1(new_n800), .B2(new_n1222), .C1(new_n773), .C2(new_n801), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n785), .A2(G128), .B1(new_n841), .B2(new_n1168), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n1161), .B2(new_n787), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n790), .A2(G132), .B1(G137), .B2(new_n807), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1226), .B(KEYINPUT115), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n1225), .B(new_n1227), .C1(G150), .C2(new_n798), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1223), .B1(new_n1229), .B2(KEYINPUT59), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(KEYINPUT59), .B2(new_n1229), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n760), .A2(new_n282), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1232), .B(new_n788), .C1(G33), .C2(G41), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1050), .B1(new_n844), .B2(new_n800), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n1234), .B(new_n1232), .C1(G58), .C2(new_n965), .ZN(new_n1235));
  XOR2_X1   g1035(.A(new_n1235), .B(KEYINPUT114), .Z(new_n1236));
  OAI22_X1  g1036(.A1(new_n791), .A2(new_n579), .B1(new_n787), .B2(new_n543), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n786), .A2(new_n362), .B1(new_n356), .B2(new_n793), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n1237), .B(new_n1238), .C1(G68), .C2(new_n798), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1236), .A2(KEYINPUT58), .A3(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1236), .A2(new_n1239), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT58), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1231), .A2(new_n1233), .A3(new_n1240), .A4(new_n1243), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n1219), .B(new_n1220), .C1(new_n768), .C2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1218), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1217), .A2(new_n1248), .ZN(G375));
  OAI211_X1 g1049(.A(new_n1113), .B(new_n1120), .C1(new_n1117), .C2(new_n933), .ZN(new_n1250));
  XOR2_X1   g1050(.A(new_n1008), .B(KEYINPUT120), .Z(new_n1251));
  NAND3_X1  g1051(.A1(new_n1122), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n931), .A2(new_n765), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n754), .B1(G68), .B2(new_n837), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1254), .B(KEYINPUT121), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n760), .B1(G50), .B2(new_n798), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n787), .A2(new_n856), .B1(new_n777), .B2(new_n1051), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(G150), .B2(new_n807), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n785), .A2(G137), .B1(G58), .B2(new_n965), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n790), .A2(new_n1168), .B1(new_n816), .B2(G128), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1256), .A2(new_n1258), .A3(new_n1259), .A4(new_n1260), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n791), .A2(new_n543), .B1(new_n793), .B2(new_n362), .ZN(new_n1262));
  OR2_X1    g1062(.A1(new_n1262), .A2(KEYINPUT122), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(KEYINPUT122), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n787), .A2(new_n839), .B1(new_n800), .B2(new_n595), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n267), .B(new_n1265), .C1(G97), .C2(new_n841), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n774), .A2(G77), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1263), .A2(new_n1264), .A3(new_n1266), .A4(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1055), .B1(G283), .B2(new_n785), .ZN(new_n1269));
  XOR2_X1   g1069(.A(new_n1269), .B(KEYINPUT123), .Z(new_n1270));
  OAI21_X1  g1070(.A(new_n1261), .B1(new_n1268), .B2(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1255), .B1(new_n1271), .B2(new_n768), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n1118), .A2(new_n752), .B1(new_n1253), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1252), .A2(new_n1273), .ZN(G381));
  INV_X1    g1074(.A(G384), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1104), .A2(new_n1275), .ZN(new_n1276));
  OR4_X1    g1076(.A1(G396), .A2(new_n1276), .A3(G393), .A4(G381), .ZN(new_n1277));
  OR4_X1    g1077(.A1(G387), .A2(new_n1277), .A3(G375), .A4(G378), .ZN(G407));
  NAND2_X1  g1078(.A1(new_n675), .A2(G213), .ZN(new_n1279));
  OR3_X1    g1079(.A1(G375), .A2(G378), .A3(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(G407), .A2(new_n1280), .A3(G213), .ZN(G409));
  XNOR2_X1  g1081(.A(G393), .B(new_n823), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1012), .B1(new_n1011), .B2(new_n1028), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1034), .A2(KEYINPUT107), .A3(new_n1035), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(G390), .B1(new_n1286), .B2(new_n985), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n985), .ZN(new_n1288));
  AOI211_X1 g1088(.A(new_n1288), .B(new_n1104), .C1(new_n1284), .C2(new_n1285), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1283), .B1(new_n1287), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(G387), .A2(new_n1104), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1286), .A2(new_n985), .A3(G390), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1291), .A2(new_n1282), .A3(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1290), .A2(new_n1293), .ZN(new_n1294));
  AOI221_X4 g1094(.A(new_n1247), .B1(new_n1151), .B2(new_n1175), .C1(new_n1213), .C2(new_n1216), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1203), .A2(new_n1208), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1246), .B1(new_n1296), .B2(new_n751), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1214), .A2(new_n1211), .A3(new_n1209), .A4(new_n1251), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1297), .B1(new_n1298), .B2(KEYINPUT124), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1212), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT124), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1300), .A2(new_n1301), .A3(new_n1214), .A4(new_n1251), .ZN(new_n1302));
  AOI21_X1  g1102(.A(G378), .B1(new_n1299), .B2(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1279), .B1(new_n1295), .B2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT60), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1250), .A2(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n695), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT125), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1250), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1308), .B1(new_n1309), .B2(KEYINPUT60), .ZN(new_n1310));
  NOR3_X1   g1110(.A1(new_n1250), .A2(KEYINPUT125), .A3(new_n1305), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n1306), .B(new_n1307), .C1(new_n1310), .C2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n1273), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1275), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1312), .A2(G384), .A3(new_n1273), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n675), .A2(G213), .A3(G2897), .ZN(new_n1316));
  AND3_X1   g1116(.A1(new_n1314), .A2(new_n1315), .A3(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1316), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  AOI211_X1 g1119(.A(KEYINPUT61), .B(new_n1294), .C1(new_n1304), .C2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  OAI211_X1 g1122(.A(new_n1279), .B(new_n1322), .C1(new_n1295), .C2(new_n1303), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT63), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(KEYINPUT126), .ZN(new_n1326));
  OR2_X1    g1126(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT126), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1323), .A2(new_n1328), .A3(new_n1324), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1320), .A2(new_n1326), .A3(new_n1327), .A4(new_n1329), .ZN(new_n1330));
  AOI21_X1  g1130(.A(KEYINPUT61), .B1(new_n1304), .B2(new_n1319), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1217), .A2(G378), .A3(new_n1248), .ZN(new_n1332));
  AND2_X1   g1132(.A1(new_n1299), .A2(new_n1302), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1332), .B1(new_n1333), .B2(G378), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT62), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1334), .A2(new_n1335), .A3(new_n1279), .A4(new_n1322), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1323), .A2(KEYINPUT62), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1331), .A2(new_n1336), .A3(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1338), .A2(new_n1294), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1330), .A2(new_n1339), .ZN(G405));
  NAND3_X1  g1140(.A1(G375), .A2(new_n1151), .A3(new_n1175), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1341), .A2(new_n1332), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(new_n1322), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1341), .A2(new_n1332), .A3(new_n1321), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  XNOR2_X1  g1145(.A(new_n1345), .B(new_n1294), .ZN(G402));
endmodule


