//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 1 1 1 1 1 1 1 1 1 1 1 0 0 1 0 0 0 0 1 0 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n542, new_n543,
    new_n544, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n560, new_n561, new_n562,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n589, new_n590, new_n591, new_n592, new_n595, new_n596, new_n598,
    new_n599, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1095, new_n1096;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G221), .A3(G220), .A4(G218), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  XOR2_X1   g029(.A(G325), .B(KEYINPUT66), .Z(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n463), .A2(G137), .B1(G101), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n467), .B1(new_n462), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(G160));
  OAI21_X1  g047(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n473));
  INV_X1    g048(.A(G112), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n473), .B1(new_n474), .B2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n462), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT67), .ZN(new_n479));
  AOI211_X1 g054(.A(new_n475), .B(new_n479), .C1(G136), .C2(new_n463), .ZN(G162));
  NAND2_X1  g055(.A1(KEYINPUT4), .A2(G138), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT3), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(new_n464), .ZN(new_n483));
  NAND2_X1  g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(G102), .A2(G2104), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n476), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(G126), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n489), .B1(new_n483), .B2(new_n484), .ZN(new_n490));
  NAND2_X1  g065(.A1(G114), .A2(G2104), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(G2105), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  OAI211_X1 g068(.A(G138), .B(new_n476), .C1(new_n460), .C2(new_n461), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n488), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  XNOR2_X1  g073(.A(KEYINPUT5), .B(G543), .ZN(new_n499));
  XNOR2_X1  g074(.A(KEYINPUT6), .B(G651), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G88), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G50), .ZN(new_n504));
  OAI22_X1  g079(.A1(new_n501), .A2(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n499), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n505), .A2(new_n508), .ZN(G166));
  NAND3_X1  g084(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n510));
  XNOR2_X1  g085(.A(new_n510), .B(KEYINPUT7), .ZN(new_n511));
  INV_X1    g086(.A(G51), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n503), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n499), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n500), .A2(G89), .ZN(new_n515));
  NAND2_X1  g090(.A1(G63), .A2(G651), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT68), .ZN(new_n518));
  OR3_X1    g093(.A1(new_n513), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n513), .B2(new_n517), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(G168));
  AOI22_X1  g096(.A1(new_n499), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n522), .A2(new_n507), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT69), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n501), .ZN(new_n526));
  INV_X1    g101(.A(new_n503), .ZN(new_n527));
  AOI22_X1  g102(.A1(G90), .A2(new_n526), .B1(new_n527), .B2(G52), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n523), .A2(new_n524), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(G171));
  NAND2_X1  g106(.A1(new_n499), .A2(G56), .ZN(new_n532));
  NAND2_X1  g107(.A1(G68), .A2(G543), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n507), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(KEYINPUT70), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(KEYINPUT70), .ZN(new_n536));
  AOI22_X1  g111(.A1(G81), .A2(new_n526), .B1(new_n527), .B2(G43), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G860), .ZN(G153));
  NAND4_X1  g115(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g116(.A1(G1), .A2(G3), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT8), .ZN(new_n543));
  NAND4_X1  g118(.A1(G319), .A2(G483), .A3(G661), .A4(new_n543), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT71), .ZN(G188));
  INV_X1    g120(.A(G53), .ZN(new_n546));
  OAI21_X1  g121(.A(KEYINPUT9), .B1(new_n503), .B2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT9), .ZN(new_n548));
  NAND4_X1  g123(.A1(new_n500), .A2(new_n548), .A3(G53), .A4(G543), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n547), .A2(new_n549), .B1(new_n526), .B2(G91), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n499), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n551), .A2(new_n507), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(KEYINPUT72), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT72), .ZN(new_n554));
  NOR3_X1   g129(.A1(new_n551), .A2(new_n554), .A3(new_n507), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n550), .B1(new_n553), .B2(new_n555), .ZN(G299));
  INV_X1    g131(.A(G171), .ZN(G301));
  AND2_X1   g132(.A1(new_n519), .A2(new_n520), .ZN(G286));
  INV_X1    g133(.A(G166), .ZN(G303));
  OAI21_X1  g134(.A(G651), .B1(new_n499), .B2(G74), .ZN(new_n560));
  INV_X1    g135(.A(G49), .ZN(new_n561));
  INV_X1    g136(.A(G87), .ZN(new_n562));
  OAI221_X1 g137(.A(new_n560), .B1(new_n503), .B2(new_n561), .C1(new_n562), .C2(new_n501), .ZN(G288));
  INV_X1    g138(.A(G86), .ZN(new_n564));
  INV_X1    g139(.A(G48), .ZN(new_n565));
  OAI22_X1  g140(.A1(new_n501), .A2(new_n564), .B1(new_n503), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n499), .A2(G61), .ZN(new_n568));
  NAND2_X1  g143(.A1(G73), .A2(G543), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n507), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT73), .ZN(new_n571));
  AND2_X1   g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n570), .A2(new_n571), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n567), .B1(new_n572), .B2(new_n573), .ZN(G305));
  AOI22_X1  g149(.A1(G85), .A2(new_n526), .B1(new_n527), .B2(G47), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n499), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n507), .B2(new_n576), .ZN(G290));
  NAND2_X1  g152(.A1(new_n526), .A2(G92), .ZN(new_n578));
  XOR2_X1   g153(.A(new_n578), .B(KEYINPUT10), .Z(new_n579));
  NAND2_X1  g154(.A1(G79), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G66), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n514), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(G651), .B1(new_n527), .B2(G54), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(G868), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n586), .B1(new_n585), .B2(G171), .ZN(G284));
  OAI21_X1  g162(.A(new_n586), .B1(new_n585), .B2(G171), .ZN(G321));
  NAND2_X1  g163(.A1(G286), .A2(G868), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n589), .A2(KEYINPUT74), .ZN(new_n590));
  INV_X1    g165(.A(G299), .ZN(new_n591));
  OAI211_X1 g166(.A(new_n589), .B(KEYINPUT74), .C1(new_n591), .C2(G868), .ZN(new_n592));
  AND2_X1   g167(.A1(new_n590), .A2(new_n592), .ZN(G297));
  XNOR2_X1  g168(.A(G297), .B(KEYINPUT75), .ZN(G280));
  INV_X1    g169(.A(new_n584), .ZN(new_n595));
  INV_X1    g170(.A(G559), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n596), .B2(G860), .ZN(G148));
  NAND2_X1  g172(.A1(new_n538), .A2(new_n585), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n584), .A2(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(new_n585), .ZN(G323));
  XNOR2_X1  g175(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g176(.A1(new_n463), .A2(G135), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT76), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n477), .A2(G123), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT77), .ZN(new_n605));
  OR2_X1    g180(.A1(G99), .A2(G2105), .ZN(new_n606));
  OAI211_X1 g181(.A(new_n606), .B(G2104), .C1(G111), .C2(new_n476), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n603), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT78), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n609), .A2(G2096), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(G2096), .ZN(new_n611));
  INV_X1    g186(.A(new_n462), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(new_n465), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT13), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(G2100), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n610), .A2(new_n611), .A3(new_n616), .ZN(G156));
  XOR2_X1   g192(.A(G2451), .B(G2454), .Z(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT16), .ZN(new_n619));
  XNOR2_X1  g194(.A(G1341), .B(G1348), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT14), .ZN(new_n622));
  XNOR2_X1  g197(.A(G2427), .B(G2438), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2430), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT15), .B(G2435), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n622), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(new_n625), .B2(new_n624), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n621), .B(new_n627), .Z(new_n628));
  XNOR2_X1  g203(.A(G2443), .B(G2446), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n630), .A2(new_n631), .A3(G14), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT79), .Z(G401));
  XOR2_X1   g208(.A(G2084), .B(G2090), .Z(new_n634));
  XNOR2_X1  g209(.A(G2067), .B(G2678), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G2072), .B(G2078), .Z(new_n637));
  NOR2_X1   g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT18), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n637), .B(KEYINPUT17), .ZN(new_n640));
  INV_X1    g215(.A(new_n634), .ZN(new_n641));
  INV_X1    g216(.A(new_n635), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n641), .A2(new_n637), .A3(new_n642), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(new_n636), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n639), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2096), .B(G2100), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(G227));
  XOR2_X1   g223(.A(G1971), .B(G1976), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT19), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1956), .B(G2474), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1961), .B(G1966), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AND2_X1   g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  NOR3_X1   g229(.A1(new_n650), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n650), .A2(new_n653), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT20), .Z(new_n657));
  AOI211_X1 g232(.A(new_n655), .B(new_n657), .C1(new_n650), .C2(new_n654), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1991), .B(G1996), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1981), .B(G1986), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(G229));
  INV_X1    g240(.A(G16), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(G22), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n667), .B1(G166), .B2(new_n666), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G1971), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(G23), .ZN(new_n670));
  INV_X1    g245(.A(G288), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n670), .B1(new_n671), .B2(new_n666), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT82), .Z(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT33), .B(G1976), .Z(new_n675));
  AOI21_X1  g250(.A(new_n669), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  MUX2_X1   g251(.A(G6), .B(G305), .S(G16), .Z(new_n677));
  XOR2_X1   g252(.A(KEYINPUT32), .B(G1981), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT81), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n677), .B(new_n679), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n676), .B(new_n680), .C1(new_n675), .C2(new_n674), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n681), .A2(KEYINPUT34), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(KEYINPUT34), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n463), .A2(G131), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n477), .A2(G119), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n476), .A2(G107), .ZN(new_n686));
  OAI21_X1  g261(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n684), .B(new_n685), .C1(new_n686), .C2(new_n687), .ZN(new_n688));
  MUX2_X1   g263(.A(G25), .B(new_n688), .S(G29), .Z(new_n689));
  XOR2_X1   g264(.A(KEYINPUT35), .B(G1991), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  MUX2_X1   g266(.A(G24), .B(G290), .S(G16), .Z(new_n692));
  XOR2_X1   g267(.A(KEYINPUT80), .B(G1986), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NAND4_X1  g269(.A1(new_n682), .A2(new_n683), .A3(new_n691), .A4(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT36), .Z(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT84), .B(KEYINPUT24), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(G29), .B1(new_n698), .B2(G34), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G34), .B2(new_n698), .ZN(new_n700));
  INV_X1    g275(.A(G29), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(G160), .B2(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT85), .Z(new_n703));
  NAND2_X1  g278(.A1(new_n666), .A2(G21), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G168), .B2(new_n666), .ZN(new_n705));
  AOI22_X1  g280(.A1(new_n703), .A2(G2084), .B1(G1966), .B2(new_n705), .ZN(new_n706));
  OAI221_X1 g281(.A(new_n706), .B1(new_n701), .B2(new_n609), .C1(G2084), .C2(new_n703), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n666), .A2(G5), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G171), .B2(new_n666), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT91), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n707), .B1(new_n710), .B2(G1961), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n705), .A2(G1966), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT90), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n711), .B(new_n713), .C1(G1961), .C2(new_n710), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n701), .A2(G27), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G164), .B2(new_n701), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT92), .Z(new_n717));
  NOR2_X1   g292(.A1(new_n717), .A2(G2078), .ZN(new_n718));
  NOR2_X1   g293(.A1(G162), .A2(new_n701), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(new_n701), .B2(G35), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT29), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n718), .B1(new_n722), .B2(G2090), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n595), .A2(G16), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G4), .B2(G16), .ZN(new_n725));
  INV_X1    g300(.A(G1348), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT25), .ZN(new_n727));
  NAND2_X1  g302(.A1(G103), .A2(G2104), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n727), .B1(new_n728), .B2(G2105), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n476), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n463), .A2(G139), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n612), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(new_n476), .B2(new_n732), .ZN(new_n733));
  MUX2_X1   g308(.A(G33), .B(new_n733), .S(G29), .Z(new_n734));
  NOR2_X1   g309(.A1(new_n734), .A2(G2072), .ZN(new_n735));
  AOI22_X1  g310(.A1(new_n725), .A2(new_n726), .B1(KEYINPUT83), .B2(new_n735), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT31), .B(G11), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT88), .B(G28), .ZN(new_n738));
  AOI21_X1  g313(.A(G29), .B1(new_n738), .B2(KEYINPUT30), .ZN(new_n739));
  OAI22_X1  g314(.A1(new_n739), .A2(KEYINPUT89), .B1(KEYINPUT30), .B2(new_n738), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n739), .A2(KEYINPUT89), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n737), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n734), .B2(G2072), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n736), .B(new_n743), .C1(new_n726), .C2(new_n725), .ZN(new_n744));
  NOR2_X1   g319(.A1(G16), .A2(G19), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n539), .B2(G16), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G1341), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n666), .A2(G20), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT23), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n591), .B2(new_n666), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G1956), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n701), .A2(G32), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n477), .A2(G129), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT86), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n463), .A2(G141), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n465), .A2(G105), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT87), .ZN(new_n758));
  NAND3_X1  g333(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT26), .ZN(new_n760));
  NOR3_X1   g335(.A1(new_n756), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n754), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n752), .B1(new_n762), .B2(new_n701), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT27), .B(G1996), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n701), .A2(G26), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT28), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n463), .A2(G140), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n477), .A2(G128), .ZN(new_n769));
  OR2_X1    g344(.A1(G104), .A2(G2105), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n770), .B(G2104), .C1(G116), .C2(new_n476), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n768), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n767), .B1(new_n773), .B2(new_n701), .ZN(new_n774));
  INV_X1    g349(.A(G2067), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n765), .B(new_n776), .C1(KEYINPUT83), .C2(new_n735), .ZN(new_n777));
  NOR4_X1   g352(.A1(new_n744), .A2(new_n747), .A3(new_n751), .A4(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(G2090), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n721), .A2(new_n779), .B1(G2078), .B2(new_n717), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n723), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  NOR3_X1   g356(.A1(new_n696), .A2(new_n714), .A3(new_n781), .ZN(G311));
  INV_X1    g357(.A(G311), .ZN(G150));
  AOI22_X1  g358(.A1(G93), .A2(new_n526), .B1(new_n527), .B2(G55), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n499), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n785), .A2(new_n507), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT93), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n788), .A2(new_n538), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n539), .A2(new_n787), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT38), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n595), .A2(G559), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n794), .A2(KEYINPUT39), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n794), .A2(KEYINPUT39), .ZN(new_n796));
  NOR3_X1   g371(.A1(new_n795), .A2(new_n796), .A3(G860), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n788), .A2(G860), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT37), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n797), .A2(new_n799), .ZN(G145));
  XNOR2_X1  g375(.A(new_n762), .B(new_n733), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n477), .A2(G130), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n476), .A2(G118), .ZN(new_n803));
  OAI21_X1  g378(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G142), .B2(new_n463), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(new_n614), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n801), .B(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(G164), .B(new_n772), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(new_n688), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n808), .B(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n609), .B(G160), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G162), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n811), .B(new_n813), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT94), .B(G37), .Z(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT95), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g393(.A1(new_n788), .A2(new_n585), .ZN(new_n819));
  XNOR2_X1  g394(.A(G290), .B(new_n671), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT96), .ZN(new_n821));
  XNOR2_X1  g396(.A(G305), .B(G303), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n822), .A2(KEYINPUT96), .A3(new_n820), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT42), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n791), .B(new_n599), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n584), .B(G299), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(KEYINPUT41), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n829), .B1(new_n830), .B2(new_n827), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n826), .B(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n819), .B1(new_n832), .B2(new_n585), .ZN(G295));
  OAI21_X1  g408(.A(new_n819), .B1(new_n832), .B2(new_n585), .ZN(G331));
  INV_X1    g409(.A(KEYINPUT44), .ZN(new_n835));
  OAI21_X1  g410(.A(G171), .B1(G286), .B2(KEYINPUT97), .ZN(new_n836));
  AND3_X1   g411(.A1(new_n519), .A2(KEYINPUT97), .A3(new_n520), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n837), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n789), .A2(new_n790), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n791), .A2(new_n839), .A3(new_n838), .ZN(new_n843));
  INV_X1    g418(.A(new_n828), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT99), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n825), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT98), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n843), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n791), .A2(KEYINPUT98), .A3(new_n839), .A4(new_n838), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n850), .A2(new_n842), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(new_n830), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n847), .A2(new_n848), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n825), .A2(KEYINPUT100), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT100), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n856), .B1(new_n823), .B2(new_n824), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT41), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n844), .A2(KEYINPUT101), .A3(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(new_n830), .B2(KEYINPUT101), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n861), .B1(new_n843), .B2(new_n842), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n852), .A2(new_n828), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n858), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT43), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n854), .A2(new_n864), .A3(new_n865), .A4(new_n815), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT102), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(G37), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n854), .A2(new_n869), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n855), .A2(new_n857), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n871), .B1(new_n853), .B2(new_n847), .ZN(new_n872));
  OAI21_X1  g447(.A(KEYINPUT43), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n868), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n866), .A2(new_n867), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n835), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n870), .A2(new_n872), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n877), .A2(KEYINPUT43), .ZN(new_n878));
  AND4_X1   g453(.A1(KEYINPUT43), .A2(new_n854), .A3(new_n864), .A4(new_n815), .ZN(new_n879));
  OAI21_X1  g454(.A(KEYINPUT44), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n876), .A2(new_n880), .ZN(G397));
  NAND3_X1  g456(.A1(new_n466), .A2(G40), .A3(new_n470), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT45), .ZN(new_n884));
  INV_X1    g459(.A(G1384), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n497), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n883), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT103), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n888), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n762), .B(G1996), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n772), .B(new_n775), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n690), .ZN(new_n896));
  NOR3_X1   g471(.A1(new_n895), .A2(new_n896), .A3(new_n688), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n772), .A2(G2067), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n892), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT46), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n900), .B1(new_n891), .B2(G1996), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT125), .ZN(new_n902));
  OAI211_X1 g477(.A(new_n762), .B(new_n894), .C1(new_n900), .C2(G1996), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n892), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT47), .ZN(new_n906));
  INV_X1    g481(.A(new_n895), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n688), .B(new_n690), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n892), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(KEYINPUT126), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n891), .A2(G1986), .A3(G290), .ZN(new_n912));
  XOR2_X1   g487(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n913));
  XNOR2_X1  g488(.A(new_n912), .B(new_n913), .ZN(new_n914));
  OAI221_X1 g489(.A(new_n899), .B1(new_n905), .B2(new_n906), .C1(new_n911), .C2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n915), .B1(new_n906), .B2(new_n905), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT114), .ZN(new_n917));
  INV_X1    g492(.A(G8), .ZN(new_n918));
  NOR2_X1   g493(.A1(G166), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT55), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT106), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n922), .B1(KEYINPUT55), .B2(new_n919), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n920), .A2(KEYINPUT106), .A3(new_n921), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT50), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n497), .A2(new_n926), .A3(new_n885), .ZN(new_n927));
  XOR2_X1   g502(.A(new_n927), .B(KEYINPUT104), .Z(new_n928));
  AOI21_X1  g503(.A(new_n882), .B1(new_n886), .B2(KEYINPUT50), .ZN(new_n929));
  XNOR2_X1  g504(.A(KEYINPUT105), .B(G2090), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n481), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n932), .B1(new_n460), .B2(new_n461), .ZN(new_n933));
  AOI21_X1  g508(.A(G2105), .B1(new_n933), .B2(new_n486), .ZN(new_n934));
  OAI21_X1  g509(.A(G126), .B1(new_n460), .B2(new_n461), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n476), .B1(new_n935), .B2(new_n491), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(G1384), .B1(new_n937), .B2(new_n496), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n882), .B1(new_n938), .B2(KEYINPUT45), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n886), .A2(new_n884), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(G1971), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n918), .B1(new_n931), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT113), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n925), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n946), .B1(new_n945), .B2(new_n944), .ZN(new_n947));
  INV_X1    g522(.A(G2084), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n928), .A2(new_n948), .A3(new_n929), .ZN(new_n949));
  OR2_X1    g524(.A1(new_n949), .A2(KEYINPUT112), .ZN(new_n950));
  INV_X1    g525(.A(G1966), .ZN(new_n951));
  AOI22_X1  g526(.A1(new_n949), .A2(KEYINPUT112), .B1(new_n951), .B2(new_n941), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n918), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n953), .A2(KEYINPUT63), .A3(G168), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n947), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n923), .A2(new_n924), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n944), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n883), .A2(new_n938), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(G8), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n959), .B1(G1976), .B2(new_n671), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT52), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(KEYINPUT107), .B(G1976), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT52), .B1(G288), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n962), .B1(new_n960), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(G1981), .B1(new_n566), .B2(new_n570), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n966), .B1(G305), .B2(G1981), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT108), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT49), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  OAI211_X1 g544(.A(KEYINPUT108), .B(new_n966), .C1(G305), .C2(G1981), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n959), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OAI211_X1 g546(.A(KEYINPUT49), .B(new_n966), .C1(G305), .C2(G1981), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT109), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n972), .B(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT110), .ZN(new_n975));
  AND3_X1   g550(.A1(new_n971), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n975), .B1(new_n971), .B2(new_n974), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n957), .B(new_n965), .C1(new_n976), .C2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n917), .B1(new_n955), .B2(new_n979), .ZN(new_n980));
  NOR4_X1   g555(.A1(new_n947), .A2(new_n954), .A3(new_n978), .A4(KEYINPUT114), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n883), .B1(new_n938), .B2(new_n926), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT111), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n927), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n497), .A2(KEYINPUT111), .A3(new_n926), .A4(new_n885), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n982), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AOI22_X1  g561(.A1(new_n986), .A2(new_n930), .B1(new_n942), .B2(new_n941), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n925), .B1(new_n918), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n979), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n953), .A2(G168), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI22_X1  g566(.A1(new_n980), .A2(new_n981), .B1(new_n991), .B2(KEYINPUT63), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n993), .B1(new_n941), .B2(G2078), .ZN(new_n994));
  OR3_X1    g569(.A1(new_n941), .A2(new_n993), .A3(G2078), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n928), .A2(new_n929), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n994), .B(new_n995), .C1(new_n996), .C2(G1961), .ZN(new_n997));
  AND4_X1   g572(.A1(G171), .A2(new_n979), .A3(new_n988), .A4(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT123), .ZN(new_n1000));
  AOI211_X1 g575(.A(new_n1000), .B(new_n918), .C1(new_n950), .C2(new_n952), .ZN(new_n1001));
  NOR2_X1   g576(.A1(G168), .A2(new_n918), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n999), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1002), .B1(KEYINPUT123), .B2(new_n999), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n990), .B1(new_n953), .B2(new_n1004), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n1003), .A2(new_n1005), .A3(KEYINPUT62), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT62), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n998), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  OR2_X1    g583(.A1(new_n976), .A2(new_n977), .ZN(new_n1009));
  INV_X1    g584(.A(G1976), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1009), .A2(new_n1010), .A3(new_n671), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1011), .B1(G1981), .B2(G305), .ZN(new_n1012));
  INV_X1    g587(.A(new_n959), .ZN(new_n1013));
  INV_X1    g588(.A(new_n957), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1009), .A2(new_n965), .ZN(new_n1015));
  AOI22_X1  g590(.A1(new_n1012), .A2(new_n1013), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n992), .A2(new_n1008), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT124), .ZN(new_n1019));
  NAND3_X1  g594(.A1(G171), .A2(new_n1019), .A3(KEYINPUT54), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1020), .B1(KEYINPUT54), .B2(G171), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n997), .B(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1018), .A2(new_n988), .A3(new_n979), .A4(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n996), .A2(G1348), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n958), .A2(G2067), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n1025), .B(KEYINPUT118), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  OR2_X1    g602(.A1(new_n595), .A2(KEYINPUT121), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n595), .A2(KEYINPUT121), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1027), .A2(KEYINPUT60), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1027), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT60), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1030), .B(new_n1033), .C1(new_n1034), .C2(new_n1028), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n885), .ZN(new_n1036));
  XNOR2_X1  g611(.A(KEYINPUT56), .B(G2072), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n940), .A2(new_n883), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n939), .A2(KEYINPUT116), .A3(new_n940), .A4(new_n1037), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n984), .A2(new_n985), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(new_n929), .ZN(new_n1045));
  INV_X1    g620(.A(G1956), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1043), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  AOI211_X1 g622(.A(KEYINPUT115), .B(G1956), .C1(new_n1044), .C2(new_n929), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1042), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT57), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1051), .B(new_n550), .C1(new_n553), .C2(new_n555), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1049), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT117), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT115), .B1(new_n986), .B2(G1956), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1045), .A2(new_n1043), .A3(new_n1046), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1053), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1055), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1059), .B(new_n1055), .C1(new_n1047), .C2(new_n1048), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1054), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT61), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G1996), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n939), .A2(new_n1066), .A3(new_n940), .ZN(new_n1067));
  XOR2_X1   g642(.A(KEYINPUT58), .B(G1341), .Z(new_n1068));
  NAND2_X1  g643(.A1(new_n958), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n538), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g645(.A(new_n1070), .B(KEYINPUT59), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1064), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1071), .B1(new_n1072), .B2(new_n1054), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT120), .B1(new_n1065), .B2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1059), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT117), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n1076), .A2(new_n1061), .B1(new_n1049), .B2(new_n1053), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1073), .B(KEYINPUT120), .C1(new_n1077), .C2(KEYINPUT61), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1035), .B1(new_n1074), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1054), .B1(new_n1027), .B2(new_n584), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT119), .ZN(new_n1083));
  XNOR2_X1  g658(.A(new_n1082), .B(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1080), .A2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1023), .B1(new_n1085), .B2(KEYINPUT122), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT122), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1080), .A2(new_n1087), .A3(new_n1084), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1017), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n909), .ZN(new_n1090));
  XOR2_X1   g665(.A(G290), .B(G1986), .Z(new_n1091));
  AOI21_X1  g666(.A(new_n891), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n916), .B1(new_n1089), .B2(new_n1092), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g668(.A1(G401), .A2(new_n458), .A3(G227), .ZN(new_n1095));
  AND2_X1   g669(.A1(new_n664), .A2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g670(.A(new_n817), .B(new_n1096), .C1(new_n874), .C2(new_n875), .ZN(G225));
  INV_X1    g671(.A(G225), .ZN(G308));
endmodule


