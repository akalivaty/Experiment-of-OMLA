//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 1 1 0 0 1 0 0 1 0 0 0 1 0 1 0 0 1 1 0 1 1 0 0 0 0 1 0 1 1 1 0 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n806, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G169gat), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n205), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n206), .A2(G197gat), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  AOI21_X1  g008(.A(G197gat), .B1(new_n206), .B2(new_n207), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT88), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n204), .B(new_n205), .ZN(new_n212));
  INV_X1    g011(.A(G197gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT88), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n214), .A2(new_n215), .A3(new_n208), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n211), .A2(KEYINPUT12), .A3(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT12), .B1(new_n211), .B2(new_n216), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G50gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G43gat), .ZN(new_n222));
  INV_X1    g021(.A(G43gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(G50gat), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT89), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT15), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n222), .A2(new_n224), .A3(KEYINPUT89), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT14), .ZN(new_n233));
  INV_X1    g032(.A(G29gat), .ZN(new_n234));
  INV_X1    g033(.A(G36gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT90), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT90), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n238), .A2(new_n233), .A3(new_n234), .A4(new_n235), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n232), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  OAI22_X1  g039(.A1(new_n240), .A2(KEYINPUT91), .B1(new_n234), .B2(new_n235), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT91), .ZN(new_n242));
  AOI211_X1 g041(.A(new_n242), .B(new_n232), .C1(new_n237), .C2(new_n239), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n230), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n224), .A2(KEYINPUT92), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(new_n222), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n224), .A2(KEYINPUT92), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n226), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n236), .A2(new_n231), .B1(G29gat), .B2(G36gat), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n229), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n244), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT17), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G15gat), .B(G22gat), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT16), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n254), .B1(new_n255), .B2(G1gat), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n256), .B1(G1gat), .B2(new_n254), .ZN(new_n257));
  XOR2_X1   g056(.A(new_n257), .B(G8gat), .Z(new_n258));
  NAND3_X1  g057(.A1(new_n244), .A2(KEYINPUT17), .A3(new_n250), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n253), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n258), .ZN(new_n261));
  AOI22_X1  g060(.A1(new_n261), .A2(new_n251), .B1(G229gat), .B2(G233gat), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT93), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n263), .A2(KEYINPUT18), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n260), .A2(new_n262), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(G229gat), .A2(G233gat), .ZN(new_n267));
  XOR2_X1   g066(.A(new_n267), .B(KEYINPUT13), .Z(new_n268));
  INV_X1    g067(.A(new_n251), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n269), .A2(new_n258), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n261), .A2(new_n251), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n268), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n266), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n265), .B1(new_n260), .B2(new_n262), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n220), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n211), .A2(new_n216), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT12), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(new_n217), .ZN(new_n279));
  INV_X1    g078(.A(new_n274), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n279), .A2(new_n280), .A3(new_n272), .A4(new_n266), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n275), .A2(new_n281), .A3(KEYINPUT94), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT94), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n220), .B(new_n283), .C1(new_n274), .C2(new_n273), .ZN(new_n284));
  AND3_X1   g083(.A1(new_n282), .A2(new_n284), .A3(KEYINPUT95), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT95), .B1(new_n282), .B2(new_n284), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G232gat), .A2(G233gat), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n289), .A2(KEYINPUT41), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n290), .B(KEYINPUT101), .ZN(new_n291));
  INV_X1    g090(.A(G134gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n293), .B(G162gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n289), .A2(KEYINPUT41), .ZN(new_n295));
  NAND2_X1  g094(.A1(G85gat), .A2(G92gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n296), .B(KEYINPUT7), .ZN(new_n297));
  NAND2_X1  g096(.A1(G99gat), .A2(G106gat), .ZN(new_n298));
  INV_X1    g097(.A(G85gat), .ZN(new_n299));
  INV_X1    g098(.A(G92gat), .ZN(new_n300));
  AOI22_X1  g099(.A1(KEYINPUT8), .A2(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G99gat), .ZN(new_n303));
  INV_X1    g102(.A(G106gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n302), .A2(new_n298), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n298), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n297), .A2(new_n307), .A3(new_n301), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n295), .B1(new_n269), .B2(new_n309), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n253), .A2(new_n259), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(new_n309), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT102), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT102), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n311), .A2(new_n314), .A3(new_n309), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n310), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT103), .ZN(new_n317));
  XNOR2_X1  g116(.A(G190gat), .B(G218gat), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n316), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT103), .B1(new_n316), .B2(new_n319), .ZN(new_n321));
  AOI211_X1 g120(.A(new_n318), .B(new_n310), .C1(new_n313), .C2(new_n315), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n294), .B(new_n320), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT104), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n313), .A2(new_n315), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n324), .B(new_n318), .C1(new_n325), .C2(new_n310), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT104), .B1(new_n316), .B2(new_n319), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n294), .B1(new_n316), .B2(new_n319), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n323), .A2(new_n329), .ZN(new_n330));
  XOR2_X1   g129(.A(G71gat), .B(G78gat), .Z(new_n331));
  XNOR2_X1  g130(.A(G57gat), .B(G64gat), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT9), .B1(new_n333), .B2(KEYINPUT96), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT96), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n331), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n331), .A2(new_n332), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(KEYINPUT97), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT98), .B(KEYINPUT21), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(G231gat), .A2(G233gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n344), .B(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G127gat), .B(G155gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n347), .B(KEYINPUT20), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n346), .B(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT100), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n342), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n337), .A2(KEYINPUT100), .A3(new_n341), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n351), .A2(KEYINPUT21), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(new_n258), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(G183gat), .ZN(new_n355));
  INV_X1    g154(.A(G183gat), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n353), .A2(new_n356), .A3(new_n258), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n349), .B(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT99), .B(KEYINPUT19), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(G211gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n359), .B(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT105), .B1(new_n330), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n361), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n359), .B(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT105), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n365), .A2(new_n323), .A3(new_n329), .A4(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT10), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n309), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n351), .A2(new_n369), .A3(new_n352), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT106), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT106), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n351), .A2(new_n369), .A3(new_n372), .A4(new_n352), .ZN(new_n373));
  OR2_X1    g172(.A1(new_n342), .A2(new_n309), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n342), .A2(new_n309), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n374), .A2(new_n368), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n371), .A2(new_n373), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(G230gat), .A2(G233gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n374), .A2(new_n375), .ZN(new_n380));
  INV_X1    g179(.A(new_n378), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G176gat), .B(G204gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n384), .B(G148gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(KEYINPUT107), .B(G120gat), .ZN(new_n386));
  XOR2_X1   g185(.A(new_n385), .B(new_n386), .Z(new_n387));
  OR2_X1    g186(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n383), .A2(new_n387), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n363), .A2(new_n367), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(G228gat), .A2(G233gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(G155gat), .A2(G162gat), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(G155gat), .A2(G162gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  XOR2_X1   g196(.A(KEYINPUT75), .B(KEYINPUT2), .Z(new_n398));
  INV_X1    g197(.A(G148gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(G141gat), .ZN(new_n400));
  INV_X1    g199(.A(G141gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(G148gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n397), .B1(new_n398), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n401), .A2(KEYINPUT76), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT76), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(G141gat), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(new_n407), .A3(G148gat), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT2), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n409), .ZN(new_n410));
  AOI22_X1  g209(.A1(new_n408), .A2(new_n400), .B1(new_n396), .B2(new_n410), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n404), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT3), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT29), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G197gat), .B(G204gat), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT22), .ZN(new_n416));
  INV_X1    g215(.A(G211gat), .ZN(new_n417));
  INV_X1    g216(.A(G218gat), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  XOR2_X1   g219(.A(G211gat), .B(G218gat), .Z(new_n421));
  XNOR2_X1  g220(.A(new_n420), .B(new_n421), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n414), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT29), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n412), .B1(new_n425), .B2(new_n413), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n393), .B1(new_n423), .B2(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(KEYINPUT81), .ZN(new_n428));
  XOR2_X1   g227(.A(new_n422), .B(KEYINPUT71), .Z(new_n429));
  OAI211_X1 g228(.A(G228gat), .B(G233gat), .C1(new_n429), .C2(new_n414), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n427), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  XNOR2_X1  g230(.A(KEYINPUT31), .B(G50gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n432), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n434), .B(new_n427), .C1(new_n428), .C2(new_n430), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(G78gat), .B(G106gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n437), .B(G22gat), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n433), .A2(new_n438), .A3(new_n435), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(KEYINPUT82), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT82), .B1(new_n440), .B2(new_n441), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(G127gat), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n446), .A2(G134gat), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n292), .A2(G127gat), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT68), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n292), .A2(G127gat), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n446), .A2(G134gat), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT68), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT1), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n454), .B1(G113gat), .B2(G120gat), .ZN(new_n455));
  AND2_X1   g254(.A1(G113gat), .A2(G120gat), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n449), .A2(new_n453), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT69), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT69), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n449), .A2(new_n460), .A3(new_n453), .A4(new_n457), .ZN(new_n461));
  INV_X1    g260(.A(new_n457), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n450), .A2(new_n451), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n459), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n412), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT77), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n412), .A2(new_n459), .A3(new_n461), .A4(new_n464), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(G225gat), .A2(G233gat), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n465), .A2(KEYINPUT77), .A3(new_n466), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n470), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n469), .A2(KEYINPUT4), .ZN(new_n475));
  AOI22_X1  g274(.A1(new_n458), .A2(KEYINPUT69), .B1(new_n463), .B2(new_n462), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT4), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n476), .A2(new_n477), .A3(new_n461), .A4(new_n412), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT3), .B1(new_n404), .B2(new_n411), .ZN(new_n479));
  XNOR2_X1  g278(.A(G141gat), .B(G148gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(KEYINPUT75), .B(KEYINPUT2), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n396), .B(new_n395), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  AND2_X1   g281(.A1(new_n408), .A2(new_n400), .ZN(new_n483));
  AND2_X1   g282(.A1(new_n410), .A2(new_n396), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n482), .B(new_n413), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n479), .A2(new_n485), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n475), .A2(new_n478), .B1(new_n465), .B2(new_n486), .ZN(new_n487));
  AOI22_X1  g286(.A1(new_n474), .A2(KEYINPUT5), .B1(new_n487), .B2(new_n471), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n475), .A2(new_n478), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n486), .A2(new_n465), .ZN(new_n490));
  AND4_X1   g289(.A1(KEYINPUT5), .A2(new_n489), .A3(new_n471), .A4(new_n490), .ZN(new_n491));
  XOR2_X1   g290(.A(G57gat), .B(G85gat), .Z(new_n492));
  XNOR2_X1  g291(.A(G1gat), .B(G29gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n492), .B(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n495));
  XOR2_X1   g294(.A(new_n494), .B(new_n495), .Z(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NOR3_X1   g296(.A1(new_n488), .A2(new_n491), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT6), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n497), .B1(new_n488), .B2(new_n491), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT79), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT6), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT79), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n504), .B(new_n497), .C1(new_n488), .C2(new_n491), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n502), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT80), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n498), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n502), .A2(KEYINPUT80), .A3(new_n503), .A4(new_n505), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n500), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(G226gat), .ZN(new_n511));
  INV_X1    g310(.A(G233gat), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT27), .B1(new_n356), .B2(KEYINPUT67), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT67), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT27), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n517), .A3(G183gat), .ZN(new_n518));
  INV_X1    g317(.A(G190gat), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n515), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT28), .ZN(new_n521));
  XNOR2_X1  g320(.A(KEYINPUT27), .B(G183gat), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n521), .A2(G190gat), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n520), .A2(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(G169gat), .A2(G176gat), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT26), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(G169gat), .A2(G176gat), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(G183gat), .A2(G190gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OR2_X1    g331(.A1(new_n524), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n525), .A2(KEYINPUT66), .A3(KEYINPUT23), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT25), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n536), .B(new_n529), .C1(new_n525), .C2(KEYINPUT23), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT66), .B1(new_n525), .B2(KEYINPUT23), .ZN(new_n538));
  NOR3_X1   g337(.A1(new_n535), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT65), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g341(.A1(KEYINPUT65), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT24), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n531), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n356), .A2(new_n519), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n542), .A2(new_n543), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n545), .A2(new_n540), .A3(new_n546), .ZN(new_n548));
  INV_X1    g347(.A(G176gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n205), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT23), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n525), .A2(KEYINPUT23), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n548), .A2(new_n529), .A3(new_n552), .A4(new_n553), .ZN(new_n554));
  AOI22_X1  g353(.A1(new_n539), .A2(new_n547), .B1(new_n554), .B2(KEYINPUT25), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n514), .B1(new_n533), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(KEYINPUT25), .ZN(new_n557));
  INV_X1    g356(.A(new_n537), .ZN(new_n558));
  INV_X1    g357(.A(new_n538), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n547), .A2(new_n558), .A3(new_n534), .A4(new_n559), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n557), .B(new_n560), .C1(new_n524), .C2(new_n532), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n424), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n556), .B1(new_n514), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(new_n422), .ZN(new_n564));
  XNOR2_X1  g363(.A(G8gat), .B(G36gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(G64gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(new_n300), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT29), .B1(new_n533), .B2(new_n555), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT72), .B1(new_n568), .B2(new_n513), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT72), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n562), .A2(new_n570), .A3(new_n514), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n556), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n564), .B(new_n567), .C1(new_n572), .C2(new_n429), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT30), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n556), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n570), .B1(new_n562), .B2(new_n514), .ZN(new_n577));
  AOI211_X1 g376(.A(KEYINPUT72), .B(new_n513), .C1(new_n561), .C2(new_n424), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n429), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n581), .A2(KEYINPUT30), .A3(new_n564), .A4(new_n567), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n564), .B1(new_n572), .B2(new_n429), .ZN(new_n583));
  INV_X1    g382(.A(new_n567), .ZN(new_n584));
  AOI22_X1  g383(.A1(new_n582), .A2(KEYINPUT73), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g384(.A1(new_n579), .A2(new_n580), .B1(new_n422), .B2(new_n563), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT73), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n586), .A2(new_n587), .A3(KEYINPUT30), .A4(new_n567), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT74), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(KEYINPUT73), .B1(new_n573), .B2(new_n574), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n583), .A2(new_n584), .ZN(new_n591));
  AND4_X1   g390(.A1(KEYINPUT74), .A2(new_n590), .A3(new_n588), .A4(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n575), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n445), .B1(new_n510), .B2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G15gat), .B(G43gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(G71gat), .B(G99gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  OR3_X1    g396(.A1(new_n561), .A2(new_n465), .A3(KEYINPUT70), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n561), .A2(new_n465), .ZN(new_n599));
  OAI21_X1  g398(.A(KEYINPUT70), .B1(new_n561), .B2(new_n465), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G227gat), .A2(G233gat), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n602), .B(KEYINPUT64), .Z(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT33), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n597), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(KEYINPUT32), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI211_X1 g407(.A(new_n604), .B(KEYINPUT32), .C1(new_n605), .C2(new_n597), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n601), .A2(new_n603), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n611), .B(KEYINPUT34), .Z(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n611), .B(KEYINPUT34), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n614), .A2(new_n609), .A3(new_n608), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT36), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  AND3_X1   g417(.A1(new_n594), .A2(KEYINPUT83), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT83), .B1(new_n594), .B2(new_n618), .ZN(new_n620));
  XOR2_X1   g419(.A(KEYINPUT85), .B(KEYINPUT38), .Z(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n567), .B1(new_n583), .B2(KEYINPUT37), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT87), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(KEYINPUT86), .B(KEYINPUT37), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n586), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n627), .B1(new_n623), .B2(new_n624), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n622), .B1(new_n625), .B2(new_n628), .ZN(new_n629));
  AOI211_X1 g428(.A(new_n567), .B(new_n622), .C1(new_n586), .C2(new_n626), .ZN(new_n630));
  OAI22_X1  g429(.A1(new_n579), .A2(new_n580), .B1(new_n422), .B2(new_n563), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(KEYINPUT37), .ZN(new_n632));
  AOI22_X1  g431(.A1(new_n630), .A2(new_n632), .B1(new_n586), .B2(new_n567), .ZN(new_n633));
  INV_X1    g432(.A(new_n498), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n502), .A2(new_n634), .A3(new_n503), .A4(new_n505), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n629), .A2(new_n633), .A3(new_n499), .A4(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n440), .A2(new_n441), .ZN(new_n637));
  INV_X1    g436(.A(new_n487), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT84), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n638), .A2(new_n639), .A3(new_n472), .ZN(new_n640));
  OAI21_X1  g439(.A(KEYINPUT84), .B1(new_n487), .B2(new_n471), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n470), .A2(new_n473), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n471), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n640), .A2(KEYINPUT39), .A3(new_n641), .A4(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(new_n497), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT40), .ZN(new_n646));
  AOI21_X1  g445(.A(KEYINPUT39), .B1(new_n640), .B2(new_n641), .ZN(new_n647));
  OR3_X1    g446(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n585), .A2(new_n575), .A3(new_n588), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n646), .B1(new_n645), .B2(new_n647), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n648), .A2(new_n649), .A3(new_n634), .A4(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n636), .A2(new_n637), .A3(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NOR3_X1   g452(.A1(new_n619), .A2(new_n620), .A3(new_n653), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n613), .A2(new_n615), .ZN(new_n655));
  INV_X1    g454(.A(new_n649), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n655), .A2(new_n637), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n635), .A2(new_n499), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT35), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n506), .A2(new_n507), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n662), .A2(new_n634), .A3(new_n509), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(new_n499), .ZN(new_n664));
  INV_X1    g463(.A(new_n637), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n665), .A2(new_n616), .ZN(new_n666));
  INV_X1    g465(.A(new_n575), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n590), .A2(new_n588), .A3(new_n591), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT74), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n585), .A2(KEYINPUT74), .A3(new_n588), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n667), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n664), .A2(new_n666), .A3(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n661), .B1(KEYINPUT35), .B2(new_n673), .ZN(new_n674));
  OAI211_X1 g473(.A(new_n287), .B(new_n392), .C1(new_n654), .C2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT108), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n287), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT83), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT82), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n637), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n442), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n682), .B1(new_n664), .B2(new_n672), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n616), .B(KEYINPUT36), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n679), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n594), .A2(KEYINPUT83), .A3(new_n618), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n685), .A2(new_n686), .A3(new_n652), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n673), .A2(KEYINPUT35), .ZN(new_n688));
  INV_X1    g487(.A(new_n661), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n678), .B1(new_n687), .B2(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n691), .A2(KEYINPUT108), .A3(new_n392), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n510), .ZN(new_n694));
  XOR2_X1   g493(.A(KEYINPUT109), .B(G1gat), .Z(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1324gat));
  XOR2_X1   g495(.A(KEYINPUT16), .B(G8gat), .Z(new_n697));
  NAND3_X1  g496(.A1(new_n693), .A2(new_n649), .A3(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT42), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n693), .A2(KEYINPUT42), .A3(new_n649), .A4(new_n697), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n594), .A2(new_n618), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n653), .B1(new_n702), .B2(new_n679), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n674), .B1(new_n703), .B2(new_n686), .ZN(new_n704));
  NOR4_X1   g503(.A1(new_n704), .A2(new_n676), .A3(new_n678), .A4(new_n391), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT108), .B1(new_n691), .B2(new_n392), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(G8gat), .B1(new_n707), .B2(new_n656), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n700), .A2(new_n701), .A3(new_n708), .ZN(G1325gat));
  OR3_X1    g508(.A1(new_n707), .A2(G15gat), .A3(new_n616), .ZN(new_n710));
  OR2_X1    g509(.A1(new_n618), .A2(KEYINPUT110), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n618), .A2(KEYINPUT110), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(G15gat), .B1(new_n707), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n710), .A2(new_n714), .ZN(G1326gat));
  XNOR2_X1  g514(.A(KEYINPUT43), .B(G22gat), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT111), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n718), .B1(new_n693), .B2(new_n445), .ZN(new_n719));
  AOI211_X1 g518(.A(KEYINPUT111), .B(new_n682), .C1(new_n677), .C2(new_n692), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n717), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(KEYINPUT111), .B1(new_n707), .B2(new_n682), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n693), .A2(new_n718), .A3(new_n445), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n722), .A2(new_n716), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n721), .A2(new_n724), .ZN(G1327gat));
  INV_X1    g524(.A(new_n390), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n365), .A2(new_n726), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n282), .A2(new_n284), .A3(KEYINPUT112), .ZN(new_n728));
  AOI21_X1  g527(.A(KEYINPUT112), .B1(new_n282), .B2(new_n284), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  XOR2_X1   g530(.A(new_n731), .B(KEYINPUT113), .Z(new_n732));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n594), .A2(new_n652), .A3(new_n618), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n733), .B(new_n330), .C1(new_n734), .C2(new_n674), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT114), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n594), .A2(new_n652), .A3(new_n618), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n690), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n739), .A2(KEYINPUT114), .A3(new_n733), .A4(new_n330), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n330), .ZN(new_n742));
  OAI21_X1  g541(.A(KEYINPUT44), .B1(new_n704), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n732), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n234), .B1(new_n744), .B2(new_n510), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n727), .A2(new_n330), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n664), .A2(G29gat), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n691), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT45), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n749), .B(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(KEYINPUT115), .B1(new_n745), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n749), .B(KEYINPUT45), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT115), .ZN(new_n754));
  AOI211_X1 g553(.A(new_n664), .B(new_n732), .C1(new_n741), .C2(new_n743), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n753), .B(new_n754), .C1(new_n755), .C2(new_n234), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n752), .A2(new_n756), .ZN(G1328gat));
  AOI21_X1  g556(.A(new_n235), .B1(new_n744), .B2(new_n649), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n656), .A2(G36gat), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n691), .A2(new_n747), .A3(new_n759), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT46), .ZN(new_n761));
  OAI21_X1  g560(.A(KEYINPUT116), .B1(new_n758), .B2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT46), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n760), .B(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT116), .ZN(new_n765));
  AOI211_X1 g564(.A(new_n656), .B(new_n732), .C1(new_n741), .C2(new_n743), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n764), .B(new_n765), .C1(new_n766), .C2(new_n235), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n762), .A2(new_n767), .ZN(G1329gat));
  AND4_X1   g567(.A1(new_n223), .A2(new_n691), .A3(new_n655), .A4(new_n747), .ZN(new_n769));
  INV_X1    g568(.A(new_n713), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n744), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n769), .B1(new_n771), .B2(G43gat), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n223), .B1(new_n744), .B2(new_n684), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT47), .ZN(new_n774));
  OR2_X1    g573(.A1(new_n769), .A2(new_n774), .ZN(new_n775));
  OAI22_X1  g574(.A1(new_n772), .A2(KEYINPUT47), .B1(new_n773), .B2(new_n775), .ZN(G1330gat));
  AND4_X1   g575(.A1(new_n221), .A2(new_n691), .A3(new_n445), .A4(new_n747), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n744), .A2(new_n445), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n777), .B1(new_n778), .B2(G50gat), .ZN(new_n779));
  XNOR2_X1  g578(.A(KEYINPUT117), .B(KEYINPUT48), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n221), .B1(new_n744), .B2(new_n665), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT48), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n777), .A2(new_n782), .ZN(new_n783));
  OAI22_X1  g582(.A1(new_n779), .A2(new_n780), .B1(new_n781), .B2(new_n783), .ZN(G1331gat));
  INV_X1    g583(.A(new_n730), .ZN(new_n785));
  AND4_X1   g584(.A1(new_n363), .A2(new_n367), .A3(new_n785), .A4(new_n726), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n739), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(new_n510), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g588(.A(new_n656), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(KEYINPUT118), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(KEYINPUT119), .ZN(new_n793));
  NOR2_X1   g592(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n793), .B(new_n794), .ZN(G1333gat));
  INV_X1    g594(.A(G71gat), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n796), .B1(new_n787), .B2(new_n770), .ZN(new_n797));
  AND4_X1   g596(.A1(new_n796), .A2(new_n739), .A3(new_n655), .A4(new_n786), .ZN(new_n798));
  OR3_X1    g597(.A1(new_n797), .A2(new_n798), .A3(KEYINPUT120), .ZN(new_n799));
  OAI21_X1  g598(.A(KEYINPUT120), .B1(new_n797), .B2(new_n798), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT50), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n799), .A2(KEYINPUT50), .A3(new_n800), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(G1334gat));
  NAND2_X1  g604(.A1(new_n787), .A2(new_n445), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g606(.A1(new_n730), .A2(new_n365), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n726), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n809), .B1(new_n741), .B2(new_n743), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n299), .B1(new_n810), .B2(new_n510), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n739), .A2(new_n330), .A3(new_n808), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(KEYINPUT51), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT51), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n739), .A2(new_n814), .A3(new_n330), .A4(new_n808), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n813), .A2(new_n726), .A3(new_n815), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n816), .A2(G85gat), .A3(new_n664), .ZN(new_n817));
  OR2_X1    g616(.A1(new_n811), .A2(new_n817), .ZN(G1336gat));
  AOI21_X1  g617(.A(new_n300), .B1(new_n810), .B2(new_n649), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n816), .A2(G92gat), .A3(new_n656), .ZN(new_n820));
  OAI21_X1  g619(.A(KEYINPUT52), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n816), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n822), .A2(new_n300), .A3(new_n649), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n824));
  AOI211_X1 g623(.A(new_n656), .B(new_n809), .C1(new_n741), .C2(new_n743), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n823), .B(new_n824), .C1(new_n825), .C2(new_n300), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n821), .A2(new_n826), .ZN(G1337gat));
  AOI21_X1  g626(.A(G99gat), .B1(new_n822), .B2(new_n655), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n713), .A2(new_n303), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n828), .B1(new_n810), .B2(new_n829), .ZN(G1338gat));
  NOR2_X1   g629(.A1(new_n637), .A2(G106gat), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n816), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n810), .A2(new_n445), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n833), .B1(new_n834), .B2(G106gat), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n836), .B1(new_n816), .B2(new_n832), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n304), .B1(new_n810), .B2(new_n665), .ZN(new_n838));
  OAI22_X1  g637(.A1(new_n835), .A2(new_n836), .B1(new_n837), .B2(new_n838), .ZN(G1339gat));
  NAND2_X1  g638(.A1(new_n282), .A2(new_n284), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT112), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT55), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n371), .A2(new_n376), .A3(new_n381), .A4(new_n373), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n379), .A2(KEYINPUT54), .A3(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n377), .A2(new_n847), .A3(new_n378), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n387), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n843), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n845), .A2(KEYINPUT55), .A3(new_n387), .A4(new_n848), .ZN(new_n851));
  AND3_X1   g650(.A1(new_n850), .A2(new_n388), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n282), .A2(new_n284), .A3(KEYINPUT112), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n842), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n270), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n267), .B1(new_n855), .B2(new_n260), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n270), .A2(new_n271), .A3(new_n268), .ZN(new_n857));
  OAI22_X1  g656(.A1(new_n856), .A2(new_n857), .B1(new_n209), .B2(new_n210), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n281), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n390), .A2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n330), .B1(new_n854), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n850), .A2(new_n388), .A3(new_n851), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(new_n859), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n330), .A2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n362), .B1(new_n862), .B2(new_n866), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n363), .A2(new_n367), .A3(new_n785), .A4(new_n390), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n445), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n869), .A2(new_n510), .A3(new_n655), .A4(new_n656), .ZN(new_n870));
  INV_X1    g669(.A(G113gat), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n870), .A2(new_n871), .A3(new_n678), .ZN(new_n872));
  AOI211_X1 g671(.A(new_n664), .B(new_n657), .C1(new_n867), .C2(new_n868), .ZN(new_n873));
  AOI21_X1  g672(.A(G113gat), .B1(new_n873), .B2(new_n730), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n872), .A2(new_n874), .ZN(G1340gat));
  INV_X1    g674(.A(G120gat), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n870), .A2(new_n876), .A3(new_n390), .ZN(new_n877));
  AOI21_X1  g676(.A(G120gat), .B1(new_n873), .B2(new_n726), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n877), .A2(new_n878), .ZN(G1341gat));
  OAI21_X1  g678(.A(G127gat), .B1(new_n870), .B2(new_n362), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n873), .A2(new_n446), .A3(new_n365), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(G1342gat));
  NAND3_X1  g681(.A1(new_n873), .A2(new_n292), .A3(new_n330), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n883), .A2(KEYINPUT56), .ZN(new_n884));
  OAI21_X1  g683(.A(G134gat), .B1(new_n870), .B2(new_n742), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(KEYINPUT56), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(G1343gat));
  AND2_X1   g686(.A1(new_n405), .A2(new_n407), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT57), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n728), .A2(new_n729), .A3(new_n863), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n742), .B1(new_n891), .B2(new_n860), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n365), .B1(new_n892), .B2(new_n865), .ZN(new_n893));
  AND4_X1   g692(.A1(new_n363), .A2(new_n367), .A3(new_n785), .A4(new_n390), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n890), .B(new_n665), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n618), .A2(new_n510), .A3(new_n656), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT95), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n840), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n282), .A2(new_n284), .A3(KEYINPUT95), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n899), .A2(new_n852), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n330), .B1(new_n901), .B2(new_n861), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n362), .B1(new_n902), .B2(new_n866), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n682), .B1(new_n903), .B2(new_n868), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n895), .B(new_n897), .C1(new_n890), .C2(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n889), .B1(new_n905), .B2(new_n678), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT58), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n664), .B1(new_n867), .B2(new_n868), .ZN(new_n908));
  AOI211_X1 g707(.A(new_n637), .B(new_n649), .C1(new_n711), .C2(new_n712), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n287), .A2(new_n401), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n910), .B(KEYINPUT121), .ZN(new_n911));
  AND3_X1   g710(.A1(new_n908), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n906), .A2(new_n907), .A3(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT122), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n889), .B1(new_n905), .B2(new_n785), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n913), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n915), .B1(new_n917), .B2(KEYINPUT58), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n285), .A2(new_n286), .A3(new_n863), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n742), .B1(new_n919), .B2(new_n860), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n365), .B1(new_n920), .B2(new_n865), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n445), .B1(new_n921), .B2(new_n894), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(KEYINPUT57), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n923), .A2(new_n730), .A3(new_n895), .A4(new_n897), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n912), .B1(new_n924), .B2(new_n889), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n925), .A2(KEYINPUT122), .A3(new_n907), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n914), .B1(new_n918), .B2(new_n926), .ZN(G1344gat));
  INV_X1    g726(.A(KEYINPUT59), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n928), .B(G148gat), .C1(new_n905), .C2(new_n390), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT124), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n391), .A2(new_n287), .ZN(new_n931));
  OAI211_X1 g730(.A(new_n890), .B(new_n445), .C1(new_n931), .C2(new_n921), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n726), .B1(new_n896), .B2(KEYINPUT123), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n933), .B1(new_n896), .B2(KEYINPUT123), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n637), .B1(new_n867), .B2(new_n868), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n932), .B(new_n934), .C1(new_n890), .C2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(G148gat), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n930), .B1(new_n937), .B2(KEYINPUT59), .ZN(new_n938));
  AOI211_X1 g737(.A(KEYINPUT124), .B(new_n928), .C1(new_n936), .C2(G148gat), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n929), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n908), .A2(new_n909), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n941), .A2(new_n399), .A3(new_n726), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n940), .A2(new_n942), .ZN(G1345gat));
  OAI21_X1  g742(.A(G155gat), .B1(new_n905), .B2(new_n362), .ZN(new_n944));
  INV_X1    g743(.A(G155gat), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n941), .A2(new_n945), .A3(new_n365), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n944), .A2(new_n946), .ZN(G1346gat));
  OAI21_X1  g746(.A(G162gat), .B1(new_n905), .B2(new_n742), .ZN(new_n948));
  INV_X1    g747(.A(G162gat), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n941), .A2(new_n949), .A3(new_n330), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(G1347gat));
  NAND4_X1  g750(.A1(new_n869), .A2(new_n664), .A3(new_n655), .A4(new_n649), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n952), .A2(new_n205), .A3(new_n678), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n867), .A2(new_n868), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(new_n664), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n656), .B1(new_n955), .B2(KEYINPUT125), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT125), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n954), .A2(new_n957), .A3(new_n664), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n956), .A2(new_n666), .A3(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(new_n730), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n953), .B1(new_n961), .B2(new_n205), .ZN(G1348gat));
  OAI21_X1  g761(.A(G176gat), .B1(new_n952), .B2(new_n390), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n726), .A2(new_n549), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n963), .B1(new_n959), .B2(new_n964), .ZN(G1349gat));
  OAI21_X1  g764(.A(G183gat), .B1(new_n952), .B2(new_n362), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n365), .A2(new_n522), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n966), .B1(new_n959), .B2(new_n967), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n968), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g768(.A1(new_n960), .A2(new_n519), .A3(new_n330), .ZN(new_n970));
  OAI21_X1  g769(.A(G190gat), .B1(new_n952), .B2(new_n742), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n971), .A2(KEYINPUT61), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n971), .A2(KEYINPUT61), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n970), .B1(new_n972), .B2(new_n973), .ZN(G1351gat));
  OR2_X1    g773(.A1(new_n935), .A2(new_n890), .ZN(new_n975));
  NOR3_X1   g774(.A1(new_n770), .A2(new_n510), .A3(new_n656), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n975), .A2(new_n932), .A3(new_n976), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n977), .A2(new_n213), .A3(new_n678), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n770), .A2(new_n637), .ZN(new_n979));
  AND3_X1   g778(.A1(new_n956), .A2(new_n979), .A3(new_n958), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(new_n730), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n978), .B1(new_n981), .B2(new_n213), .ZN(G1352gat));
  OR2_X1    g781(.A1(new_n977), .A2(new_n390), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n390), .A2(G204gat), .ZN(new_n984));
  NAND4_X1  g783(.A1(new_n956), .A2(new_n979), .A3(new_n958), .A4(new_n984), .ZN(new_n985));
  AOI22_X1  g784(.A1(new_n983), .A2(G204gat), .B1(KEYINPUT62), .B2(new_n985), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT126), .ZN(new_n987));
  OR3_X1    g786(.A1(new_n985), .A2(new_n987), .A3(KEYINPUT62), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n987), .B1(new_n985), .B2(KEYINPUT62), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n986), .A2(new_n988), .A3(new_n989), .ZN(G1353gat));
  NAND4_X1  g789(.A1(new_n975), .A2(new_n365), .A3(new_n932), .A4(new_n976), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n991), .A2(G211gat), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT63), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n991), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n994), .A2(KEYINPUT127), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g795(.A(KEYINPUT63), .B1(new_n991), .B2(G211gat), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT127), .ZN(new_n998));
  NOR2_X1   g797(.A1(new_n362), .A2(G211gat), .ZN(new_n999));
  AOI22_X1  g798(.A1(new_n997), .A2(new_n998), .B1(new_n980), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n996), .A2(new_n1000), .ZN(G1354gat));
  NOR3_X1   g800(.A1(new_n977), .A2(new_n418), .A3(new_n742), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n980), .A2(new_n330), .ZN(new_n1003));
  AOI21_X1  g802(.A(new_n1002), .B1(new_n1003), .B2(new_n418), .ZN(G1355gat));
endmodule


