//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 0 1 0 0 1 0 1 1 0 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 1 0 1 0 0 1 0 0 1 1 0 0 0 0 0 0 0 0 1 0 1 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n826, new_n827, new_n828,
    new_n829, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n970, new_n971;
  OAI21_X1  g000(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT23), .ZN(new_n203));
  INV_X1    g002(.A(G169gat), .ZN(new_n204));
  INV_X1    g003(.A(G176gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT65), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g008(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n210));
  AOI22_X1  g009(.A1(new_n202), .A2(new_n206), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n212), .B(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(KEYINPUT67), .B(G190gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n215), .B1(new_n216), .B2(G183gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n211), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT25), .ZN(new_n219));
  OR4_X1    g018(.A1(KEYINPUT69), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT69), .B1(new_n221), .B2(KEYINPUT26), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(KEYINPUT26), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n220), .A2(new_n222), .A3(new_n223), .A4(new_n207), .ZN(new_n224));
  INV_X1    g023(.A(new_n216), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT28), .ZN(new_n226));
  INV_X1    g025(.A(G183gat), .ZN(new_n227));
  OR3_X1    g026(.A1(new_n227), .A2(KEYINPUT68), .A3(KEYINPUT27), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT27), .B1(new_n227), .B2(KEYINPUT68), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n225), .A2(new_n226), .A3(new_n228), .A4(new_n229), .ZN(new_n230));
  XOR2_X1   g029(.A(KEYINPUT27), .B(G183gat), .Z(new_n231));
  OAI21_X1  g030(.A(KEYINPUT28), .B1(new_n231), .B2(new_n216), .ZN(new_n232));
  NAND2_X1  g031(.A1(G183gat), .A2(G190gat), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n224), .A2(new_n230), .A3(new_n232), .A4(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT25), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n215), .B1(G183gat), .B2(G190gat), .ZN(new_n236));
  OR2_X1    g035(.A1(new_n236), .A2(new_n212), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT64), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n206), .A2(new_n202), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n238), .B1(new_n239), .B2(new_n207), .ZN(new_n240));
  AND2_X1   g039(.A1(G169gat), .A2(G176gat), .ZN(new_n241));
  AOI211_X1 g040(.A(KEYINPUT64), .B(new_n241), .C1(new_n206), .C2(new_n202), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n235), .B(new_n237), .C1(new_n240), .C2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n219), .A2(new_n234), .A3(new_n243), .ZN(new_n244));
  AND2_X1   g043(.A1(G226gat), .A2(G233gat), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT29), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n244), .A2(new_n248), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n219), .A2(new_n234), .A3(new_n243), .A4(new_n246), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G197gat), .B(G204gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(KEYINPUT22), .ZN(new_n253));
  NAND2_X1  g052(.A1(G211gat), .A2(G218gat), .ZN(new_n254));
  OR2_X1    g053(.A1(G211gat), .A2(G218gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n253), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT74), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT22), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n254), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(new_n252), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT74), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n253), .A2(new_n261), .A3(new_n254), .A4(new_n255), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n257), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n251), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n249), .A2(new_n250), .A3(new_n263), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(new_n266), .A3(KEYINPUT75), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT75), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n251), .A2(new_n268), .A3(new_n264), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G8gat), .B(G36gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT76), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n272), .B(G64gat), .Z(new_n273));
  XNOR2_X1  g072(.A(new_n273), .B(G92gat), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT30), .B1(new_n270), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n274), .B1(new_n267), .B2(new_n269), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(KEYINPUT30), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT77), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n277), .A2(KEYINPUT77), .A3(KEYINPUT30), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n279), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  AND2_X1   g084(.A1(G155gat), .A2(G162gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(G155gat), .A2(G162gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n288), .B(KEYINPUT78), .ZN(new_n289));
  XNOR2_X1  g088(.A(G141gat), .B(G148gat), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G155gat), .A2(G162gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT2), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT79), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n296), .B1(new_n286), .B2(new_n287), .ZN(new_n297));
  INV_X1    g096(.A(G155gat), .ZN(new_n298));
  INV_X1    g097(.A(G162gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n300), .A2(KEYINPUT79), .A3(new_n292), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT80), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n293), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n292), .A2(KEYINPUT80), .A3(KEYINPUT2), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n302), .A2(new_n306), .A3(new_n291), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n307), .A2(KEYINPUT81), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT81), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n290), .B1(new_n297), .B2(new_n301), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n309), .B1(new_n310), .B2(new_n306), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n295), .B1(new_n308), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT3), .ZN(new_n313));
  XOR2_X1   g112(.A(G127gat), .B(G134gat), .Z(new_n314));
  INV_X1    g113(.A(KEYINPUT70), .ZN(new_n315));
  XNOR2_X1  g114(.A(G113gat), .B(G120gat), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n314), .B(new_n315), .C1(KEYINPUT1), .C2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G113gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G120gat), .ZN(new_n319));
  INV_X1    g118(.A(G120gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G113gat), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT1), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G127gat), .B(G134gat), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT70), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n317), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT1), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT72), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n319), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n318), .A2(KEYINPUT72), .A3(G120gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  OR2_X1    g129(.A1(KEYINPUT71), .A2(G120gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(KEYINPUT71), .A2(G120gat), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n318), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n326), .B(new_n323), .C1(new_n330), .C2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n325), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT82), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n325), .A2(KEYINPUT82), .A3(new_n334), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT3), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n340), .B(new_n295), .C1(new_n308), .C2(new_n311), .ZN(new_n341));
  AND3_X1   g140(.A1(new_n313), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT86), .ZN(new_n343));
  NOR3_X1   g142(.A1(new_n312), .A2(KEYINPUT4), .A3(new_n335), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT4), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n307), .A2(KEYINPUT81), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n310), .A2(new_n309), .A3(new_n306), .ZN(new_n347));
  AOI22_X1  g146(.A1(new_n346), .A2(new_n347), .B1(new_n294), .B2(new_n289), .ZN(new_n348));
  INV_X1    g147(.A(new_n335), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n345), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n343), .B1(new_n344), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT4), .B1(new_n312), .B2(new_n335), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n348), .A2(new_n345), .A3(new_n349), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n352), .A2(KEYINPUT86), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n342), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G225gat), .A2(G233gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n357), .A2(KEYINPUT5), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT5), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n348), .A2(new_n349), .ZN(new_n361));
  AND3_X1   g160(.A1(new_n325), .A2(KEYINPUT82), .A3(new_n334), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT82), .B1(new_n325), .B2(new_n334), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n361), .B1(new_n364), .B2(new_n348), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n360), .B1(new_n365), .B2(new_n357), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n352), .A2(new_n353), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n313), .A2(new_n339), .A3(new_n341), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n367), .A2(new_n356), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT83), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n366), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n370), .B1(new_n366), .B2(new_n369), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n359), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G57gat), .B(G85gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n374), .B(G29gat), .ZN(new_n375));
  XOR2_X1   g174(.A(KEYINPUT84), .B(KEYINPUT0), .Z(new_n376));
  XNOR2_X1  g175(.A(new_n375), .B(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT85), .B(G1gat), .ZN(new_n378));
  XOR2_X1   g177(.A(new_n377), .B(new_n378), .Z(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n373), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT6), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n379), .B(new_n359), .C1(new_n371), .C2(new_n372), .ZN(new_n383));
  AND3_X1   g182(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n373), .A2(KEYINPUT6), .A3(new_n380), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n285), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G78gat), .B(G106gat), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n263), .B1(new_n341), .B2(new_n247), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n263), .A2(new_n247), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n348), .B1(new_n391), .B2(new_n340), .ZN(new_n392));
  NAND2_X1  g191(.A1(G228gat), .A2(G233gat), .ZN(new_n393));
  NOR3_X1   g192(.A1(new_n390), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT29), .B1(new_n348), .B2(new_n340), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n256), .A2(new_n260), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT3), .B1(new_n397), .B2(new_n247), .ZN(new_n398));
  OAI22_X1  g197(.A1(new_n396), .A2(new_n263), .B1(new_n348), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT88), .B1(new_n399), .B2(new_n393), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n348), .A2(new_n398), .ZN(new_n401));
  OAI211_X1 g200(.A(KEYINPUT88), .B(new_n393), .C1(new_n390), .C2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n395), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(G22gat), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n393), .B1(new_n390), .B2(new_n401), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT88), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n402), .ZN(new_n409));
  INV_X1    g208(.A(G22gat), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n410), .A3(new_n395), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n405), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT87), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n389), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  AOI211_X1 g213(.A(KEYINPUT87), .B(new_n388), .C1(new_n405), .C2(new_n411), .ZN(new_n415));
  XNOR2_X1  g214(.A(KEYINPUT31), .B(G50gat), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NOR3_X1   g216(.A1(new_n414), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n410), .B1(new_n409), .B2(new_n395), .ZN(new_n419));
  AOI211_X1 g218(.A(G22gat), .B(new_n394), .C1(new_n408), .C2(new_n402), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n413), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n388), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n412), .A2(new_n413), .A3(new_n389), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n416), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n387), .B1(new_n418), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n244), .A2(new_n349), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n335), .A2(new_n219), .A3(new_n234), .A4(new_n243), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(G227gat), .ZN(new_n429));
  INV_X1    g228(.A(G233gat), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n426), .A2(new_n431), .A3(new_n427), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT32), .ZN(new_n435));
  XNOR2_X1  g234(.A(G15gat), .B(G43gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n436), .B(G71gat), .ZN(new_n437));
  INV_X1    g236(.A(G99gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT33), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n434), .A2(KEYINPUT73), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT73), .B1(new_n434), .B2(new_n440), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n435), .B(new_n439), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT34), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n439), .A2(KEYINPUT33), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n434), .A2(KEYINPUT32), .A3(new_n445), .ZN(new_n446));
  AND3_X1   g245(.A1(new_n443), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n444), .B1(new_n443), .B2(new_n446), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n433), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n443), .A2(new_n446), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT34), .ZN(new_n451));
  INV_X1    g250(.A(new_n433), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n443), .A2(new_n444), .A3(new_n446), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT36), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n455), .B(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n417), .B1(new_n414), .B2(new_n415), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n422), .A2(new_n423), .A3(new_n416), .ZN(new_n459));
  OR2_X1    g258(.A1(new_n365), .A2(new_n357), .ZN(new_n460));
  OAI211_X1 g259(.A(KEYINPUT39), .B(new_n460), .C1(new_n355), .C2(new_n356), .ZN(new_n461));
  NOR3_X1   g260(.A1(new_n344), .A2(new_n350), .A3(new_n343), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT86), .B1(new_n352), .B2(new_n353), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n368), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT39), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n464), .A2(new_n465), .A3(new_n357), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n461), .A2(new_n466), .A3(KEYINPUT40), .A4(new_n379), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n461), .A2(new_n379), .A3(new_n466), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT90), .ZN(new_n469));
  XOR2_X1   g268(.A(KEYINPUT89), .B(KEYINPUT40), .Z(new_n470));
  AND3_X1   g269(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n469), .B1(new_n468), .B2(new_n470), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n467), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n284), .A2(new_n381), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n458), .B(new_n459), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT37), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n275), .B1(new_n270), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n477), .B1(new_n476), .B2(new_n270), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n277), .B1(new_n478), .B2(KEYINPUT38), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT38), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n265), .A2(new_n266), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n477), .B(new_n481), .C1(new_n476), .C2(new_n482), .ZN(new_n483));
  AND4_X1   g282(.A1(new_n385), .A2(new_n479), .A3(new_n480), .A4(new_n483), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n425), .B(new_n457), .C1(new_n475), .C2(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n284), .B1(new_n480), .B2(new_n385), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n449), .A2(new_n454), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n458), .A2(new_n486), .A3(new_n487), .A4(new_n459), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT35), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n418), .A2(new_n424), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n491), .A2(KEYINPUT35), .A3(new_n487), .A4(new_n486), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n485), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(KEYINPUT94), .B(KEYINPUT17), .ZN(new_n494));
  OAI22_X1  g293(.A1(KEYINPUT91), .A2(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(KEYINPUT91), .A2(KEYINPUT14), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(G29gat), .ZN(new_n499));
  INV_X1    g298(.A(G36gat), .ZN(new_n500));
  AND4_X1   g299(.A1(KEYINPUT91), .A2(new_n499), .A3(new_n500), .A4(KEYINPUT14), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT92), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(G50gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(G43gat), .ZN(new_n504));
  INV_X1    g303(.A(G43gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(G50gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(new_n506), .A3(KEYINPUT15), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n499), .A2(new_n500), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT91), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT14), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n508), .A2(new_n511), .A3(new_n496), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT92), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n499), .A2(new_n500), .A3(KEYINPUT91), .A4(KEYINPUT14), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n504), .A2(new_n506), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT15), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n516), .A2(new_n517), .B1(G29gat), .B2(G36gat), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n502), .A2(new_n507), .A3(new_n515), .A4(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT93), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n512), .B(new_n514), .C1(new_n499), .C2(new_n500), .ZN(new_n521));
  INV_X1    g320(.A(new_n507), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n519), .A2(new_n520), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n520), .B1(new_n519), .B2(new_n523), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n494), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(G15gat), .B(G22gat), .ZN(new_n527));
  INV_X1    g326(.A(G1gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT16), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n530), .B1(G1gat), .B2(new_n527), .ZN(new_n531));
  XOR2_X1   g330(.A(new_n531), .B(G8gat), .Z(new_n532));
  NAND3_X1  g331(.A1(new_n519), .A2(KEYINPUT17), .A3(new_n523), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n526), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n532), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n535), .B1(new_n524), .B2(new_n525), .ZN(new_n536));
  NAND2_X1  g335(.A1(G229gat), .A2(G233gat), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n534), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT18), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n524), .A2(new_n525), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(new_n532), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n536), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n537), .B(KEYINPUT13), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n534), .A2(new_n536), .A3(KEYINPUT18), .A4(new_n537), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n540), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G113gat), .B(G141gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(G197gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT11), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(new_n204), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(KEYINPUT12), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n548), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n540), .A2(new_n553), .A3(new_n546), .A4(new_n547), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(G230gat), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n559), .A2(new_n430), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(G57gat), .B(G64gat), .Z(new_n562));
  OR2_X1    g361(.A1(G71gat), .A2(G78gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(G71gat), .A2(G78gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n562), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G57gat), .B(G64gat), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n564), .B(new_n563), .C1(new_n569), .C2(new_n566), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(G85gat), .ZN(new_n572));
  INV_X1    g371(.A(G92gat), .ZN(new_n573));
  OAI21_X1  g372(.A(KEYINPUT7), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT7), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n575), .A2(G85gat), .A3(G92gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G99gat), .A2(G106gat), .ZN(new_n578));
  AOI22_X1  g377(.A1(KEYINPUT8), .A2(new_n578), .B1(new_n572), .B2(new_n573), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(G99gat), .B(G106gat), .Z(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n577), .A2(new_n581), .A3(new_n579), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT97), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n571), .A2(new_n583), .A3(new_n584), .A4(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n568), .A2(new_n570), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT97), .B1(new_n577), .B2(new_n579), .ZN(new_n589));
  INV_X1    g388(.A(new_n584), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n581), .B1(new_n577), .B2(new_n579), .ZN(new_n591));
  OAI22_X1  g390(.A1(new_n588), .A2(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT10), .B1(new_n587), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n583), .A2(new_n584), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n594), .A2(KEYINPUT10), .A3(new_n571), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n561), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n587), .A2(new_n560), .A3(new_n592), .ZN(new_n598));
  XNOR2_X1  g397(.A(G120gat), .B(G148gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(new_n205), .ZN(new_n600));
  INV_X1    g399(.A(G204gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n597), .A2(new_n598), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT98), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n603), .B1(new_n597), .B2(new_n598), .ZN(new_n607));
  OR3_X1    g406(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n606), .B1(new_n605), .B2(new_n607), .ZN(new_n609));
  AND2_X1   g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n558), .A2(new_n610), .ZN(new_n611));
  AND2_X1   g410(.A1(new_n493), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n594), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n526), .A2(new_n613), .A3(new_n533), .ZN(new_n614));
  NAND3_X1  g413(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n594), .B1(new_n524), .B2(new_n525), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(G190gat), .ZN(new_n618));
  INV_X1    g417(.A(G190gat), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n614), .A2(new_n619), .A3(new_n615), .A4(new_n616), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(G218gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n618), .A2(G218gat), .A3(new_n620), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n623), .A2(KEYINPUT96), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G134gat), .B(G162gat), .ZN(new_n628));
  INV_X1    g427(.A(new_n626), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n623), .A2(KEYINPUT96), .A3(new_n629), .A4(new_n624), .ZN(new_n630));
  AND3_X1   g429(.A1(new_n627), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n628), .B1(new_n627), .B2(new_n630), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT21), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n532), .B1(new_n634), .B2(new_n588), .ZN(new_n635));
  XOR2_X1   g434(.A(G127gat), .B(G155gat), .Z(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  AND2_X1   g436(.A1(G231gat), .A2(G233gat), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n641), .A2(new_n634), .A3(new_n588), .ZN(new_n642));
  OAI211_X1 g441(.A(new_n639), .B(new_n640), .C1(KEYINPUT21), .C2(new_n571), .ZN(new_n643));
  XNOR2_X1  g442(.A(G183gat), .B(G211gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT20), .ZN(new_n645));
  XNOR2_X1  g444(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  AND3_X1   g446(.A1(new_n642), .A2(new_n643), .A3(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n647), .B1(new_n642), .B2(new_n643), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n633), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n612), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n384), .A2(new_n386), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(new_n528), .ZN(G1324gat));
  NOR2_X1   g456(.A1(new_n653), .A2(new_n285), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(G8gat), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT42), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT16), .B(G8gat), .ZN(new_n662));
  OR3_X1    g461(.A1(new_n659), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n662), .B(KEYINPUT99), .Z(new_n664));
  NAND2_X1  g463(.A1(new_n658), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT100), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n665), .A2(new_n666), .A3(new_n661), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n666), .B1(new_n665), .B2(new_n661), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n660), .B(new_n663), .C1(new_n668), .C2(new_n669), .ZN(G1325gat));
  INV_X1    g469(.A(new_n653), .ZN(new_n671));
  AOI21_X1  g470(.A(G15gat), .B1(new_n671), .B2(new_n487), .ZN(new_n672));
  INV_X1    g471(.A(new_n457), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(G15gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT101), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n672), .B1(new_n671), .B2(new_n675), .ZN(G1326gat));
  NOR2_X1   g475(.A1(new_n653), .A2(new_n491), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT43), .B(G22gat), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1327gat));
  NAND2_X1  g478(.A1(new_n493), .A2(new_n633), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n651), .A2(new_n611), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n682), .A2(new_n499), .A3(new_n654), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT45), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n680), .A2(KEYINPUT44), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n493), .A2(new_n686), .A3(new_n633), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n681), .B(KEYINPUT102), .Z(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(G29gat), .B1(new_n690), .B2(new_n655), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n684), .A2(new_n691), .ZN(G1328gat));
  OAI21_X1  g491(.A(G36gat), .B1(new_n690), .B2(new_n285), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n682), .A2(new_n500), .A3(new_n284), .ZN(new_n694));
  OR2_X1    g493(.A1(new_n694), .A2(KEYINPUT103), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT46), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(KEYINPUT103), .ZN(new_n697));
  AND3_X1   g496(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n696), .B1(new_n695), .B2(new_n697), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n693), .B1(new_n698), .B2(new_n699), .ZN(G1329gat));
  NAND2_X1  g499(.A1(new_n627), .A2(new_n630), .ZN(new_n701));
  INV_X1    g500(.A(new_n628), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n627), .A2(new_n628), .A3(new_n630), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n488), .B(KEYINPUT35), .ZN(new_n706));
  AOI211_X1 g505(.A(KEYINPUT44), .B(new_n705), .C1(new_n706), .C2(new_n485), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n686), .B1(new_n493), .B2(new_n633), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n673), .B(new_n689), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(KEYINPUT104), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT104), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n688), .A2(new_n711), .A3(new_n673), .A4(new_n689), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n710), .A2(new_n712), .A3(G43gat), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n682), .A2(new_n505), .A3(new_n487), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n713), .A2(KEYINPUT47), .A3(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n714), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n716), .B1(new_n709), .B2(G43gat), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n715), .B1(KEYINPUT47), .B2(new_n717), .ZN(G1330gat));
  INV_X1    g517(.A(new_n491), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n688), .A2(new_n719), .A3(new_n689), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(G50gat), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT105), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n682), .A2(new_n503), .A3(new_n719), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT48), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n723), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n721), .B(new_n724), .C1(new_n722), .C2(KEYINPUT48), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(G1331gat));
  INV_X1    g528(.A(new_n610), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n650), .B(new_n558), .C1(new_n631), .C2(new_n632), .ZN(new_n731));
  AOI211_X1 g530(.A(new_n730), .B(new_n731), .C1(new_n706), .C2(new_n485), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n654), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g533(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n732), .A2(new_n284), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT106), .ZN(new_n737));
  NOR2_X1   g536(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(G1333gat));
  NAND3_X1  g538(.A1(new_n732), .A2(G71gat), .A3(new_n673), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n732), .A2(new_n487), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n741), .B2(G71gat), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g542(.A1(new_n732), .A2(new_n719), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g544(.A1(new_n650), .A2(new_n557), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n688), .A2(new_n654), .A3(new_n610), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(G85gat), .ZN(new_n748));
  INV_X1    g547(.A(new_n746), .ZN(new_n749));
  OR3_X1    g548(.A1(new_n680), .A2(KEYINPUT51), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(KEYINPUT51), .B1(new_n680), .B2(new_n749), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n750), .A2(new_n572), .A3(new_n751), .A4(new_n610), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n748), .B1(new_n655), .B2(new_n752), .ZN(G1336gat));
  OAI211_X1 g552(.A(new_n610), .B(new_n746), .C1(new_n707), .C2(new_n708), .ZN(new_n754));
  OAI21_X1  g553(.A(G92gat), .B1(new_n754), .B2(new_n285), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n285), .A2(G92gat), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n750), .A2(new_n610), .A3(new_n751), .A4(new_n756), .ZN(new_n757));
  AOI211_X1 g556(.A(KEYINPUT107), .B(KEYINPUT52), .C1(new_n755), .C2(new_n757), .ZN(new_n758));
  OR2_X1    g557(.A1(KEYINPUT107), .A2(KEYINPUT52), .ZN(new_n759));
  NAND2_X1  g558(.A1(KEYINPUT107), .A2(KEYINPUT52), .ZN(new_n760));
  AND4_X1   g559(.A1(new_n759), .A2(new_n755), .A3(new_n760), .A4(new_n757), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n758), .A2(new_n761), .ZN(G1337gat));
  NOR3_X1   g561(.A1(new_n754), .A2(new_n438), .A3(new_n457), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n750), .A2(new_n610), .A3(new_n751), .A4(new_n487), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n763), .B1(new_n438), .B2(new_n764), .ZN(G1338gat));
  OAI21_X1  g564(.A(G106gat), .B1(new_n754), .B2(new_n491), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT108), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n491), .A2(G106gat), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n750), .A2(new_n610), .A3(new_n751), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n768), .A2(new_n771), .A3(KEYINPUT53), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n766), .B(new_n770), .C1(new_n767), .C2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(G1339gat));
  INV_X1    g574(.A(KEYINPUT10), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n586), .A2(new_n570), .A3(new_n568), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n777), .A2(new_n594), .ZN(new_n778));
  AOI22_X1  g577(.A1(new_n571), .A2(new_n586), .B1(new_n583), .B2(new_n584), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n776), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n780), .A2(new_n560), .A3(new_n595), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n781), .A2(new_n597), .A3(KEYINPUT54), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n783), .B(new_n561), .C1(new_n593), .C2(new_n596), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n782), .A2(KEYINPUT55), .A3(new_n602), .A4(new_n784), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n785), .A2(new_n604), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n784), .A2(new_n602), .ZN(new_n787));
  AOI211_X1 g586(.A(KEYINPUT109), .B(KEYINPUT55), .C1(new_n787), .C2(new_n782), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT109), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n782), .A2(new_n602), .A3(new_n784), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT55), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n786), .B1(new_n788), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(KEYINPUT110), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT110), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n795), .B(new_n786), .C1(new_n788), .C2(new_n792), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n558), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n543), .A2(new_n545), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n537), .B1(new_n534), .B2(new_n536), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n552), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(KEYINPUT111), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT111), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n802), .B(new_n552), .C1(new_n798), .C2(new_n799), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n801), .A2(new_n556), .A3(new_n803), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n730), .A2(new_n804), .ZN(new_n805));
  OAI22_X1  g604(.A1(new_n631), .A2(new_n632), .B1(new_n797), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n804), .B1(new_n794), .B2(new_n796), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n703), .A2(new_n704), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n650), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n731), .A2(new_n610), .ZN(new_n810));
  OR2_X1    g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n719), .A2(new_n455), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n811), .A2(new_n654), .A3(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n813), .A2(new_n284), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(KEYINPUT112), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT112), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n816), .B1(new_n813), .B2(new_n284), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(G113gat), .B1(new_n818), .B2(new_n558), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n814), .A2(new_n318), .A3(new_n557), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(G1340gat));
  OAI21_X1  g620(.A(G120gat), .B1(new_n818), .B2(new_n730), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n331), .A2(new_n332), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n814), .A2(new_n823), .A3(new_n610), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(G1341gat));
  NAND4_X1  g624(.A1(new_n815), .A2(G127gat), .A3(new_n817), .A4(new_n650), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n826), .A2(KEYINPUT113), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n826), .A2(KEYINPUT113), .ZN(new_n828));
  AOI21_X1  g627(.A(G127gat), .B1(new_n814), .B2(new_n650), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(G1342gat));
  NOR2_X1   g629(.A1(new_n813), .A2(G134gat), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n633), .A2(new_n285), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(KEYINPUT114), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  XOR2_X1   g633(.A(new_n834), .B(KEYINPUT56), .Z(new_n835));
  OAI21_X1  g634(.A(G134gat), .B1(new_n818), .B2(new_n705), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(G1343gat));
  INV_X1    g636(.A(new_n804), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n610), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n790), .A2(new_n791), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n557), .A2(new_n786), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n705), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n650), .B1(new_n843), .B2(new_n808), .ZN(new_n844));
  OAI211_X1 g643(.A(KEYINPUT57), .B(new_n719), .C1(new_n844), .C2(new_n810), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(KEYINPUT116), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n703), .A2(new_n704), .A3(new_n807), .ZN(new_n847));
  AOI22_X1  g646(.A1(new_n703), .A2(new_n704), .B1(new_n839), .B2(new_n841), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n651), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n849), .B1(new_n610), .B2(new_n731), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n850), .A2(new_n851), .A3(KEYINPUT57), .A4(new_n719), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n719), .B1(new_n809), .B2(new_n810), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n846), .A2(new_n852), .A3(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n655), .A2(new_n284), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(KEYINPUT115), .A3(new_n457), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(KEYINPUT115), .B1(new_n857), .B2(new_n457), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n856), .A2(new_n557), .A3(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT120), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n856), .A2(KEYINPUT120), .A3(new_n557), .A4(new_n861), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n864), .A2(G141gat), .A3(new_n865), .ZN(new_n866));
  XOR2_X1   g665(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n867));
  OAI21_X1  g666(.A(new_n654), .B1(new_n809), .B2(new_n810), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT117), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n673), .A2(new_n491), .ZN(new_n871));
  OAI211_X1 g670(.A(KEYINPUT117), .B(new_n654), .C1(new_n809), .C2(new_n810), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT118), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n870), .A2(KEYINPUT118), .A3(new_n871), .A4(new_n872), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n284), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n558), .A2(G141gat), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n867), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n866), .A2(new_n879), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n862), .A2(G141gat), .ZN(new_n881));
  NOR4_X1   g680(.A1(new_n873), .A2(G141gat), .A3(new_n558), .A4(new_n284), .ZN(new_n882));
  OAI21_X1  g681(.A(KEYINPUT58), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n880), .A2(new_n883), .ZN(G1344gat));
  INV_X1    g683(.A(G148gat), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n877), .A2(new_n885), .A3(new_n610), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n856), .A2(new_n861), .ZN(new_n887));
  AOI211_X1 g686(.A(KEYINPUT59), .B(new_n885), .C1(new_n887), .C2(new_n610), .ZN(new_n888));
  INV_X1    g687(.A(new_n793), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n633), .A2(new_n889), .A3(new_n838), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n650), .B1(new_n890), .B2(new_n843), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n854), .B(new_n719), .C1(new_n891), .C2(new_n810), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n853), .A2(KEYINPUT57), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(new_n893), .A3(new_n610), .ZN(new_n894));
  INV_X1    g693(.A(new_n861), .ZN(new_n895));
  OAI21_X1  g694(.A(G148gat), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n896), .A2(new_n897), .A3(KEYINPUT59), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n897), .B1(new_n896), .B2(KEYINPUT59), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n886), .B1(new_n888), .B2(new_n900), .ZN(G1345gat));
  AOI21_X1  g700(.A(G155gat), .B1(new_n877), .B2(new_n650), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n856), .A2(new_n861), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n903), .A2(new_n298), .A3(new_n651), .ZN(new_n904));
  OAI21_X1  g703(.A(KEYINPUT122), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n887), .A2(G155gat), .A3(new_n650), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT122), .ZN(new_n907));
  AOI211_X1 g706(.A(new_n651), .B(new_n284), .C1(new_n875), .C2(new_n876), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n906), .B(new_n907), .C1(new_n908), .C2(G155gat), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n905), .A2(new_n909), .ZN(G1346gat));
  OAI21_X1  g709(.A(G162gat), .B1(new_n903), .B2(new_n705), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n875), .A2(new_n876), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n912), .A2(new_n299), .A3(new_n833), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(G1347gat));
  NAND2_X1  g713(.A1(new_n655), .A2(new_n284), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n811), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n812), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n918), .A2(new_n558), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(new_n204), .ZN(G1348gat));
  INV_X1    g719(.A(new_n918), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(new_n610), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT123), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n922), .A2(new_n923), .A3(G176gat), .ZN(new_n924));
  XOR2_X1   g723(.A(KEYINPUT123), .B(G176gat), .Z(new_n925));
  OAI21_X1  g724(.A(new_n924), .B1(new_n922), .B2(new_n925), .ZN(G1349gat));
  INV_X1    g725(.A(KEYINPUT60), .ZN(new_n927));
  INV_X1    g726(.A(new_n231), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n917), .A2(new_n650), .A3(new_n928), .A4(new_n812), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT124), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(G183gat), .B1(new_n918), .B2(new_n651), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n932), .A2(new_n929), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n927), .B(new_n931), .C1(new_n933), .C2(new_n930), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n930), .B1(new_n932), .B2(new_n929), .ZN(new_n935));
  INV_X1    g734(.A(new_n931), .ZN(new_n936));
  OAI21_X1  g735(.A(KEYINPUT60), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n934), .A2(new_n937), .ZN(G1350gat));
  AOI21_X1  g737(.A(new_n619), .B1(new_n921), .B2(new_n633), .ZN(new_n939));
  OR2_X1    g738(.A1(new_n939), .A2(KEYINPUT61), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n921), .A2(new_n633), .A3(new_n225), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(KEYINPUT61), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(G1351gat));
  AND2_X1   g742(.A1(new_n892), .A2(new_n893), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n916), .A2(new_n457), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(G197gat), .B1(new_n947), .B2(new_n558), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n811), .A2(new_n719), .A3(new_n946), .ZN(new_n949));
  OR3_X1    g748(.A1(new_n949), .A2(G197gat), .A3(new_n558), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT125), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n951), .B(new_n952), .ZN(G1352gat));
  INV_X1    g752(.A(KEYINPUT126), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n954), .B1(new_n947), .B2(new_n730), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n944), .A2(KEYINPUT126), .A3(new_n610), .A4(new_n946), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n955), .A2(G204gat), .A3(new_n956), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n949), .A2(G204gat), .A3(new_n730), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n958), .B(KEYINPUT62), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n957), .A2(new_n959), .ZN(G1353gat));
  INV_X1    g759(.A(KEYINPUT127), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT63), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI211_X1 g762(.A(G211gat), .B(new_n963), .C1(new_n947), .C2(new_n651), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n961), .A2(new_n962), .ZN(new_n965));
  OR2_X1    g764(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OR3_X1    g765(.A1(new_n949), .A2(G211gat), .A3(new_n651), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n964), .A2(new_n965), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(G1354gat));
  NOR3_X1   g768(.A1(new_n947), .A2(new_n622), .A3(new_n705), .ZN(new_n970));
  OR2_X1    g769(.A1(new_n949), .A2(new_n705), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n970), .B1(new_n622), .B2(new_n971), .ZN(G1355gat));
endmodule


