//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 0 1 1 1 1 0 1 0 0 1 0 0 1 1 1 0 0 0 0 1 1 1 0 1 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014;
  OR2_X1    g000(.A1(KEYINPUT69), .A2(G237), .ZN(new_n187));
  NAND2_X1  g001(.A1(KEYINPUT69), .A2(G237), .ZN(new_n188));
  AOI21_X1  g002(.A(G953), .B1(new_n187), .B2(new_n188), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G210), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT27), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT26), .B(G101), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n190), .B(KEYINPUT27), .ZN(new_n195));
  INV_X1    g009(.A(new_n193), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(new_n197), .ZN(new_n198));
  OR2_X1    g012(.A1(KEYINPUT66), .A2(G116), .ZN(new_n199));
  NAND2_X1  g013(.A1(KEYINPUT66), .A2(G116), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(G119), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G116), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(G119), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n201), .A2(new_n204), .ZN(new_n205));
  XOR2_X1   g019(.A(KEYINPUT2), .B(G113), .Z(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT67), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  AND2_X1   g022(.A1(KEYINPUT66), .A2(G116), .ZN(new_n209));
  NOR2_X1   g023(.A1(KEYINPUT66), .A2(G116), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n203), .B1(new_n211), .B2(G119), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n213), .A3(new_n206), .ZN(new_n214));
  AOI22_X1  g028(.A1(new_n208), .A2(new_n214), .B1(new_n205), .B2(new_n207), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G143), .ZN(new_n217));
  INV_X1    g031(.A(G143), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G128), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n216), .A2(G143), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n217), .A2(new_n219), .A3(G128), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n222), .B(new_n225), .C1(new_n223), .C2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G131), .ZN(new_n228));
  INV_X1    g042(.A(G137), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(G134), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT11), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n232), .B1(G134), .B2(new_n229), .ZN(new_n233));
  INV_X1    g047(.A(G134), .ZN(new_n234));
  NOR3_X1   g048(.A1(new_n234), .A2(KEYINPUT11), .A3(G137), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n228), .B(new_n231), .C1(new_n233), .C2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT64), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n237), .B1(new_n229), .B2(G134), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n229), .A2(G134), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n234), .A2(KEYINPUT64), .A3(G137), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G131), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n227), .A2(new_n236), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(KEYINPUT0), .A2(G128), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n217), .A2(new_n219), .A3(new_n244), .ZN(new_n245));
  XOR2_X1   g059(.A(KEYINPUT0), .B(G128), .Z(new_n246));
  XNOR2_X1  g060(.A(G143), .B(G146), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT11), .B1(new_n234), .B2(G137), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n232), .A2(new_n229), .A3(G134), .ZN(new_n250));
  AOI211_X1 g064(.A(G131), .B(new_n230), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n250), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n228), .B1(new_n252), .B2(new_n231), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n248), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT68), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT68), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n256), .B(new_n248), .C1(new_n251), .C2(new_n253), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n243), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n198), .B1(new_n215), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n227), .A2(new_n236), .A3(new_n242), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n254), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n262), .A2(KEYINPUT30), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n252), .A2(new_n231), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G131), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(new_n236), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n256), .B1(new_n266), .B2(new_n248), .ZN(new_n267));
  INV_X1    g081(.A(new_n257), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n261), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n263), .B1(new_n269), .B2(KEYINPUT30), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n259), .B(new_n260), .C1(new_n270), .C2(new_n215), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n242), .A2(new_n236), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n266), .A2(new_n248), .B1(new_n273), .B2(new_n227), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT30), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n276), .B1(new_n258), .B2(new_n275), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n213), .B1(new_n212), .B2(new_n206), .ZN(new_n278));
  AND4_X1   g092(.A1(new_n213), .A2(new_n206), .A3(new_n201), .A4(new_n204), .ZN(new_n279));
  OAI22_X1  g093(.A1(new_n278), .A2(new_n279), .B1(new_n212), .B2(new_n206), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n260), .B1(new_n281), .B2(new_n259), .ZN(new_n282));
  OAI21_X1  g096(.A(KEYINPUT31), .B1(new_n272), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n259), .B1(new_n270), .B2(new_n215), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT31), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT71), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n287), .B1(new_n274), .B2(new_n215), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n215), .B(new_n261), .C1(new_n267), .C2(new_n268), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n262), .A2(KEYINPUT71), .A3(new_n280), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT28), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT72), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT72), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n291), .A2(new_n294), .A3(KEYINPUT28), .ZN(new_n295));
  AOI21_X1  g109(.A(KEYINPUT28), .B1(new_n274), .B2(new_n215), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n293), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n283), .A2(new_n286), .B1(new_n198), .B2(new_n298), .ZN(new_n299));
  NOR2_X1   g113(.A1(G472), .A2(G902), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NOR3_X1   g115(.A1(new_n299), .A2(KEYINPUT32), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT32), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n284), .A2(KEYINPUT70), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n285), .B1(new_n304), .B2(new_n271), .ZN(new_n305));
  INV_X1    g119(.A(new_n286), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n291), .A2(new_n294), .A3(KEYINPUT28), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n294), .B1(new_n291), .B2(KEYINPUT28), .ZN(new_n308));
  NOR3_X1   g122(.A1(new_n307), .A2(new_n308), .A3(new_n296), .ZN(new_n309));
  INV_X1    g123(.A(new_n198), .ZN(new_n310));
  OAI22_X1  g124(.A1(new_n305), .A2(new_n306), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n303), .B1(new_n311), .B2(new_n300), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n293), .A2(new_n310), .A3(new_n295), .A4(new_n297), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n281), .A2(new_n289), .ZN(new_n315));
  AOI21_X1  g129(.A(KEYINPUT29), .B1(new_n315), .B2(new_n198), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n289), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n255), .A2(new_n257), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n215), .B1(new_n319), .B2(new_n261), .ZN(new_n320));
  OAI21_X1  g134(.A(KEYINPUT28), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n310), .A2(KEYINPUT29), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n297), .A3(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G902), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n317), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n313), .B1(new_n327), .B2(G472), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n325), .B1(new_n314), .B2(new_n316), .ZN(new_n329));
  INV_X1    g143(.A(G472), .ZN(new_n330));
  NOR3_X1   g144(.A1(new_n329), .A2(KEYINPUT73), .A3(new_n330), .ZN(new_n331));
  OAI22_X1  g145(.A1(new_n302), .A2(new_n312), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT22), .B(G137), .ZN(new_n333));
  INV_X1    g147(.A(G953), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n334), .A2(G221), .A3(G234), .ZN(new_n335));
  XOR2_X1   g149(.A(new_n333), .B(new_n335), .Z(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G119), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G128), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n221), .A2(G119), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT74), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT74), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n339), .A2(new_n340), .A3(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT24), .B(G110), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n342), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT75), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n347), .B(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n340), .A2(KEYINPUT78), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT78), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(new_n221), .A3(G119), .ZN(new_n352));
  OAI22_X1  g166(.A1(new_n221), .A2(G119), .B1(KEYINPUT77), .B2(KEYINPUT23), .ZN(new_n353));
  AND2_X1   g167(.A1(KEYINPUT77), .A2(KEYINPUT23), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n350), .B(new_n352), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT76), .ZN(new_n356));
  NAND2_X1  g170(.A1(KEYINPUT23), .A2(G119), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n356), .B1(new_n357), .B2(G128), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n221), .A2(KEYINPUT76), .A3(KEYINPUT23), .A4(G119), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT16), .ZN(new_n362));
  INV_X1    g176(.A(G140), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(new_n363), .A3(G125), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(G125), .ZN(new_n365));
  INV_X1    g179(.A(G125), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G140), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n364), .B1(new_n368), .B2(new_n362), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n216), .ZN(new_n370));
  OAI211_X1 g184(.A(G146), .B(new_n364), .C1(new_n368), .C2(new_n362), .ZN(new_n371));
  AOI22_X1  g185(.A1(G110), .A2(new_n361), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n349), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n365), .A2(new_n367), .A3(new_n216), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  XOR2_X1   g189(.A(KEYINPUT79), .B(G110), .Z(new_n376));
  NAND4_X1  g190(.A1(new_n355), .A2(new_n360), .A3(KEYINPUT80), .A4(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n342), .A2(new_n344), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n345), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n355), .A2(new_n360), .A3(new_n376), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT80), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n375), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n337), .B1(new_n373), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n380), .A2(new_n383), .ZN(new_n386));
  INV_X1    g200(.A(new_n375), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n349), .A2(new_n372), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n389), .A3(new_n336), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n385), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G217), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n392), .B1(G234), .B2(new_n324), .ZN(new_n393));
  NOR3_X1   g207(.A1(new_n391), .A2(G902), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n385), .A2(new_n390), .A3(new_n324), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT25), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n385), .A2(new_n390), .A3(KEYINPUT25), .A4(new_n324), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n394), .B1(new_n399), .B2(new_n393), .ZN(new_n400));
  XNOR2_X1  g214(.A(G113), .B(G122), .ZN(new_n401));
  INV_X1    g215(.A(G104), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n401), .B(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n368), .A2(G146), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n374), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n189), .A2(G143), .A3(G214), .ZN(new_n407));
  AND2_X1   g221(.A1(KEYINPUT69), .A2(G237), .ZN(new_n408));
  NOR2_X1   g222(.A1(KEYINPUT69), .A2(G237), .ZN(new_n409));
  OAI211_X1 g223(.A(G214), .B(new_n334), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n218), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(KEYINPUT18), .A2(G131), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n406), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n410), .B(G143), .ZN(new_n416));
  OAI21_X1  g230(.A(KEYINPUT88), .B1(new_n416), .B2(new_n413), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT88), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n412), .A2(new_n418), .A3(new_n414), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n415), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n368), .B(KEYINPUT19), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n371), .B1(new_n421), .B2(G146), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n412), .A2(G131), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n407), .A2(new_n411), .A3(new_n228), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n404), .B1(new_n420), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n370), .A2(new_n371), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n228), .B1(new_n407), .B2(new_n411), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n427), .B1(KEYINPUT17), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT17), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n423), .A2(new_n430), .A3(new_n424), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n416), .A2(new_n413), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n418), .B1(new_n412), .B2(new_n414), .ZN(new_n434));
  AOI211_X1 g248(.A(KEYINPUT88), .B(new_n413), .C1(new_n407), .C2(new_n411), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n406), .B(new_n433), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n432), .A2(new_n436), .A3(new_n403), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n426), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(G475), .A2(G902), .ZN(new_n439));
  XOR2_X1   g253(.A(new_n439), .B(KEYINPUT89), .Z(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(KEYINPUT90), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT20), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n432), .A2(new_n436), .A3(new_n403), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n403), .B1(new_n432), .B2(new_n436), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n324), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(G475), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n440), .B1(new_n426), .B2(new_n437), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(KEYINPUT90), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(KEYINPUT20), .B1(new_n449), .B2(KEYINPUT90), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n444), .B(new_n448), .C1(new_n451), .C2(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n218), .A2(G128), .ZN(new_n454));
  OAI21_X1  g268(.A(G134), .B1(new_n454), .B2(KEYINPUT13), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n218), .A2(G128), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n221), .A2(G143), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n455), .A2(new_n458), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n199), .A2(G122), .A3(new_n200), .ZN(new_n461));
  XNOR2_X1  g275(.A(KEYINPUT82), .B(G107), .ZN(new_n462));
  OR2_X1    g276(.A1(new_n202), .A2(G122), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n462), .B1(new_n461), .B2(new_n463), .ZN(new_n465));
  OAI22_X1  g279(.A1(new_n459), .A2(new_n460), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n456), .A2(new_n457), .A3(G134), .ZN(new_n468));
  AOI21_X1  g282(.A(G134), .B1(new_n456), .B2(new_n457), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT14), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n461), .A2(new_n471), .A3(new_n463), .ZN(new_n472));
  OAI21_X1  g286(.A(G107), .B1(new_n461), .B2(new_n471), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n467), .B(new_n470), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(KEYINPUT9), .B(G234), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n475), .B(KEYINPUT81), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n334), .A2(G217), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n466), .A2(new_n474), .A3(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT91), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n466), .A2(new_n474), .ZN(new_n482));
  INV_X1    g296(.A(new_n478), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n466), .A2(new_n474), .A3(new_n478), .A4(KEYINPUT91), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n481), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n324), .ZN(new_n487));
  INV_X1    g301(.A(G478), .ZN(new_n488));
  OR2_X1    g302(.A1(new_n488), .A2(KEYINPUT15), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n487), .B(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n453), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(G234), .A2(G237), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n493), .A2(G902), .A3(G953), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(KEYINPUT21), .B(G898), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n334), .A2(G952), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n495), .A2(new_n496), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n492), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(G214), .B1(G237), .B2(G902), .ZN(new_n501));
  INV_X1    g315(.A(G107), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT82), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT82), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G107), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT3), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n503), .A2(new_n505), .A3(new_n506), .A4(G104), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n506), .B1(new_n502), .B2(G104), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n502), .A2(G104), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT4), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n511), .A2(new_n512), .A3(G101), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n511), .A2(G101), .ZN(new_n514));
  INV_X1    g328(.A(G101), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n507), .A2(new_n510), .A3(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n514), .A2(KEYINPUT4), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n280), .A2(new_n513), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n212), .A2(KEYINPUT5), .ZN(new_n519));
  INV_X1    g333(.A(G113), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT5), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n520), .B1(new_n203), .B2(new_n521), .ZN(new_n522));
  AOI22_X1  g336(.A1(new_n208), .A2(new_n214), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT83), .ZN(new_n524));
  AOI21_X1  g338(.A(G104), .B1(new_n503), .B2(new_n505), .ZN(new_n525));
  INV_X1    g339(.A(new_n509), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n524), .B(G101), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n516), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n509), .B1(new_n462), .B2(G104), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n524), .B1(new_n529), .B2(G101), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n523), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g346(.A(G110), .B(G122), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n518), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G224), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n535), .A2(G953), .ZN(new_n536));
  XOR2_X1   g350(.A(KEYINPUT65), .B(KEYINPUT1), .Z(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(G128), .A3(new_n247), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n538), .A2(new_n366), .A3(new_n225), .A4(new_n222), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT86), .ZN(new_n540));
  OAI22_X1  g354(.A1(new_n539), .A2(new_n540), .B1(new_n366), .B2(new_n248), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n539), .A2(new_n540), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n536), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT7), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n544), .B1(new_n541), .B2(new_n542), .ZN(new_n545));
  AND3_X1   g359(.A1(new_n534), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n503), .A2(new_n505), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n526), .B1(new_n547), .B2(new_n402), .ZN(new_n548));
  OAI21_X1  g362(.A(KEYINPUT83), .B1(new_n548), .B2(new_n515), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n549), .A2(new_n516), .A3(new_n527), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT87), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n523), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  XOR2_X1   g366(.A(new_n533), .B(KEYINPUT8), .Z(new_n553));
  NOR2_X1   g367(.A1(new_n550), .A2(new_n551), .ZN(new_n554));
  INV_X1    g368(.A(new_n523), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR3_X1   g370(.A1(new_n541), .A2(new_n542), .A3(new_n536), .ZN(new_n557));
  AOI22_X1  g371(.A1(new_n552), .A2(new_n556), .B1(new_n557), .B2(KEYINPUT7), .ZN(new_n558));
  AOI21_X1  g372(.A(G902), .B1(new_n546), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n518), .A2(new_n532), .ZN(new_n560));
  INV_X1    g374(.A(new_n533), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT6), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n563), .A2(KEYINPUT85), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n562), .A2(new_n534), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n557), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n543), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n560), .B(new_n561), .C1(KEYINPUT85), .C2(new_n563), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n565), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(G210), .B1(G237), .B2(G902), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n559), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n570), .B1(new_n559), .B2(new_n569), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n501), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(G469), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n531), .A2(KEYINPUT10), .A3(new_n227), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n218), .A2(KEYINPUT1), .A3(G146), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n222), .B(new_n576), .C1(new_n223), .C2(new_n226), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n549), .A2(new_n516), .A3(new_n577), .A4(new_n527), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT10), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n517), .A2(new_n248), .A3(new_n513), .ZN(new_n581));
  INV_X1    g395(.A(new_n266), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n575), .A2(new_n580), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(G110), .B(G140), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n334), .A2(G227), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n584), .B(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n227), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n589), .B1(new_n528), .B2(new_n530), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n590), .A2(KEYINPUT84), .A3(new_n578), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT84), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n550), .A2(new_n592), .A3(new_n589), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n591), .A2(KEYINPUT12), .A3(new_n266), .A4(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n591), .A2(new_n266), .A3(new_n593), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT12), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n588), .B1(new_n594), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n575), .A2(new_n580), .A3(new_n581), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n266), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n587), .B1(new_n600), .B2(new_n583), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n574), .B(new_n324), .C1(new_n598), .C2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n600), .A2(new_n587), .A3(new_n583), .ZN(new_n603));
  INV_X1    g417(.A(new_n583), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n604), .B1(new_n597), .B2(new_n594), .ZN(new_n605));
  OAI211_X1 g419(.A(G469), .B(new_n603), .C1(new_n605), .C2(new_n587), .ZN(new_n606));
  NAND2_X1  g420(.A1(G469), .A2(G902), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n602), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(G221), .B1(new_n476), .B2(G902), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n500), .A2(new_n573), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n332), .A2(new_n400), .A3(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(G101), .ZN(G3));
  AND3_X1   g427(.A1(new_n608), .A2(new_n400), .A3(new_n609), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n311), .A2(new_n300), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n283), .A2(new_n286), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n298), .A2(new_n198), .ZN(new_n617));
  AOI21_X1  g431(.A(G902), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  OAI211_X1 g432(.A(new_n614), .B(new_n615), .C1(new_n618), .C2(new_n330), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT92), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n311), .A2(new_n324), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(G472), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n623), .A2(KEYINPUT92), .A3(new_n615), .A4(new_n614), .ZN(new_n624));
  INV_X1    g438(.A(new_n501), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n559), .A2(new_n569), .ZN(new_n626));
  INV_X1    g440(.A(new_n570), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n559), .A2(new_n569), .A3(new_n570), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n625), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n499), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n438), .A2(new_n441), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT90), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n634), .A2(KEYINPUT20), .A3(new_n450), .ZN(new_n635));
  AOI22_X1  g449(.A1(new_n442), .A2(new_n443), .B1(G475), .B2(new_n447), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n324), .A2(G478), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT33), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n482), .B2(new_n483), .ZN(new_n639));
  AOI221_X4 g453(.A(new_n637), .B1(new_n639), .B2(new_n479), .C1(new_n486), .C2(new_n638), .ZN(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT93), .B(G478), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n642), .B1(new_n486), .B2(new_n324), .ZN(new_n643));
  OAI21_X1  g457(.A(KEYINPUT94), .B1(new_n640), .B2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n643), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT94), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n486), .A2(new_n638), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n639), .A2(new_n479), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n645), .B(new_n646), .C1(new_n649), .C2(new_n637), .ZN(new_n650));
  AOI22_X1  g464(.A1(new_n635), .A2(new_n636), .B1(new_n644), .B2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n631), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n621), .A2(new_n624), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT34), .B(G104), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT95), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n654), .B(new_n656), .ZN(G6));
  INV_X1    g471(.A(new_n453), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n491), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n631), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n621), .A2(new_n624), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT35), .B(G107), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G9));
  NAND2_X1  g477(.A1(new_n388), .A2(new_n389), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT96), .ZN(new_n665));
  OR2_X1    g479(.A1(new_n337), .A2(KEYINPUT36), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n393), .A2(G902), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n399), .A2(new_n393), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n611), .A2(new_n615), .A3(new_n623), .A4(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT37), .B(G110), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(KEYINPUT97), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n672), .B(new_n674), .ZN(G12));
  NAND2_X1  g489(.A1(new_n497), .A2(new_n493), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT98), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(G900), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n678), .B1(new_n679), .B2(new_n495), .ZN(new_n680));
  NOR4_X1   g494(.A1(new_n659), .A2(new_n610), .A3(new_n573), .A4(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n332), .A2(new_n681), .A3(new_n671), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G128), .ZN(G30));
  NAND2_X1  g497(.A1(new_n453), .A2(new_n491), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n671), .A2(new_n625), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT99), .ZN(new_n686));
  OAI21_X1  g500(.A(KEYINPUT32), .B1(new_n299), .B2(new_n301), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n311), .A2(new_n303), .A3(new_n300), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n272), .A2(new_n282), .ZN(new_n690));
  OR2_X1    g504(.A1(new_n318), .A2(new_n320), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n690), .B1(new_n310), .B2(new_n692), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n693), .A2(new_n324), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n689), .B1(new_n330), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n628), .A2(new_n629), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT38), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n686), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT100), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  INV_X1    g515(.A(new_n610), .ZN(new_n702));
  XOR2_X1   g516(.A(new_n680), .B(KEYINPUT39), .Z(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g518(.A(new_n704), .B(KEYINPUT40), .Z(new_n705));
  NAND3_X1  g519(.A1(new_n700), .A2(new_n701), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G143), .ZN(G45));
  NAND2_X1  g521(.A1(new_n644), .A2(new_n650), .ZN(new_n708));
  INV_X1    g522(.A(new_n680), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n453), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g524(.A(KEYINPUT101), .B1(new_n710), .B2(new_n573), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT101), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n630), .A2(new_n712), .A3(new_n651), .A4(new_n709), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n332), .A2(new_n702), .A3(new_n671), .A4(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT102), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n669), .A2(new_n670), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n327), .A2(new_n313), .A3(G472), .ZN(new_n719));
  OAI21_X1  g533(.A(KEYINPUT73), .B1(new_n329), .B2(new_n330), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n718), .B1(new_n689), .B2(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n722), .A2(KEYINPUT102), .A3(new_n702), .A4(new_n714), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n717), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G146), .ZN(G48));
  OAI21_X1  g539(.A(new_n324), .B1(new_n598), .B2(new_n601), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(G469), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT103), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n727), .A2(new_n728), .A3(new_n602), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n726), .A2(KEYINPUT103), .A3(G469), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n609), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n332), .A2(new_n734), .A3(new_n400), .A4(new_n653), .ZN(new_n735));
  XNOR2_X1  g549(.A(KEYINPUT41), .B(G113), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G15));
  NAND4_X1  g551(.A1(new_n332), .A2(new_n734), .A3(new_n400), .A4(new_n660), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G116), .ZN(G18));
  INV_X1    g553(.A(new_n500), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n731), .A2(new_n630), .A3(new_n609), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n332), .A2(new_n740), .A3(new_n671), .A4(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G119), .ZN(G21));
  AND2_X1   g557(.A1(new_n321), .A2(new_n297), .ZN(new_n744));
  OAI22_X1  g558(.A1(new_n305), .A2(new_n306), .B1(new_n310), .B2(new_n744), .ZN(new_n745));
  AOI22_X1  g559(.A1(new_n622), .A2(G472), .B1(new_n300), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n631), .A2(new_n684), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n734), .A2(new_n746), .A3(new_n747), .A4(new_n400), .ZN(new_n748));
  XNOR2_X1  g562(.A(KEYINPUT104), .B(G122), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(G24));
  INV_X1    g564(.A(new_n710), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n741), .A2(new_n746), .A3(new_n671), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G125), .ZN(G27));
  NAND4_X1  g567(.A1(new_n628), .A2(new_n501), .A3(new_n629), .A4(new_n609), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n607), .B(KEYINPUT105), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n602), .A2(new_n606), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(KEYINPUT106), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT106), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n602), .A2(new_n606), .A3(new_n758), .A4(new_n755), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n754), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n332), .A2(new_n400), .A3(new_n751), .A4(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT42), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g577(.A(KEYINPUT107), .B1(new_n302), .B2(new_n312), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT107), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n687), .A2(new_n688), .A3(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n764), .A2(new_n721), .A3(new_n766), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n760), .A2(KEYINPUT42), .A3(new_n751), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(new_n400), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n763), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT108), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n763), .A2(new_n769), .A3(KEYINPUT108), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(new_n228), .ZN(G33));
  NOR2_X1   g589(.A1(new_n659), .A2(new_n680), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n332), .A2(new_n400), .A3(new_n776), .A4(new_n760), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G134), .ZN(G36));
  OAI21_X1  g592(.A(new_n603), .B1(new_n605), .B2(new_n587), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT45), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n574), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n781), .B1(new_n780), .B2(new_n779), .ZN(new_n782));
  XOR2_X1   g596(.A(new_n782), .B(KEYINPUT109), .Z(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(KEYINPUT46), .A3(new_n755), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n602), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n785), .A2(KEYINPUT110), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT46), .B1(new_n783), .B2(new_n755), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT110), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n788), .B1(new_n784), .B2(new_n602), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n786), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n790), .A2(new_n733), .ZN(new_n791));
  INV_X1    g605(.A(new_n708), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(new_n453), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(KEYINPUT43), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n623), .A2(new_n615), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(new_n795), .A3(new_n671), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT44), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n696), .A2(new_n625), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n800), .B1(new_n796), .B2(new_n797), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n791), .A2(new_n703), .A3(new_n798), .A4(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G137), .ZN(G39));
  INV_X1    g617(.A(KEYINPUT47), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n804), .B1(new_n790), .B2(new_n733), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n789), .A2(new_n787), .ZN(new_n806));
  OAI211_X1 g620(.A(KEYINPUT47), .B(new_n609), .C1(new_n806), .C2(new_n786), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NOR4_X1   g622(.A1(new_n332), .A2(new_n400), .A3(new_n710), .A4(new_n800), .ZN(new_n809));
  XOR2_X1   g623(.A(new_n809), .B(KEYINPUT111), .Z(new_n810));
  NAND2_X1  g624(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(KEYINPUT112), .B(G140), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n811), .B(new_n812), .ZN(G42));
  AND4_X1   g627(.A1(new_n678), .A2(new_n794), .A3(new_n734), .A4(new_n799), .ZN(new_n814));
  XOR2_X1   g628(.A(new_n814), .B(KEYINPUT117), .Z(new_n815));
  NAND2_X1  g629(.A1(new_n767), .A2(new_n400), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(KEYINPUT48), .ZN(new_n818));
  INV_X1    g632(.A(new_n741), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n794), .A2(new_n400), .A3(new_n678), .A4(new_n746), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n689), .B(new_n400), .C1(new_n330), .C2(new_n694), .ZN(new_n821));
  INV_X1    g635(.A(new_n734), .ZN(new_n822));
  OR4_X1    g636(.A1(new_n676), .A2(new_n821), .A3(new_n822), .A4(new_n800), .ZN(new_n823));
  OAI221_X1 g637(.A(new_n497), .B1(new_n819), .B2(new_n820), .C1(new_n823), .C2(new_n652), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n818), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n746), .A2(new_n671), .ZN(new_n826));
  OR2_X1    g640(.A1(new_n815), .A2(new_n826), .ZN(new_n827));
  NOR4_X1   g641(.A1(new_n820), .A2(new_n501), .A3(new_n697), .A4(new_n822), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(KEYINPUT50), .ZN(new_n829));
  OR3_X1    g643(.A1(new_n823), .A2(new_n453), .A3(new_n708), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n827), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n805), .B(new_n807), .C1(new_n609), .C2(new_n732), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n820), .A2(new_n800), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n825), .B1(new_n834), .B2(KEYINPUT51), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n827), .A2(KEYINPUT51), .A3(new_n829), .A4(new_n830), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n832), .A2(KEYINPUT118), .ZN(new_n837));
  INV_X1    g651(.A(new_n833), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n838), .B1(new_n832), .B2(KEYINPUT118), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n836), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  OR2_X1    g654(.A1(new_n835), .A2(new_n840), .ZN(new_n841));
  OR3_X1    g655(.A1(new_n453), .A2(KEYINPUT113), .A3(new_n490), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT113), .B1(new_n453), .B2(new_n490), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n844), .A2(new_n631), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n621), .A2(new_n624), .A3(new_n845), .ZN(new_n846));
  AND4_X1   g660(.A1(new_n612), .A2(new_n654), .A3(new_n846), .A4(new_n672), .ZN(new_n847));
  AND4_X1   g661(.A1(new_n735), .A2(new_n738), .A3(new_n742), .A4(new_n748), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n799), .A2(new_n492), .A3(new_n709), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n332), .A2(new_n702), .A3(new_n671), .A4(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n746), .A2(new_n671), .A3(new_n751), .A4(new_n760), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n777), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n847), .A2(new_n848), .A3(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(KEYINPUT114), .B1(new_n774), .B2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n654), .A2(new_n846), .A3(new_n612), .A4(new_n672), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n735), .A2(new_n738), .A3(new_n742), .A4(new_n748), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n856), .A2(new_n857), .A3(new_n852), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT114), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n858), .A2(new_n859), .A3(new_n772), .A4(new_n773), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n855), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n682), .A2(new_n752), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n757), .A2(new_n759), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n630), .A2(new_n491), .A3(new_n453), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n709), .A2(new_n609), .ZN(new_n866));
  NOR4_X1   g680(.A1(new_n864), .A2(new_n865), .A3(new_n671), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n695), .ZN(new_n868));
  AOI211_X1 g682(.A(new_n610), .B(new_n718), .C1(new_n689), .C2(new_n721), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT102), .B1(new_n869), .B2(new_n714), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n715), .A2(new_n716), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n863), .B(new_n868), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  XNOR2_X1  g686(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT53), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n862), .B1(new_n717), .B2(new_n723), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT52), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n877), .A2(new_n878), .A3(new_n868), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n875), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  AND4_X1   g694(.A1(new_n878), .A2(new_n724), .A3(new_n863), .A4(new_n868), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n878), .B1(new_n877), .B2(new_n868), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n855), .A2(new_n883), .A3(new_n860), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  OAI221_X1 g699(.A(KEYINPUT54), .B1(new_n861), .B2(new_n880), .C1(new_n885), .C2(new_n876), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n884), .A2(new_n876), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n876), .B1(new_n763), .B2(new_n769), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n875), .A2(new_n858), .A3(new_n879), .A4(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT116), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AND4_X1   g705(.A1(new_n847), .A2(new_n888), .A3(new_n848), .A4(new_n853), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n892), .A2(KEYINPUT116), .A3(new_n879), .A4(new_n875), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT54), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n887), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n886), .A2(new_n896), .ZN(new_n897));
  OAI22_X1  g711(.A1(new_n841), .A2(new_n897), .B1(G952), .B2(G953), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n731), .B(KEYINPUT49), .Z(new_n899));
  NAND3_X1  g713(.A1(new_n793), .A2(new_n501), .A3(new_n609), .ZN(new_n900));
  OR4_X1    g714(.A1(new_n697), .A2(new_n899), .A3(new_n821), .A4(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n898), .A2(new_n901), .ZN(G75));
  INV_X1    g716(.A(KEYINPUT120), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n887), .A2(new_n894), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT119), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n904), .A2(new_n905), .A3(G210), .A4(G902), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n565), .A2(new_n568), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n907), .B(new_n567), .Z(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT55), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n909), .A2(KEYINPUT56), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n324), .B1(new_n887), .B2(new_n894), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n905), .B1(new_n912), .B2(G210), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n334), .A2(G952), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT56), .B1(new_n912), .B2(G210), .ZN(new_n917));
  INV_X1    g731(.A(new_n909), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n903), .B1(new_n914), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n904), .A2(G210), .A3(G902), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT56), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n915), .B1(new_n923), .B2(new_n909), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n921), .A2(KEYINPUT119), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n925), .A2(new_n906), .A3(new_n910), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n924), .A2(KEYINPUT120), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n920), .A2(new_n927), .ZN(G51));
  INV_X1    g742(.A(KEYINPUT121), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n896), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n887), .A2(new_n894), .A3(KEYINPUT121), .A4(new_n895), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n904), .A2(KEYINPUT54), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n755), .B(KEYINPUT57), .Z(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OR2_X1    g749(.A1(new_n598), .A2(new_n601), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(new_n912), .ZN(new_n938));
  OR2_X1    g752(.A1(new_n938), .A2(new_n783), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n915), .B1(new_n937), .B2(new_n939), .ZN(G54));
  NAND2_X1  g754(.A1(KEYINPUT58), .A2(G475), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT122), .Z(new_n942));
  NAND2_X1  g756(.A1(new_n912), .A2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n438), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n916), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT123), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n946), .B1(new_n943), .B2(new_n944), .ZN(new_n947));
  AOI211_X1 g761(.A(KEYINPUT123), .B(new_n438), .C1(new_n912), .C2(new_n942), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n945), .A2(new_n947), .A3(new_n948), .ZN(G60));
  XOR2_X1   g763(.A(KEYINPUT124), .B(KEYINPUT59), .Z(new_n950));
  NOR2_X1   g764(.A1(new_n488), .A2(new_n324), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n952), .B1(new_n886), .B2(new_n896), .ZN(new_n953));
  INV_X1    g767(.A(new_n649), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n916), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n649), .A2(new_n952), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n955), .B1(new_n933), .B2(new_n956), .ZN(G63));
  NAND2_X1  g771(.A1(G217), .A2(G902), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT125), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT60), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n904), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n667), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT126), .ZN(new_n963));
  AOI21_X1  g777(.A(KEYINPUT61), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n915), .B1(new_n961), .B2(new_n667), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n904), .A2(new_n960), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n391), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n964), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(KEYINPUT126), .B1(new_n961), .B2(new_n667), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n967), .B(new_n965), .C1(new_n970), .C2(KEYINPUT61), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n969), .A2(new_n971), .ZN(G66));
  NAND2_X1  g786(.A1(new_n847), .A2(new_n848), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n334), .ZN(new_n974));
  OAI21_X1  g788(.A(G953), .B1(new_n496), .B2(new_n535), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n907), .B1(G898), .B2(new_n334), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n976), .B(new_n977), .ZN(G69));
  INV_X1    g792(.A(new_n811), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n816), .A2(new_n865), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n791), .A2(new_n703), .A3(new_n980), .ZN(new_n981));
  AND4_X1   g795(.A1(new_n772), .A2(new_n773), .A3(new_n777), .A4(new_n877), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n802), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n979), .A2(new_n983), .A3(G953), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n679), .A2(new_n334), .ZN(new_n985));
  OR2_X1    g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(G227), .A2(G900), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n270), .B(new_n421), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n986), .A2(G953), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n988), .B1(new_n984), .B2(new_n985), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n987), .A2(G953), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n706), .A2(new_n877), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(KEYINPUT62), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT127), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n993), .B(new_n994), .ZN(new_n995));
  OR2_X1    g809(.A1(new_n992), .A2(KEYINPUT62), .ZN(new_n996));
  AOI211_X1 g810(.A(new_n800), .B(new_n704), .C1(new_n652), .C2(new_n844), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n997), .A2(new_n332), .A3(new_n400), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n996), .A2(new_n811), .A3(new_n802), .A4(new_n998), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n995), .A2(new_n999), .ZN(new_n1000));
  OR2_X1    g814(.A1(new_n988), .A2(G953), .ZN(new_n1001));
  OAI211_X1 g815(.A(new_n990), .B(new_n991), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n989), .A2(new_n1002), .ZN(G72));
  AOI21_X1  g817(.A(new_n198), .B1(new_n281), .B2(new_n289), .ZN(new_n1004));
  NOR3_X1   g818(.A1(new_n995), .A2(new_n999), .A3(new_n973), .ZN(new_n1005));
  NAND2_X1  g819(.A1(G472), .A2(G902), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1006), .B(KEYINPUT63), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1004), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n315), .A2(new_n310), .ZN(new_n1009));
  NOR3_X1   g823(.A1(new_n979), .A2(new_n983), .A3(new_n973), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1009), .B1(new_n1010), .B2(new_n1007), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n315), .A2(new_n198), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1007), .B1(new_n690), .B2(new_n1012), .ZN(new_n1013));
  OAI221_X1 g827(.A(new_n1013), .B1(new_n861), .B2(new_n880), .C1(new_n885), .C2(new_n876), .ZN(new_n1014));
  AND4_X1   g828(.A1(new_n916), .A2(new_n1008), .A3(new_n1011), .A4(new_n1014), .ZN(G57));
endmodule


