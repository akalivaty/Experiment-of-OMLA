//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 0 1 0 1 0 1 0 0 0 0 0 0 1 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n577, new_n578, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n599, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n635, new_n638, new_n640,
    new_n641, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1174, new_n1175, new_n1176;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  INV_X1    g022(.A(G567), .ZN(new_n448));
  NOR2_X1   g023(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT65), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT66), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n453), .A2(new_n458), .B1(new_n448), .B2(new_n454), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT67), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT68), .Z(G319));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT69), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n467), .B1(new_n463), .B2(G2105), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n469), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  AOI22_X1  g046(.A1(G137), .A2(new_n466), .B1(new_n471), .B2(G101), .ZN(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n473), .B1(new_n464), .B2(new_n465), .ZN(new_n474));
  AND2_X1   g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  OAI21_X1  g050(.A(G2105), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT70), .ZN(G160));
  AND2_X1   g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NOR2_X1   g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(new_n469), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  XOR2_X1   g058(.A(new_n483), .B(KEYINPUT72), .Z(new_n484));
  XNOR2_X1  g059(.A(new_n466), .B(KEYINPUT71), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n484), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n492), .B1(new_n479), .B2(new_n480), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT73), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g070(.A(KEYINPUT3), .B(G2104), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n496), .A2(KEYINPUT73), .A3(new_n492), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n495), .A2(KEYINPUT4), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n493), .A2(new_n494), .A3(new_n499), .ZN(new_n500));
  OAI211_X1 g075(.A(G126), .B(G2105), .C1(new_n479), .C2(new_n480), .ZN(new_n501));
  OR2_X1    g076(.A1(G102), .A2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G2105), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n502), .A2(new_n504), .A3(G2104), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n498), .A2(new_n500), .A3(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT74), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(KEYINPUT74), .A2(KEYINPUT5), .A3(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n515), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n517));
  AND2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n510), .A2(new_n516), .B1(new_n517), .B2(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  INV_X1    g097(.A(G543), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT6), .B(G651), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT76), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OR2_X1    g101(.A1(KEYINPUT6), .A2(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n527), .A2(KEYINPUT76), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G51), .ZN(new_n532));
  AND3_X1   g107(.A1(KEYINPUT74), .A2(KEYINPUT5), .A3(G543), .ZN(new_n533));
  AOI21_X1  g108(.A(KEYINPUT5), .B1(KEYINPUT74), .B2(G543), .ZN(new_n534));
  OAI21_X1  g109(.A(KEYINPUT75), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT75), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n513), .A2(new_n536), .A3(new_n514), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n538), .A2(G63), .A3(G651), .ZN(new_n539));
  XOR2_X1   g114(.A(KEYINPUT77), .B(KEYINPUT7), .Z(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n540), .B(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n533), .A2(new_n534), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n520), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G89), .ZN(new_n545));
  NAND4_X1  g120(.A1(new_n532), .A2(new_n539), .A3(new_n542), .A4(new_n545), .ZN(G286));
  INV_X1    g121(.A(G286), .ZN(G168));
  NAND2_X1  g122(.A1(new_n538), .A2(G64), .ZN(new_n548));
  NAND2_X1  g123(.A1(G77), .A2(G543), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n510), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n544), .A2(G90), .ZN(new_n551));
  XOR2_X1   g126(.A(KEYINPUT78), .B(G52), .Z(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n530), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(G171));
  OAI21_X1  g129(.A(new_n525), .B1(new_n518), .B2(new_n519), .ZN(new_n555));
  NAND4_X1  g130(.A1(new_n529), .A2(new_n555), .A3(G43), .A4(G543), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n515), .A2(G81), .A3(new_n524), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(KEYINPUT79), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT79), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n556), .A2(new_n560), .A3(new_n557), .ZN(new_n561));
  NAND2_X1  g136(.A1(G68), .A2(G543), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n535), .A2(new_n537), .ZN(new_n563));
  INV_X1    g138(.A(G56), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n559), .A2(new_n561), .B1(G651), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT80), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n565), .A2(G651), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n560), .B1(new_n556), .B2(new_n557), .ZN(new_n570));
  AND3_X1   g145(.A1(new_n556), .A2(new_n560), .A3(new_n557), .ZN(new_n571));
  OAI211_X1 g146(.A(new_n569), .B(new_n567), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G860), .ZN(G153));
  NAND4_X1  g150(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g151(.A1(G1), .A2(G3), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT8), .ZN(new_n578));
  NAND4_X1  g153(.A1(G319), .A2(G483), .A3(G661), .A4(new_n578), .ZN(G188));
  INV_X1    g154(.A(G78), .ZN(new_n580));
  OR3_X1    g155(.A1(new_n580), .A2(new_n523), .A3(KEYINPUT81), .ZN(new_n581));
  OAI21_X1  g156(.A(KEYINPUT81), .B1(new_n580), .B2(new_n523), .ZN(new_n582));
  XNOR2_X1  g157(.A(KEYINPUT82), .B(G65), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n581), .B(new_n582), .C1(new_n543), .C2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(G651), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n529), .A2(new_n555), .A3(G53), .A4(G543), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT9), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n526), .A2(KEYINPUT9), .A3(G53), .A4(new_n529), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n544), .A2(G91), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n585), .A2(new_n588), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(KEYINPUT83), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n584), .A2(G651), .B1(new_n544), .B2(G91), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT83), .ZN(new_n594));
  NAND4_X1  g169(.A1(new_n593), .A2(new_n594), .A3(new_n588), .A4(new_n589), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G299));
  INV_X1    g172(.A(G171), .ZN(G301));
  NAND3_X1  g173(.A1(new_n515), .A2(G87), .A3(new_n524), .ZN(new_n599));
  NAND4_X1  g174(.A1(new_n529), .A2(new_n555), .A3(G49), .A4(G543), .ZN(new_n600));
  AOI21_X1  g175(.A(G74), .B1(new_n535), .B2(new_n537), .ZN(new_n601));
  OAI211_X1 g176(.A(new_n599), .B(new_n600), .C1(new_n601), .C2(new_n510), .ZN(G288));
  NAND2_X1  g177(.A1(G73), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G61), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n543), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(G651), .ZN(new_n606));
  NAND2_X1  g181(.A1(G48), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G86), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n543), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(new_n524), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n606), .A2(new_n610), .ZN(G305));
  NAND2_X1  g186(.A1(new_n538), .A2(G60), .ZN(new_n612));
  NAND2_X1  g187(.A1(G72), .A2(G543), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n510), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(G47), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n515), .A2(new_n524), .ZN(new_n616));
  XNOR2_X1  g191(.A(KEYINPUT84), .B(G85), .ZN(new_n617));
  OAI22_X1  g192(.A1(new_n530), .A2(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(G290));
  NAND2_X1  g195(.A1(G301), .A2(G868), .ZN(new_n621));
  NAND2_X1  g196(.A1(G79), .A2(G543), .ZN(new_n622));
  INV_X1    g197(.A(G66), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n543), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G651), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n526), .A2(G54), .A3(new_n529), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(G92), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n616), .A2(new_n628), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n629), .A2(KEYINPUT10), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(KEYINPUT10), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n627), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n621), .B1(G868), .B2(new_n632), .ZN(G321));
  XOR2_X1   g208(.A(G321), .B(KEYINPUT85), .Z(G284));
  NAND2_X1  g209(.A1(G286), .A2(G868), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(new_n596), .B2(G868), .ZN(G297));
  XOR2_X1   g211(.A(G297), .B(KEYINPUT86), .Z(G280));
  INV_X1    g212(.A(G559), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n632), .B1(new_n638), .B2(G860), .ZN(G148));
  NAND2_X1  g214(.A1(new_n632), .A2(new_n638), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(G868), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(new_n574), .B2(G868), .ZN(G323));
  XNOR2_X1  g217(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g218(.A1(new_n485), .A2(G135), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n482), .A2(G123), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n469), .A2(G111), .ZN(new_n646));
  OAI21_X1  g221(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n647));
  OAI211_X1 g222(.A(new_n644), .B(new_n645), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT88), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2096), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n471), .A2(new_n496), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT12), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT13), .ZN(new_n653));
  XOR2_X1   g228(.A(KEYINPUT87), .B(G2100), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n650), .A2(new_n655), .ZN(G156));
  XOR2_X1   g231(.A(G2451), .B(G2454), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT16), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1341), .B(G1348), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT89), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n658), .B(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT14), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2427), .B(G2438), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2430), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT15), .B(G2435), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n666), .B1(new_n665), .B2(new_n664), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n661), .B(new_n667), .Z(new_n668));
  XNOR2_X1  g243(.A(G2443), .B(G2446), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  AND3_X1   g246(.A1(new_n670), .A2(G14), .A3(new_n671), .ZN(G401));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  XNOR2_X1  g248(.A(G2067), .B(G2678), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(KEYINPUT18), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2072), .B(G2078), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G2096), .B(G2100), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT90), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n678), .B(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT18), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n675), .A2(KEYINPUT17), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n673), .A2(new_n674), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n682), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n681), .B(new_n685), .Z(G227));
  XOR2_X1   g261(.A(G1971), .B(G1976), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1956), .B(G2474), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1961), .B(G1966), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n689), .A2(new_n690), .ZN(new_n693));
  NOR3_X1   g268(.A1(new_n688), .A2(new_n693), .A3(new_n691), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n688), .A2(new_n693), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT91), .B(KEYINPUT20), .Z(new_n696));
  AOI211_X1 g271(.A(new_n692), .B(new_n694), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(new_n695), .B2(new_n696), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT92), .Z(new_n699));
  XNOR2_X1  g274(.A(G1991), .B(G1996), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n699), .B(new_n704), .ZN(G229));
  INV_X1    g280(.A(G16), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G24), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(new_n619), .B2(new_n706), .ZN(new_n708));
  INV_X1    g283(.A(G1986), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n485), .A2(G131), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n482), .A2(G119), .ZN(new_n712));
  NOR2_X1   g287(.A1(G95), .A2(G2105), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT93), .ZN(new_n714));
  OAI21_X1  g289(.A(G2104), .B1(new_n469), .B2(G107), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n711), .B(new_n712), .C1(new_n714), .C2(new_n715), .ZN(new_n716));
  MUX2_X1   g291(.A(G25), .B(new_n716), .S(G29), .Z(new_n717));
  XOR2_X1   g292(.A(KEYINPUT35), .B(G1991), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  MUX2_X1   g294(.A(G6), .B(G305), .S(G16), .Z(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT32), .ZN(new_n721));
  INV_X1    g296(.A(G1981), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G288), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n724), .A2(new_n706), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(new_n706), .B2(G23), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT33), .B(G1976), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n706), .A2(G22), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G166), .B2(new_n706), .ZN(new_n730));
  INV_X1    g305(.A(G1971), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n726), .A2(new_n727), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n723), .A2(new_n728), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n710), .B(new_n719), .C1(new_n734), .C2(KEYINPUT34), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT94), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n734), .A2(KEYINPUT34), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT36), .ZN(new_n739));
  INV_X1    g314(.A(G29), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G35), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G162), .B2(new_n740), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT29), .Z(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G2090), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT30), .B(G28), .ZN(new_n745));
  OR2_X1    g320(.A1(KEYINPUT31), .A2(G11), .ZN(new_n746));
  NAND2_X1  g321(.A1(KEYINPUT31), .A2(G11), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n745), .A2(new_n740), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n482), .A2(G129), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n471), .A2(G105), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT26), .Z(new_n752));
  NAND3_X1  g327(.A1(new_n749), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n485), .B2(G141), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n754), .A2(new_n740), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n740), .B2(G32), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT27), .B(G1996), .ZN(new_n757));
  OAI221_X1 g332(.A(new_n748), .B1(new_n740), .B2(new_n648), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(G164), .A2(G29), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G27), .B2(G29), .ZN(new_n760));
  INV_X1    g335(.A(G2078), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n756), .A2(new_n757), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n761), .B2(new_n760), .ZN(new_n763));
  INV_X1    g338(.A(G1348), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n632), .A2(G16), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G4), .B2(G16), .ZN(new_n766));
  AOI211_X1 g341(.A(new_n758), .B(new_n763), .C1(new_n764), .C2(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(G34), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n768), .A2(KEYINPUT24), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n768), .A2(KEYINPUT24), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n740), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G160), .B2(new_n740), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G2084), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n740), .A2(G26), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT28), .Z(new_n775));
  NAND2_X1  g350(.A1(new_n485), .A2(G140), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n482), .A2(G128), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n469), .A2(G116), .ZN(new_n778));
  OAI21_X1  g353(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n776), .B(new_n777), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n775), .B1(new_n780), .B2(G29), .ZN(new_n781));
  INV_X1    g356(.A(G2067), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n766), .A2(new_n764), .ZN(new_n784));
  NOR3_X1   g359(.A1(new_n773), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n744), .A2(new_n767), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n706), .A2(G21), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G168), .B2(new_n706), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT98), .ZN(new_n789));
  INV_X1    g364(.A(G1966), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n485), .A2(G139), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT96), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT25), .ZN(new_n795));
  NAND2_X1  g370(.A1(G115), .A2(G2104), .ZN(new_n796));
  INV_X1    g371(.A(G127), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n481), .B2(new_n797), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n798), .A2(KEYINPUT97), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n469), .B1(new_n798), .B2(KEYINPUT97), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n795), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n740), .B1(new_n793), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n740), .B2(G33), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n706), .A2(G5), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G171), .B2(new_n706), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n804), .A2(G2072), .B1(G1961), .B2(new_n806), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n806), .A2(G1961), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n807), .B(new_n808), .C1(G2072), .C2(new_n804), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT99), .B(KEYINPUT23), .Z(new_n810));
  NAND2_X1  g385(.A1(new_n706), .A2(G20), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(new_n596), .B2(new_n706), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G1956), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n574), .A2(new_n706), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n706), .B2(G19), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT95), .B(G1341), .Z(new_n817));
  AOI21_X1  g392(.A(new_n814), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(new_n816), .B2(new_n817), .ZN(new_n819));
  NOR4_X1   g394(.A1(new_n786), .A2(new_n791), .A3(new_n809), .A4(new_n819), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n739), .A2(new_n820), .ZN(G311));
  NAND2_X1  g396(.A1(new_n739), .A2(new_n820), .ZN(G150));
  NAND2_X1  g397(.A1(new_n544), .A2(G93), .ZN(new_n823));
  INV_X1    g398(.A(G55), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n530), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(G80), .A2(G543), .ZN(new_n826));
  INV_X1    g401(.A(G67), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n563), .B2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT100), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n510), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI211_X1 g405(.A(KEYINPUT100), .B(new_n826), .C1(new_n563), .C2(new_n827), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n825), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(new_n568), .B2(new_n573), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n828), .A2(new_n829), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n835), .A2(new_n831), .A3(G651), .ZN(new_n836));
  INV_X1    g411(.A(new_n825), .ZN(new_n837));
  AND3_X1   g412(.A1(new_n566), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n834), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT38), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n632), .A2(G559), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT39), .ZN(new_n844));
  AOI21_X1  g419(.A(G860), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(new_n844), .B2(new_n843), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT101), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n833), .A2(G860), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(KEYINPUT37), .Z(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(G145));
  NAND2_X1  g425(.A1(new_n793), .A2(new_n801), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n754), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n485), .A2(G142), .ZN(new_n853));
  OAI21_X1  g428(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT102), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(G118), .ZN(new_n857));
  AOI22_X1  g432(.A1(new_n854), .A2(new_n855), .B1(new_n857), .B2(G2105), .ZN(new_n858));
  AOI22_X1  g433(.A1(new_n482), .A2(G130), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n853), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n652), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n852), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n780), .B(new_n508), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n716), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n862), .B(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(G160), .B(new_n648), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(G162), .ZN(new_n867));
  AOI21_X1  g442(.A(G37), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n868), .B1(new_n867), .B2(new_n865), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(KEYINPUT103), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT103), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n868), .B(new_n871), .C1(new_n867), .C2(new_n865), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n870), .A2(KEYINPUT40), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(KEYINPUT40), .B1(new_n870), .B2(new_n872), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n873), .A2(new_n874), .ZN(G395));
  XNOR2_X1  g450(.A(G303), .B(KEYINPUT104), .ZN(new_n876));
  XNOR2_X1  g451(.A(G290), .B(new_n876), .ZN(new_n877));
  XOR2_X1   g452(.A(G305), .B(G288), .Z(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n880), .A2(KEYINPUT42), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT42), .ZN(new_n882));
  OAI21_X1  g457(.A(KEYINPUT105), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n881), .B(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n840), .B(new_n640), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT41), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n632), .A2(new_n592), .A3(new_n595), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n632), .B1(new_n592), .B2(new_n595), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n886), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n632), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n596), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n892), .A2(KEYINPUT41), .A3(new_n887), .ZN(new_n893));
  AND2_X1   g468(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n885), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n888), .A2(new_n889), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n895), .B1(new_n897), .B2(new_n885), .ZN(new_n898));
  OR2_X1    g473(.A1(new_n898), .A2(KEYINPUT106), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(KEYINPUT106), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n884), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n884), .A2(new_n900), .ZN(new_n902));
  OAI21_X1  g477(.A(G868), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n903), .B1(G868), .B2(new_n832), .ZN(G295));
  OAI21_X1  g479(.A(new_n903), .B1(G868), .B2(new_n832), .ZN(G331));
  XNOR2_X1  g480(.A(G171), .B(KEYINPUT107), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(G286), .B1(new_n834), .B2(new_n839), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n569), .B1(new_n571), .B2(new_n570), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(KEYINPUT80), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n832), .B1(new_n910), .B2(new_n572), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n911), .A2(G168), .A3(new_n838), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n907), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT108), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n893), .A2(new_n914), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n892), .A2(KEYINPUT108), .A3(KEYINPUT41), .A4(new_n887), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(new_n890), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n834), .A2(new_n839), .A3(G286), .ZN(new_n918));
  OAI21_X1  g493(.A(G168), .B1(new_n911), .B2(new_n838), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n919), .A3(new_n906), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n913), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n879), .B1(new_n921), .B2(KEYINPUT109), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n896), .B1(new_n913), .B2(new_n920), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT109), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n922), .B1(new_n921), .B2(new_n925), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n918), .A2(new_n919), .A3(new_n906), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n906), .B1(new_n918), .B2(new_n919), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n897), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n890), .A2(new_n893), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n913), .A2(new_n930), .A3(new_n920), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n929), .A2(new_n880), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(G37), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT43), .B1(new_n926), .B2(new_n934), .ZN(new_n935));
  NOR3_X1   g510(.A1(new_n927), .A2(new_n928), .A3(new_n894), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n879), .B1(new_n936), .B2(new_n923), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n937), .A2(new_n933), .A3(new_n932), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n935), .B(KEYINPUT44), .C1(KEYINPUT43), .C2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n934), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n929), .A2(new_n921), .A3(KEYINPUT109), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n941), .B(new_n879), .C1(KEYINPUT109), .C2(new_n921), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT43), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n940), .A2(new_n942), .A3(KEYINPUT110), .A4(new_n943), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n926), .A2(new_n934), .A3(KEYINPUT43), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT110), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n946), .B1(new_n938), .B2(KEYINPUT43), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n944), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n948), .A2(KEYINPUT111), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT111), .B1(new_n948), .B2(new_n949), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n939), .B1(new_n950), .B2(new_n951), .ZN(G397));
  NAND2_X1  g527(.A1(new_n471), .A2(G101), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n466), .A2(G137), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n476), .A2(G40), .A3(new_n953), .A4(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT113), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT113), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n472), .A2(new_n957), .A3(G40), .A4(new_n476), .ZN(new_n958));
  AND2_X1   g533(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  XOR2_X1   g534(.A(KEYINPUT112), .B(G1384), .Z(new_n960));
  AOI21_X1  g535(.A(KEYINPUT45), .B1(new_n508), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n780), .B(new_n782), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n962), .B1(new_n963), .B2(new_n754), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT46), .B1(new_n962), .B2(G1996), .ZN(new_n965));
  OR3_X1    g540(.A1(new_n962), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n967), .B(KEYINPUT47), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n754), .B(G1996), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n963), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n718), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n716), .A2(new_n971), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n716), .A2(new_n971), .ZN(new_n973));
  OR3_X1    g548(.A1(new_n970), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n975), .A2(new_n962), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n977), .A2(KEYINPUT126), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n977), .A2(KEYINPUT126), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n962), .A2(G1986), .A3(G290), .ZN(new_n980));
  XNOR2_X1  g555(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n981));
  XOR2_X1   g556(.A(new_n980), .B(new_n981), .Z(new_n982));
  NOR3_X1   g557(.A1(new_n978), .A2(new_n979), .A3(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n962), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n972), .B(KEYINPUT125), .ZN(new_n985));
  OAI22_X1  g560(.A1(new_n985), .A2(new_n970), .B1(G2067), .B2(new_n780), .ZN(new_n986));
  AOI211_X1 g561(.A(new_n968), .B(new_n983), .C1(new_n984), .C2(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n619), .B(G1986), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n962), .B1(new_n975), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT119), .ZN(new_n990));
  INV_X1    g565(.A(G1384), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n495), .A2(KEYINPUT4), .A3(new_n497), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n500), .A2(new_n505), .A3(new_n501), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n991), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n990), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT73), .B1(new_n496), .B2(new_n492), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n506), .B1(new_n499), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(G1384), .B1(new_n998), .B2(new_n498), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n999), .A2(KEYINPUT119), .A3(KEYINPUT45), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n994), .A2(new_n995), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n996), .A2(new_n1000), .A3(new_n959), .A4(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n790), .ZN(new_n1003));
  AOI211_X1 g578(.A(KEYINPUT50), .B(G1384), .C1(new_n998), .C2(new_n498), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n956), .A2(new_n958), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1006), .B1(new_n508), .B2(new_n991), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n1004), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G2084), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1003), .A2(new_n1010), .A3(G168), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(G8), .ZN(new_n1012));
  AOI21_X1  g587(.A(G168), .B1(new_n1003), .B2(new_n1010), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT51), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1011), .A2(new_n1015), .A3(G8), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT62), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT62), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1014), .A2(new_n1019), .A3(new_n1016), .ZN(new_n1020));
  INV_X1    g595(.A(G8), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1021), .B1(new_n959), .B2(new_n999), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n1023));
  INV_X1    g598(.A(G1976), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1023), .B1(G288), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(G651), .B1(new_n538), .B2(G74), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n600), .A2(new_n599), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1026), .A2(new_n1027), .A3(KEYINPUT115), .A4(G1976), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT52), .B1(G288), .B2(new_n1024), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1022), .A2(KEYINPUT116), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n999), .A2(new_n956), .A3(new_n958), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1029), .A2(G8), .A3(new_n1032), .A4(new_n1030), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n515), .A2(G61), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n510), .B1(new_n1036), .B2(new_n603), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n515), .A2(G86), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n520), .B1(new_n1038), .B2(new_n607), .ZN(new_n1039));
  OAI21_X1  g614(.A(G1981), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n606), .A2(new_n610), .A3(new_n722), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n1040), .A2(KEYINPUT49), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT49), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1022), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1029), .A2(G8), .A3(new_n1032), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT52), .ZN(new_n1047));
  AND4_X1   g622(.A1(new_n1031), .A2(new_n1035), .A3(new_n1045), .A4(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n956), .B(new_n958), .C1(new_n999), .C2(KEYINPUT45), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n508), .A2(KEYINPUT45), .A3(new_n960), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n731), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n999), .A2(new_n1006), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n994), .A2(KEYINPUT50), .ZN(new_n1055));
  XNOR2_X1  g630(.A(KEYINPUT114), .B(G2090), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n959), .A2(new_n1054), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1021), .B1(new_n1053), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(G303), .A2(G8), .ZN(new_n1059));
  XNOR2_X1  g634(.A(new_n1059), .B(KEYINPUT55), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1049), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1001), .A2(new_n956), .A3(new_n958), .A4(new_n1051), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1008), .A2(new_n1056), .B1(new_n1063), .B2(new_n731), .ZN(new_n1064));
  OAI211_X1 g639(.A(KEYINPUT118), .B(new_n1060), .C1(new_n1064), .C2(new_n1021), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1048), .A2(new_n1062), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  OR2_X1    g642(.A1(new_n1008), .A2(G1961), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1069), .B1(new_n1063), .B2(G2078), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n761), .A2(KEYINPUT53), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1068), .B(new_n1070), .C1(new_n1002), .C2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(G171), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1067), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1018), .A2(new_n1020), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g651(.A(KEYINPUT120), .B(KEYINPUT63), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1003), .A2(new_n1010), .ZN(new_n1078));
  NOR2_X1   g653(.A1(G286), .A2(new_n1021), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1077), .B1(new_n1067), .B2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1031), .A2(new_n1035), .A3(new_n1045), .A4(new_n1047), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  AOI22_X1  g659(.A1(new_n1022), .A2(new_n1044), .B1(new_n1046), .B2(KEYINPUT52), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1085), .A2(KEYINPUT117), .A3(new_n1031), .A4(new_n1035), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1080), .A2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1087), .A2(KEYINPUT63), .A3(new_n1089), .A4(new_n1066), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1081), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1066), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1087), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1045), .A2(new_n1024), .A3(new_n724), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(new_n1041), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n1022), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1097));
  XOR2_X1   g672(.A(new_n591), .B(KEYINPUT57), .Z(new_n1098));
  NAND3_X1  g673(.A1(new_n959), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1099));
  INV_X1    g674(.A(G1956), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g676(.A(KEYINPUT56), .B(G2072), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n959), .A2(new_n1001), .A3(new_n1051), .A4(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1098), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1099), .A2(new_n764), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n959), .A2(new_n782), .A3(new_n999), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n891), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1101), .A2(new_n1098), .A3(new_n1103), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1104), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1106), .B(KEYINPUT60), .C1(new_n1008), .C2(G1348), .ZN(new_n1111));
  OR2_X1    g686(.A1(new_n1111), .A2(KEYINPUT122), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1111), .A2(KEYINPUT122), .A3(new_n891), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n891), .B1(new_n1111), .B2(KEYINPUT122), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1112), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT60), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1108), .ZN(new_n1120));
  OAI21_X1  g695(.A(KEYINPUT61), .B1(new_n1120), .B2(new_n1104), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1103), .B1(new_n1008), .B2(G1956), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1098), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT61), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1124), .A2(new_n1125), .A3(new_n1108), .ZN(new_n1126));
  XOR2_X1   g701(.A(KEYINPUT58), .B(G1341), .Z(new_n1127));
  NAND2_X1  g702(.A1(new_n1032), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT121), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT121), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1032), .A2(new_n1130), .A3(new_n1127), .ZN(new_n1131));
  INV_X1    g706(.A(G1996), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n959), .A2(new_n1001), .A3(new_n1132), .A4(new_n1051), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1129), .A2(new_n1131), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(new_n574), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(KEYINPUT59), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT59), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1134), .A2(new_n1137), .A3(new_n574), .ZN(new_n1138));
  AOI22_X1  g713(.A1(new_n1121), .A2(new_n1126), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1110), .B1(new_n1119), .B2(new_n1139), .ZN(new_n1140));
  AND4_X1   g715(.A1(new_n1066), .A2(new_n1048), .A3(new_n1062), .A4(new_n1065), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT54), .ZN(new_n1142));
  XNOR2_X1  g717(.A(G171), .B(new_n1142), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1144));
  NOR3_X1   g719(.A1(new_n961), .A2(new_n955), .A3(new_n1071), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1143), .B1(new_n1051), .B2(new_n1145), .ZN(new_n1146));
  AOI22_X1  g721(.A1(new_n1143), .A2(new_n1072), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1017), .A2(new_n1141), .A3(new_n1147), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1091), .B(new_n1097), .C1(new_n1140), .C2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1076), .B1(new_n1149), .B2(KEYINPUT123), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1111), .A2(KEYINPUT122), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(new_n632), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1111), .A2(KEYINPUT122), .A3(new_n891), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AOI22_X1  g729(.A1(new_n1154), .A2(new_n1112), .B1(new_n1117), .B2(new_n1116), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1121), .A2(new_n1126), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1109), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1159));
  AND3_X1   g734(.A1(new_n1017), .A2(new_n1141), .A3(new_n1147), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1162), .B1(new_n1081), .B2(new_n1090), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT123), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1161), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  AOI211_X1 g740(.A(KEYINPUT124), .B(new_n989), .C1(new_n1150), .C2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT124), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1149), .A2(KEYINPUT123), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1168), .A2(new_n1165), .A3(new_n1075), .ZN(new_n1169));
  INV_X1    g744(.A(new_n989), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1167), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n987), .B1(new_n1166), .B2(new_n1171), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g747(.A(new_n460), .ZN(new_n1174));
  OR4_X1    g748(.A1(new_n1174), .A2(G229), .A3(G401), .A4(G227), .ZN(new_n1175));
  AOI21_X1  g749(.A(new_n1175), .B1(new_n870), .B2(new_n872), .ZN(new_n1176));
  AND2_X1   g750(.A1(new_n1176), .A2(new_n948), .ZN(G308));
  NAND2_X1  g751(.A1(new_n1176), .A2(new_n948), .ZN(G225));
endmodule


