

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U554 ( .A1(n786), .A2(n785), .ZN(n803) );
  NOR2_X1 U555 ( .A1(n589), .A2(n588), .ZN(n591) );
  XNOR2_X1 U556 ( .A(n594), .B(KEYINPUT75), .ZN(n521) );
  NOR2_X1 U557 ( .A1(n729), .A2(n949), .ZN(n730) );
  XOR2_X1 U558 ( .A(n731), .B(KEYINPUT98), .Z(n738) );
  INV_X1 U559 ( .A(KEYINPUT99), .ZN(n758) );
  XNOR2_X1 U560 ( .A(n758), .B(KEYINPUT30), .ZN(n759) );
  XNOR2_X1 U561 ( .A(n760), .B(n759), .ZN(n761) );
  NAND2_X1 U562 ( .A1(G8), .A2(n766), .ZN(n810) );
  NOR2_X1 U563 ( .A1(G164), .A2(G1384), .ZN(n726) );
  NOR2_X1 U564 ( .A1(n632), .A2(n545), .ZN(n650) );
  XOR2_X1 U565 ( .A(KEYINPUT17), .B(n523), .Z(n897) );
  NOR2_X1 U566 ( .A1(G651), .A2(n632), .ZN(n659) );
  NAND2_X1 U567 ( .A1(n591), .A2(n590), .ZN(n949) );
  NOR2_X1 U568 ( .A1(n541), .A2(n540), .ZN(G160) );
  INV_X1 U569 ( .A(G2104), .ZN(n526) );
  AND2_X1 U570 ( .A1(n526), .A2(G2105), .ZN(n891) );
  NAND2_X1 U571 ( .A1(n891), .A2(G126), .ZN(n522) );
  XNOR2_X1 U572 ( .A(n522), .B(KEYINPUT88), .ZN(n525) );
  NOR2_X1 U573 ( .A1(G2105), .A2(G2104), .ZN(n523) );
  NAND2_X1 U574 ( .A1(G138), .A2(n897), .ZN(n524) );
  NAND2_X1 U575 ( .A1(n525), .A2(n524), .ZN(n530) );
  NOR2_X4 U576 ( .A1(G2105), .A2(n526), .ZN(n900) );
  NAND2_X1 U577 ( .A1(G102), .A2(n900), .ZN(n528) );
  AND2_X1 U578 ( .A1(G2105), .A2(G2104), .ZN(n893) );
  NAND2_X1 U579 ( .A1(G114), .A2(n893), .ZN(n527) );
  NAND2_X1 U580 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U581 ( .A1(n530), .A2(n529), .ZN(G164) );
  INV_X1 U582 ( .A(KEYINPUT66), .ZN(n536) );
  INV_X1 U583 ( .A(KEYINPUT23), .ZN(n532) );
  NAND2_X1 U584 ( .A1(n900), .A2(G101), .ZN(n531) );
  XNOR2_X1 U585 ( .A(n532), .B(n531), .ZN(n534) );
  NAND2_X1 U586 ( .A1(n891), .A2(G125), .ZN(n533) );
  NAND2_X1 U587 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U588 ( .A(n536), .B(n535), .ZN(n538) );
  NAND2_X1 U589 ( .A1(n897), .A2(G137), .ZN(n537) );
  NAND2_X1 U590 ( .A1(n538), .A2(n537), .ZN(n541) );
  NAND2_X1 U591 ( .A1(G113), .A2(n893), .ZN(n539) );
  XNOR2_X1 U592 ( .A(KEYINPUT67), .B(n539), .ZN(n540) );
  XOR2_X1 U593 ( .A(KEYINPUT0), .B(G543), .Z(n632) );
  NAND2_X1 U594 ( .A1(n659), .A2(G52), .ZN(n544) );
  XOR2_X1 U595 ( .A(KEYINPUT68), .B(G651), .Z(n545) );
  NOR2_X1 U596 ( .A1(G543), .A2(n545), .ZN(n542) );
  XOR2_X2 U597 ( .A(KEYINPUT1), .B(n542), .Z(n653) );
  NAND2_X1 U598 ( .A1(G64), .A2(n653), .ZN(n543) );
  NAND2_X1 U599 ( .A1(n544), .A2(n543), .ZN(n550) );
  NOR2_X1 U600 ( .A1(G651), .A2(G543), .ZN(n652) );
  NAND2_X1 U601 ( .A1(G90), .A2(n652), .ZN(n547) );
  NAND2_X1 U602 ( .A1(G77), .A2(n650), .ZN(n546) );
  NAND2_X1 U603 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U604 ( .A(KEYINPUT9), .B(n548), .Z(n549) );
  NOR2_X1 U605 ( .A1(n550), .A2(n549), .ZN(G171) );
  XOR2_X1 U606 ( .A(G2451), .B(G2454), .Z(n552) );
  XNOR2_X1 U607 ( .A(G2430), .B(KEYINPUT104), .ZN(n551) );
  XNOR2_X1 U608 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U609 ( .A(n553), .B(G2446), .Z(n555) );
  XNOR2_X1 U610 ( .A(G1348), .B(G1341), .ZN(n554) );
  XNOR2_X1 U611 ( .A(n555), .B(n554), .ZN(n559) );
  XOR2_X1 U612 ( .A(G2438), .B(G2427), .Z(n557) );
  XNOR2_X1 U613 ( .A(G2443), .B(G2435), .ZN(n556) );
  XNOR2_X1 U614 ( .A(n557), .B(n556), .ZN(n558) );
  XOR2_X1 U615 ( .A(n559), .B(n558), .Z(n560) );
  AND2_X1 U616 ( .A1(G14), .A2(n560), .ZN(G401) );
  AND2_X1 U617 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U618 ( .A1(G99), .A2(n900), .ZN(n562) );
  NAND2_X1 U619 ( .A1(G111), .A2(n893), .ZN(n561) );
  NAND2_X1 U620 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U621 ( .A(KEYINPUT78), .B(n563), .ZN(n566) );
  NAND2_X1 U622 ( .A1(n891), .A2(G123), .ZN(n564) );
  XOR2_X1 U623 ( .A(KEYINPUT18), .B(n564), .Z(n565) );
  NOR2_X1 U624 ( .A1(n566), .A2(n565), .ZN(n568) );
  NAND2_X1 U625 ( .A1(n897), .A2(G135), .ZN(n567) );
  NAND2_X1 U626 ( .A1(n568), .A2(n567), .ZN(n1010) );
  XNOR2_X1 U627 ( .A(G2096), .B(n1010), .ZN(n569) );
  OR2_X1 U628 ( .A1(G2100), .A2(n569), .ZN(G156) );
  INV_X1 U629 ( .A(G57), .ZN(G237) );
  NAND2_X1 U630 ( .A1(n652), .A2(G89), .ZN(n570) );
  XNOR2_X1 U631 ( .A(n570), .B(KEYINPUT4), .ZN(n572) );
  NAND2_X1 U632 ( .A1(G76), .A2(n650), .ZN(n571) );
  NAND2_X1 U633 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U634 ( .A(n573), .B(KEYINPUT5), .ZN(n578) );
  NAND2_X1 U635 ( .A1(n659), .A2(G51), .ZN(n575) );
  NAND2_X1 U636 ( .A1(G63), .A2(n653), .ZN(n574) );
  NAND2_X1 U637 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U638 ( .A(KEYINPUT6), .B(n576), .Z(n577) );
  NAND2_X1 U639 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U640 ( .A(n579), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U641 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U642 ( .A(KEYINPUT73), .B(KEYINPUT10), .Z(n581) );
  NAND2_X1 U643 ( .A1(G7), .A2(G661), .ZN(n580) );
  XNOR2_X1 U644 ( .A(n581), .B(n580), .ZN(G223) );
  INV_X1 U645 ( .A(G223), .ZN(n836) );
  NAND2_X1 U646 ( .A1(n836), .A2(G567), .ZN(n582) );
  XOR2_X1 U647 ( .A(KEYINPUT11), .B(n582), .Z(G234) );
  NAND2_X1 U648 ( .A1(n653), .A2(G56), .ZN(n583) );
  XOR2_X1 U649 ( .A(KEYINPUT14), .B(n583), .Z(n589) );
  NAND2_X1 U650 ( .A1(n652), .A2(G81), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n584), .B(KEYINPUT12), .ZN(n586) );
  NAND2_X1 U652 ( .A1(G68), .A2(n650), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U654 ( .A(KEYINPUT13), .B(n587), .Z(n588) );
  NAND2_X1 U655 ( .A1(n659), .A2(G43), .ZN(n590) );
  INV_X1 U656 ( .A(G860), .ZN(n612) );
  OR2_X1 U657 ( .A1(n949), .A2(n612), .ZN(G153) );
  NAND2_X1 U658 ( .A1(G171), .A2(G868), .ZN(n601) );
  NAND2_X1 U659 ( .A1(n659), .A2(G54), .ZN(n593) );
  NAND2_X1 U660 ( .A1(G79), .A2(n650), .ZN(n592) );
  NAND2_X1 U661 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U662 ( .A1(G66), .A2(n653), .ZN(n595) );
  NAND2_X1 U663 ( .A1(n521), .A2(n595), .ZN(n598) );
  NAND2_X1 U664 ( .A1(n652), .A2(G92), .ZN(n596) );
  XOR2_X1 U665 ( .A(KEYINPUT74), .B(n596), .Z(n597) );
  NOR2_X1 U666 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X2 U667 ( .A(KEYINPUT15), .B(n599), .Z(n948) );
  INV_X1 U668 ( .A(G868), .ZN(n672) );
  NAND2_X1 U669 ( .A1(n948), .A2(n672), .ZN(n600) );
  NAND2_X1 U670 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U671 ( .A(KEYINPUT76), .B(n602), .Z(G284) );
  NAND2_X1 U672 ( .A1(G65), .A2(n653), .ZN(n605) );
  NAND2_X1 U673 ( .A1(G91), .A2(n652), .ZN(n603) );
  XOR2_X1 U674 ( .A(KEYINPUT71), .B(n603), .Z(n604) );
  NAND2_X1 U675 ( .A1(n605), .A2(n604), .ZN(n609) );
  NAND2_X1 U676 ( .A1(n659), .A2(G53), .ZN(n607) );
  NAND2_X1 U677 ( .A1(G78), .A2(n650), .ZN(n606) );
  NAND2_X1 U678 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U679 ( .A1(n609), .A2(n608), .ZN(n958) );
  XOR2_X1 U680 ( .A(n958), .B(KEYINPUT72), .Z(G299) );
  NOR2_X1 U681 ( .A1(G299), .A2(G868), .ZN(n611) );
  NOR2_X1 U682 ( .A1(G286), .A2(n672), .ZN(n610) );
  NOR2_X1 U683 ( .A1(n611), .A2(n610), .ZN(G297) );
  NAND2_X1 U684 ( .A1(n612), .A2(G559), .ZN(n613) );
  NAND2_X1 U685 ( .A1(n613), .A2(n948), .ZN(n614) );
  XNOR2_X1 U686 ( .A(n614), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U687 ( .A1(G559), .A2(n672), .ZN(n615) );
  NAND2_X1 U688 ( .A1(n948), .A2(n615), .ZN(n616) );
  XNOR2_X1 U689 ( .A(n616), .B(KEYINPUT77), .ZN(n618) );
  NOR2_X1 U690 ( .A1(n949), .A2(G868), .ZN(n617) );
  NOR2_X1 U691 ( .A1(n618), .A2(n617), .ZN(G282) );
  NAND2_X1 U692 ( .A1(G559), .A2(n948), .ZN(n619) );
  XNOR2_X1 U693 ( .A(n619), .B(n949), .ZN(n668) );
  NOR2_X1 U694 ( .A1(n668), .A2(G860), .ZN(n627) );
  NAND2_X1 U695 ( .A1(n659), .A2(G55), .ZN(n621) );
  NAND2_X1 U696 ( .A1(G67), .A2(n653), .ZN(n620) );
  NAND2_X1 U697 ( .A1(n621), .A2(n620), .ZN(n626) );
  NAND2_X1 U698 ( .A1(G93), .A2(n652), .ZN(n623) );
  NAND2_X1 U699 ( .A1(G80), .A2(n650), .ZN(n622) );
  NAND2_X1 U700 ( .A1(n623), .A2(n622), .ZN(n624) );
  XOR2_X1 U701 ( .A(KEYINPUT79), .B(n624), .Z(n625) );
  OR2_X1 U702 ( .A1(n626), .A2(n625), .ZN(n671) );
  XOR2_X1 U703 ( .A(n627), .B(n671), .Z(G145) );
  NAND2_X1 U704 ( .A1(G49), .A2(n659), .ZN(n629) );
  NAND2_X1 U705 ( .A1(G74), .A2(G651), .ZN(n628) );
  NAND2_X1 U706 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U707 ( .A(KEYINPUT80), .B(n630), .ZN(n631) );
  NOR2_X1 U708 ( .A1(n653), .A2(n631), .ZN(n634) );
  NAND2_X1 U709 ( .A1(n632), .A2(G87), .ZN(n633) );
  NAND2_X1 U710 ( .A1(n634), .A2(n633), .ZN(G288) );
  NAND2_X1 U711 ( .A1(G47), .A2(n659), .ZN(n635) );
  XNOR2_X1 U712 ( .A(n635), .B(KEYINPUT70), .ZN(n642) );
  NAND2_X1 U713 ( .A1(G85), .A2(n652), .ZN(n637) );
  NAND2_X1 U714 ( .A1(G72), .A2(n650), .ZN(n636) );
  NAND2_X1 U715 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U716 ( .A1(G60), .A2(n653), .ZN(n638) );
  XNOR2_X1 U717 ( .A(KEYINPUT69), .B(n638), .ZN(n639) );
  NOR2_X1 U718 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U719 ( .A1(n642), .A2(n641), .ZN(G290) );
  NAND2_X1 U720 ( .A1(G88), .A2(n652), .ZN(n644) );
  NAND2_X1 U721 ( .A1(G50), .A2(n659), .ZN(n643) );
  NAND2_X1 U722 ( .A1(n644), .A2(n643), .ZN(n647) );
  NAND2_X1 U723 ( .A1(n650), .A2(G75), .ZN(n645) );
  XOR2_X1 U724 ( .A(KEYINPUT82), .B(n645), .Z(n646) );
  NOR2_X1 U725 ( .A1(n647), .A2(n646), .ZN(n649) );
  NAND2_X1 U726 ( .A1(G62), .A2(n653), .ZN(n648) );
  NAND2_X1 U727 ( .A1(n649), .A2(n648), .ZN(G303) );
  INV_X1 U728 ( .A(G303), .ZN(G166) );
  NAND2_X1 U729 ( .A1(n650), .A2(G73), .ZN(n651) );
  XOR2_X1 U730 ( .A(KEYINPUT2), .B(n651), .Z(n658) );
  NAND2_X1 U731 ( .A1(n652), .A2(G86), .ZN(n655) );
  NAND2_X1 U732 ( .A1(G61), .A2(n653), .ZN(n654) );
  NAND2_X1 U733 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U734 ( .A(KEYINPUT81), .B(n656), .Z(n657) );
  NOR2_X1 U735 ( .A1(n658), .A2(n657), .ZN(n661) );
  NAND2_X1 U736 ( .A1(n659), .A2(G48), .ZN(n660) );
  NAND2_X1 U737 ( .A1(n661), .A2(n660), .ZN(G305) );
  XNOR2_X1 U738 ( .A(KEYINPUT83), .B(KEYINPUT19), .ZN(n663) );
  XNOR2_X1 U739 ( .A(G288), .B(G299), .ZN(n662) );
  XNOR2_X1 U740 ( .A(n663), .B(n662), .ZN(n664) );
  XOR2_X1 U741 ( .A(n671), .B(n664), .Z(n666) );
  XNOR2_X1 U742 ( .A(G290), .B(G166), .ZN(n665) );
  XNOR2_X1 U743 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U744 ( .A(n667), .B(G305), .ZN(n865) );
  XNOR2_X1 U745 ( .A(n865), .B(n668), .ZN(n669) );
  NAND2_X1 U746 ( .A1(n669), .A2(G868), .ZN(n670) );
  XNOR2_X1 U747 ( .A(n670), .B(KEYINPUT84), .ZN(n674) );
  NAND2_X1 U748 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U749 ( .A1(n674), .A2(n673), .ZN(G295) );
  NAND2_X1 U750 ( .A1(G2078), .A2(G2084), .ZN(n675) );
  XOR2_X1 U751 ( .A(KEYINPUT20), .B(n675), .Z(n676) );
  NAND2_X1 U752 ( .A1(G2090), .A2(n676), .ZN(n677) );
  XNOR2_X1 U753 ( .A(KEYINPUT21), .B(n677), .ZN(n678) );
  NAND2_X1 U754 ( .A1(n678), .A2(G2072), .ZN(G158) );
  XOR2_X1 U755 ( .A(KEYINPUT85), .B(G44), .Z(n679) );
  XNOR2_X1 U756 ( .A(KEYINPUT3), .B(n679), .ZN(G218) );
  NAND2_X1 U757 ( .A1(G132), .A2(G82), .ZN(n680) );
  XNOR2_X1 U758 ( .A(n680), .B(KEYINPUT22), .ZN(n681) );
  XNOR2_X1 U759 ( .A(n681), .B(KEYINPUT86), .ZN(n682) );
  NOR2_X1 U760 ( .A1(G218), .A2(n682), .ZN(n683) );
  NAND2_X1 U761 ( .A1(G96), .A2(n683), .ZN(n843) );
  NAND2_X1 U762 ( .A1(G2106), .A2(n843), .ZN(n687) );
  NAND2_X1 U763 ( .A1(G69), .A2(G120), .ZN(n684) );
  NOR2_X1 U764 ( .A1(G237), .A2(n684), .ZN(n685) );
  NAND2_X1 U765 ( .A1(G108), .A2(n685), .ZN(n842) );
  NAND2_X1 U766 ( .A1(G567), .A2(n842), .ZN(n686) );
  NAND2_X1 U767 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U768 ( .A(KEYINPUT87), .B(n688), .ZN(G319) );
  INV_X1 U769 ( .A(G319), .ZN(n915) );
  NAND2_X1 U770 ( .A1(G661), .A2(G483), .ZN(n689) );
  NOR2_X1 U771 ( .A1(n915), .A2(n689), .ZN(n839) );
  NAND2_X1 U772 ( .A1(n839), .A2(G36), .ZN(G176) );
  NAND2_X1 U773 ( .A1(G129), .A2(n891), .ZN(n691) );
  NAND2_X1 U774 ( .A1(G117), .A2(n893), .ZN(n690) );
  NAND2_X1 U775 ( .A1(n691), .A2(n690), .ZN(n695) );
  NAND2_X1 U776 ( .A1(G105), .A2(n900), .ZN(n692) );
  XNOR2_X1 U777 ( .A(n692), .B(KEYINPUT38), .ZN(n693) );
  XNOR2_X1 U778 ( .A(n693), .B(KEYINPUT93), .ZN(n694) );
  NOR2_X1 U779 ( .A1(n695), .A2(n694), .ZN(n697) );
  NAND2_X1 U780 ( .A1(n897), .A2(G141), .ZN(n696) );
  NAND2_X1 U781 ( .A1(n697), .A2(n696), .ZN(n888) );
  NAND2_X1 U782 ( .A1(n888), .A2(G1996), .ZN(n706) );
  NAND2_X1 U783 ( .A1(G95), .A2(n900), .ZN(n699) );
  NAND2_X1 U784 ( .A1(G107), .A2(n893), .ZN(n698) );
  NAND2_X1 U785 ( .A1(n699), .A2(n698), .ZN(n703) );
  NAND2_X1 U786 ( .A1(G119), .A2(n891), .ZN(n701) );
  NAND2_X1 U787 ( .A1(G131), .A2(n897), .ZN(n700) );
  NAND2_X1 U788 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U789 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U790 ( .A(KEYINPUT92), .B(n704), .Z(n905) );
  NAND2_X1 U791 ( .A1(n905), .A2(G1991), .ZN(n705) );
  NAND2_X1 U792 ( .A1(n706), .A2(n705), .ZN(n1005) );
  NAND2_X1 U793 ( .A1(G160), .A2(G40), .ZN(n724) );
  NOR2_X1 U794 ( .A1(n726), .A2(n724), .ZN(n830) );
  AND2_X1 U795 ( .A1(n1005), .A2(n830), .ZN(n823) );
  XOR2_X1 U796 ( .A(KEYINPUT94), .B(n823), .Z(n718) );
  XNOR2_X1 U797 ( .A(KEYINPUT37), .B(G2067), .ZN(n828) );
  XNOR2_X1 U798 ( .A(KEYINPUT91), .B(KEYINPUT36), .ZN(n717) );
  NAND2_X1 U799 ( .A1(G128), .A2(n891), .ZN(n708) );
  NAND2_X1 U800 ( .A1(G116), .A2(n893), .ZN(n707) );
  NAND2_X1 U801 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U802 ( .A(KEYINPUT35), .B(n709), .ZN(n715) );
  NAND2_X1 U803 ( .A1(G104), .A2(n900), .ZN(n711) );
  NAND2_X1 U804 ( .A1(G140), .A2(n897), .ZN(n710) );
  NAND2_X1 U805 ( .A1(n711), .A2(n710), .ZN(n713) );
  XOR2_X1 U806 ( .A(KEYINPUT34), .B(KEYINPUT90), .Z(n712) );
  XNOR2_X1 U807 ( .A(n713), .B(n712), .ZN(n714) );
  NAND2_X1 U808 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U809 ( .A(n717), .B(n716), .ZN(n912) );
  NOR2_X1 U810 ( .A1(n828), .A2(n912), .ZN(n1020) );
  NAND2_X1 U811 ( .A1(n830), .A2(n1020), .ZN(n826) );
  NAND2_X1 U812 ( .A1(n718), .A2(n826), .ZN(n817) );
  NOR2_X1 U813 ( .A1(G1971), .A2(G303), .ZN(n787) );
  XNOR2_X1 U814 ( .A(G1996), .B(KEYINPUT97), .ZN(n932) );
  INV_X1 U815 ( .A(n932), .ZN(n719) );
  AND2_X1 U816 ( .A1(n719), .A2(G40), .ZN(n720) );
  AND2_X1 U817 ( .A1(G160), .A2(n720), .ZN(n721) );
  AND2_X1 U818 ( .A1(n726), .A2(n721), .ZN(n723) );
  XOR2_X1 U819 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n722) );
  XNOR2_X1 U820 ( .A(n723), .B(n722), .ZN(n728) );
  INV_X1 U821 ( .A(n724), .ZN(n725) );
  NAND2_X1 U822 ( .A1(n726), .A2(n725), .ZN(n766) );
  NAND2_X1 U823 ( .A1(n766), .A2(G1341), .ZN(n727) );
  NAND2_X1 U824 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U825 ( .A(KEYINPUT65), .B(n730), .Z(n732) );
  NOR2_X1 U826 ( .A1(n732), .A2(n948), .ZN(n731) );
  NAND2_X1 U827 ( .A1(n732), .A2(n948), .ZN(n736) );
  INV_X1 U828 ( .A(n766), .ZN(n750) );
  NOR2_X1 U829 ( .A1(n750), .A2(G1348), .ZN(n734) );
  NOR2_X1 U830 ( .A1(G2067), .A2(n766), .ZN(n733) );
  NOR2_X1 U831 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U832 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U833 ( .A1(n738), .A2(n737), .ZN(n743) );
  NAND2_X1 U834 ( .A1(n750), .A2(G2072), .ZN(n739) );
  XNOR2_X1 U835 ( .A(n739), .B(KEYINPUT27), .ZN(n741) );
  INV_X1 U836 ( .A(G1956), .ZN(n970) );
  NOR2_X1 U837 ( .A1(n970), .A2(n750), .ZN(n740) );
  NOR2_X1 U838 ( .A1(n741), .A2(n740), .ZN(n744) );
  NAND2_X1 U839 ( .A1(n958), .A2(n744), .ZN(n742) );
  NAND2_X1 U840 ( .A1(n743), .A2(n742), .ZN(n747) );
  NOR2_X1 U841 ( .A1(n958), .A2(n744), .ZN(n745) );
  XOR2_X1 U842 ( .A(n745), .B(KEYINPUT28), .Z(n746) );
  NAND2_X1 U843 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U844 ( .A(KEYINPUT29), .B(n748), .ZN(n749) );
  INV_X1 U845 ( .A(n749), .ZN(n755) );
  OR2_X1 U846 ( .A1(n750), .A2(G1961), .ZN(n752) );
  XNOR2_X1 U847 ( .A(G2078), .B(KEYINPUT25), .ZN(n931) );
  NAND2_X1 U848 ( .A1(n750), .A2(n931), .ZN(n751) );
  NAND2_X1 U849 ( .A1(n752), .A2(n751), .ZN(n756) );
  AND2_X1 U850 ( .A1(n756), .A2(G171), .ZN(n753) );
  XOR2_X1 U851 ( .A(KEYINPUT96), .B(n753), .Z(n754) );
  NAND2_X1 U852 ( .A1(n755), .A2(n754), .ZN(n778) );
  NOR2_X1 U853 ( .A1(G171), .A2(n756), .ZN(n763) );
  NOR2_X1 U854 ( .A1(G1966), .A2(n810), .ZN(n784) );
  NOR2_X1 U855 ( .A1(G2084), .A2(n766), .ZN(n780) );
  NOR2_X1 U856 ( .A1(n784), .A2(n780), .ZN(n757) );
  NAND2_X1 U857 ( .A1(G8), .A2(n757), .ZN(n760) );
  NOR2_X1 U858 ( .A1(G168), .A2(n761), .ZN(n762) );
  NOR2_X1 U859 ( .A1(n763), .A2(n762), .ZN(n764) );
  XOR2_X1 U860 ( .A(KEYINPUT31), .B(n764), .Z(n779) );
  INV_X1 U861 ( .A(G8), .ZN(n771) );
  NOR2_X1 U862 ( .A1(G1971), .A2(n810), .ZN(n765) );
  XNOR2_X1 U863 ( .A(n765), .B(KEYINPUT100), .ZN(n768) );
  NOR2_X1 U864 ( .A1(n766), .A2(G2090), .ZN(n767) );
  NOR2_X1 U865 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U866 ( .A1(n769), .A2(G303), .ZN(n770) );
  OR2_X1 U867 ( .A1(n771), .A2(n770), .ZN(n773) );
  AND2_X1 U868 ( .A1(n779), .A2(n773), .ZN(n772) );
  NAND2_X1 U869 ( .A1(n778), .A2(n772), .ZN(n776) );
  INV_X1 U870 ( .A(n773), .ZN(n774) );
  OR2_X1 U871 ( .A1(n774), .A2(G286), .ZN(n775) );
  NAND2_X1 U872 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U873 ( .A(KEYINPUT32), .B(n777), .Z(n786) );
  NAND2_X1 U874 ( .A1(n779), .A2(n778), .ZN(n782) );
  NAND2_X1 U875 ( .A1(G8), .A2(n780), .ZN(n781) );
  NAND2_X1 U876 ( .A1(n782), .A2(n781), .ZN(n783) );
  NOR2_X1 U877 ( .A1(n784), .A2(n783), .ZN(n785) );
  NOR2_X1 U878 ( .A1(n787), .A2(n803), .ZN(n789) );
  NOR2_X1 U879 ( .A1(G288), .A2(G1976), .ZN(n788) );
  XNOR2_X1 U880 ( .A(n788), .B(KEYINPUT101), .ZN(n961) );
  NAND2_X1 U881 ( .A1(n789), .A2(n961), .ZN(n792) );
  INV_X1 U882 ( .A(KEYINPUT102), .ZN(n794) );
  NOR2_X1 U883 ( .A1(n810), .A2(n794), .ZN(n790) );
  NAND2_X1 U884 ( .A1(G1976), .A2(G288), .ZN(n956) );
  AND2_X1 U885 ( .A1(n790), .A2(n956), .ZN(n791) );
  AND2_X1 U886 ( .A1(n792), .A2(n791), .ZN(n793) );
  NOR2_X1 U887 ( .A1(n793), .A2(KEYINPUT33), .ZN(n801) );
  INV_X1 U888 ( .A(n961), .ZN(n795) );
  NAND2_X1 U889 ( .A1(n794), .A2(n795), .ZN(n798) );
  NAND2_X1 U890 ( .A1(n795), .A2(KEYINPUT33), .ZN(n796) );
  NAND2_X1 U891 ( .A1(n796), .A2(KEYINPUT102), .ZN(n797) );
  NAND2_X1 U892 ( .A1(n798), .A2(n797), .ZN(n799) );
  NOR2_X1 U893 ( .A1(n810), .A2(n799), .ZN(n800) );
  NOR2_X1 U894 ( .A1(n801), .A2(n800), .ZN(n802) );
  XOR2_X1 U895 ( .A(G1981), .B(G305), .Z(n945) );
  NAND2_X1 U896 ( .A1(n802), .A2(n945), .ZN(n815) );
  INV_X1 U897 ( .A(n803), .ZN(n806) );
  NOR2_X1 U898 ( .A1(G2090), .A2(G303), .ZN(n804) );
  NAND2_X1 U899 ( .A1(G8), .A2(n804), .ZN(n805) );
  NAND2_X1 U900 ( .A1(n806), .A2(n805), .ZN(n807) );
  NAND2_X1 U901 ( .A1(n807), .A2(n810), .ZN(n813) );
  NOR2_X1 U902 ( .A1(G1981), .A2(G305), .ZN(n808) );
  XNOR2_X1 U903 ( .A(n808), .B(KEYINPUT24), .ZN(n809) );
  XNOR2_X1 U904 ( .A(n809), .B(KEYINPUT95), .ZN(n811) );
  OR2_X1 U905 ( .A1(n811), .A2(n810), .ZN(n812) );
  AND2_X1 U906 ( .A1(n813), .A2(n812), .ZN(n814) );
  AND2_X1 U907 ( .A1(n815), .A2(n814), .ZN(n816) );
  NOR2_X1 U908 ( .A1(n817), .A2(n816), .ZN(n820) );
  XOR2_X1 U909 ( .A(G1986), .B(KEYINPUT89), .Z(n818) );
  XNOR2_X1 U910 ( .A(G290), .B(n818), .ZN(n953) );
  NAND2_X1 U911 ( .A1(n953), .A2(n830), .ZN(n819) );
  NAND2_X1 U912 ( .A1(n820), .A2(n819), .ZN(n833) );
  NOR2_X1 U913 ( .A1(G1996), .A2(n888), .ZN(n1013) );
  NOR2_X1 U914 ( .A1(G1991), .A2(n905), .ZN(n1009) );
  NOR2_X1 U915 ( .A1(G1986), .A2(G290), .ZN(n821) );
  NOR2_X1 U916 ( .A1(n1009), .A2(n821), .ZN(n822) );
  NOR2_X1 U917 ( .A1(n823), .A2(n822), .ZN(n824) );
  NOR2_X1 U918 ( .A1(n1013), .A2(n824), .ZN(n825) );
  XNOR2_X1 U919 ( .A(n825), .B(KEYINPUT39), .ZN(n827) );
  NAND2_X1 U920 ( .A1(n827), .A2(n826), .ZN(n829) );
  NAND2_X1 U921 ( .A1(n828), .A2(n912), .ZN(n1017) );
  NAND2_X1 U922 ( .A1(n829), .A2(n1017), .ZN(n831) );
  NAND2_X1 U923 ( .A1(n831), .A2(n830), .ZN(n832) );
  NAND2_X1 U924 ( .A1(n833), .A2(n832), .ZN(n835) );
  XOR2_X1 U925 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n834) );
  XNOR2_X1 U926 ( .A(n835), .B(n834), .ZN(G329) );
  NAND2_X1 U927 ( .A1(G2106), .A2(n836), .ZN(G217) );
  NAND2_X1 U928 ( .A1(G15), .A2(G2), .ZN(n837) );
  XNOR2_X1 U929 ( .A(KEYINPUT105), .B(n837), .ZN(n838) );
  NAND2_X1 U930 ( .A1(n838), .A2(G661), .ZN(G259) );
  NAND2_X1 U931 ( .A1(G1), .A2(G3), .ZN(n840) );
  NAND2_X1 U932 ( .A1(n840), .A2(n839), .ZN(n841) );
  XNOR2_X1 U933 ( .A(n841), .B(KEYINPUT106), .ZN(G188) );
  INV_X1 U935 ( .A(G132), .ZN(G219) );
  INV_X1 U936 ( .A(G120), .ZN(G236) );
  INV_X1 U937 ( .A(G82), .ZN(G220) );
  INV_X1 U938 ( .A(G69), .ZN(G235) );
  NOR2_X1 U939 ( .A1(n843), .A2(n842), .ZN(n844) );
  XNOR2_X1 U940 ( .A(n844), .B(KEYINPUT107), .ZN(G261) );
  INV_X1 U941 ( .A(G261), .ZN(G325) );
  XOR2_X1 U942 ( .A(G2100), .B(G2096), .Z(n846) );
  XNOR2_X1 U943 ( .A(KEYINPUT42), .B(G2678), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U945 ( .A(KEYINPUT43), .B(G2090), .Z(n848) );
  XNOR2_X1 U946 ( .A(G2067), .B(G2072), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U948 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U949 ( .A(G2078), .B(G2084), .ZN(n851) );
  XNOR2_X1 U950 ( .A(n852), .B(n851), .ZN(G227) );
  XOR2_X1 U951 ( .A(G1981), .B(G1966), .Z(n854) );
  XNOR2_X1 U952 ( .A(G1996), .B(G1991), .ZN(n853) );
  XNOR2_X1 U953 ( .A(n854), .B(n853), .ZN(n864) );
  XOR2_X1 U954 ( .A(KEYINPUT109), .B(KEYINPUT41), .Z(n856) );
  XNOR2_X1 U955 ( .A(G1986), .B(KEYINPUT110), .ZN(n855) );
  XNOR2_X1 U956 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U957 ( .A(G1976), .B(G1971), .Z(n858) );
  XNOR2_X1 U958 ( .A(G1956), .B(G1961), .ZN(n857) );
  XNOR2_X1 U959 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U960 ( .A(n860), .B(n859), .Z(n862) );
  XNOR2_X1 U961 ( .A(KEYINPUT108), .B(G2474), .ZN(n861) );
  XNOR2_X1 U962 ( .A(n862), .B(n861), .ZN(n863) );
  XNOR2_X1 U963 ( .A(n864), .B(n863), .ZN(G229) );
  XNOR2_X1 U964 ( .A(G286), .B(n865), .ZN(n867) );
  XNOR2_X1 U965 ( .A(n949), .B(G171), .ZN(n866) );
  XNOR2_X1 U966 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U967 ( .A(n948), .B(n868), .Z(n869) );
  NOR2_X1 U968 ( .A1(G37), .A2(n869), .ZN(n870) );
  XNOR2_X1 U969 ( .A(KEYINPUT116), .B(n870), .ZN(G397) );
  NAND2_X1 U970 ( .A1(G100), .A2(n900), .ZN(n872) );
  NAND2_X1 U971 ( .A1(G112), .A2(n893), .ZN(n871) );
  NAND2_X1 U972 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U973 ( .A(n873), .B(KEYINPUT111), .ZN(n875) );
  NAND2_X1 U974 ( .A1(G136), .A2(n897), .ZN(n874) );
  NAND2_X1 U975 ( .A1(n875), .A2(n874), .ZN(n878) );
  NAND2_X1 U976 ( .A1(n891), .A2(G124), .ZN(n876) );
  XOR2_X1 U977 ( .A(KEYINPUT44), .B(n876), .Z(n877) );
  NOR2_X1 U978 ( .A1(n878), .A2(n877), .ZN(G162) );
  NAND2_X1 U979 ( .A1(G130), .A2(n891), .ZN(n880) );
  NAND2_X1 U980 ( .A1(G118), .A2(n893), .ZN(n879) );
  NAND2_X1 U981 ( .A1(n880), .A2(n879), .ZN(n885) );
  NAND2_X1 U982 ( .A1(G106), .A2(n900), .ZN(n882) );
  NAND2_X1 U983 ( .A1(G142), .A2(n897), .ZN(n881) );
  NAND2_X1 U984 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U985 ( .A(n883), .B(KEYINPUT45), .Z(n884) );
  NOR2_X1 U986 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U987 ( .A(KEYINPUT48), .B(n886), .Z(n887) );
  XNOR2_X1 U988 ( .A(KEYINPUT46), .B(n887), .ZN(n890) );
  XNOR2_X1 U989 ( .A(n888), .B(KEYINPUT114), .ZN(n889) );
  XNOR2_X1 U990 ( .A(n890), .B(n889), .ZN(n904) );
  NAND2_X1 U991 ( .A1(n891), .A2(G127), .ZN(n892) );
  XOR2_X1 U992 ( .A(KEYINPUT113), .B(n892), .Z(n895) );
  NAND2_X1 U993 ( .A1(n893), .A2(G115), .ZN(n894) );
  NAND2_X1 U994 ( .A1(n895), .A2(n894), .ZN(n896) );
  XNOR2_X1 U995 ( .A(n896), .B(KEYINPUT47), .ZN(n899) );
  NAND2_X1 U996 ( .A1(G139), .A2(n897), .ZN(n898) );
  NAND2_X1 U997 ( .A1(n899), .A2(n898), .ZN(n903) );
  NAND2_X1 U998 ( .A1(n900), .A2(G103), .ZN(n901) );
  XOR2_X1 U999 ( .A(KEYINPUT112), .B(n901), .Z(n902) );
  NOR2_X1 U1000 ( .A1(n903), .A2(n902), .ZN(n1001) );
  XOR2_X1 U1001 ( .A(n904), .B(n1001), .Z(n907) );
  XNOR2_X1 U1002 ( .A(n905), .B(G162), .ZN(n906) );
  XNOR2_X1 U1003 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1004 ( .A(n1010), .B(n908), .ZN(n910) );
  XNOR2_X1 U1005 ( .A(G164), .B(G160), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1007 ( .A(n912), .B(n911), .Z(n913) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n913), .ZN(n914) );
  XOR2_X1 U1009 ( .A(KEYINPUT115), .B(n914), .Z(G395) );
  NOR2_X1 U1010 ( .A1(G401), .A2(n915), .ZN(n916) );
  XOR2_X1 U1011 ( .A(KEYINPUT117), .B(n916), .Z(n920) );
  NOR2_X1 U1012 ( .A1(G227), .A2(G229), .ZN(n917) );
  XOR2_X1 U1013 ( .A(KEYINPUT49), .B(n917), .Z(n918) );
  XNOR2_X1 U1014 ( .A(KEYINPUT118), .B(n918), .ZN(n919) );
  NAND2_X1 U1015 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1016 ( .A(KEYINPUT119), .B(n921), .ZN(n923) );
  NOR2_X1 U1017 ( .A1(G397), .A2(G395), .ZN(n922) );
  NAND2_X1 U1018 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1019 ( .A(KEYINPUT120), .B(n924), .ZN(G225) );
  XNOR2_X1 U1020 ( .A(KEYINPUT121), .B(G225), .ZN(G308) );
  INV_X1 U1021 ( .A(G108), .ZN(G238) );
  INV_X1 U1022 ( .A(G96), .ZN(G221) );
  XOR2_X1 U1023 ( .A(G2090), .B(G35), .Z(n927) );
  XOR2_X1 U1024 ( .A(KEYINPUT54), .B(G34), .Z(n925) );
  XNOR2_X1 U1025 ( .A(n925), .B(G2084), .ZN(n926) );
  NAND2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n942) );
  XOR2_X1 U1027 ( .A(G1991), .B(G25), .Z(n928) );
  NAND2_X1 U1028 ( .A1(n928), .A2(G28), .ZN(n938) );
  XNOR2_X1 U1029 ( .A(G2067), .B(G26), .ZN(n930) );
  XNOR2_X1 U1030 ( .A(G33), .B(G2072), .ZN(n929) );
  NOR2_X1 U1031 ( .A1(n930), .A2(n929), .ZN(n936) );
  XOR2_X1 U1032 ( .A(n931), .B(G27), .Z(n934) );
  XOR2_X1 U1033 ( .A(n932), .B(G32), .Z(n933) );
  NOR2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1036 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1037 ( .A(KEYINPUT123), .B(n939), .Z(n940) );
  XNOR2_X1 U1038 ( .A(n940), .B(KEYINPUT53), .ZN(n941) );
  NOR2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1040 ( .A(KEYINPUT55), .B(n943), .Z(n944) );
  NOR2_X1 U1041 ( .A1(G29), .A2(n944), .ZN(n998) );
  XNOR2_X1 U1042 ( .A(G16), .B(KEYINPUT56), .ZN(n969) );
  XNOR2_X1 U1043 ( .A(G1966), .B(G168), .ZN(n946) );
  NAND2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1045 ( .A(n947), .B(KEYINPUT57), .ZN(n967) );
  XNOR2_X1 U1046 ( .A(G1348), .B(n948), .ZN(n955) );
  XOR2_X1 U1047 ( .A(n949), .B(G1341), .Z(n951) );
  XNOR2_X1 U1048 ( .A(G171), .B(G1961), .ZN(n950) );
  NAND2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1050 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n965) );
  XNOR2_X1 U1052 ( .A(G166), .B(G1971), .ZN(n957) );
  NAND2_X1 U1053 ( .A1(n957), .A2(n956), .ZN(n960) );
  XOR2_X1 U1054 ( .A(n958), .B(G1956), .Z(n959) );
  NOR2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n962) );
  NAND2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(KEYINPUT124), .B(n963), .ZN(n964) );
  NOR2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1059 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1060 ( .A1(n969), .A2(n968), .ZN(n996) );
  INV_X1 U1061 ( .A(G16), .ZN(n994) );
  XOR2_X1 U1062 ( .A(G1961), .B(G5), .Z(n990) );
  XOR2_X1 U1063 ( .A(G1966), .B(G21), .Z(n980) );
  XNOR2_X1 U1064 ( .A(G20), .B(n970), .ZN(n974) );
  XNOR2_X1 U1065 ( .A(G1341), .B(G19), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(G1981), .B(G6), .ZN(n971) );
  NOR2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n977) );
  XOR2_X1 U1069 ( .A(KEYINPUT59), .B(G1348), .Z(n975) );
  XNOR2_X1 U1070 ( .A(G4), .B(n975), .ZN(n976) );
  NOR2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1072 ( .A(KEYINPUT60), .B(n978), .ZN(n979) );
  NAND2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n988) );
  XNOR2_X1 U1074 ( .A(G1971), .B(G22), .ZN(n982) );
  XNOR2_X1 U1075 ( .A(G23), .B(G1976), .ZN(n981) );
  NOR2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n985) );
  XNOR2_X1 U1077 ( .A(G1986), .B(KEYINPUT125), .ZN(n983) );
  XNOR2_X1 U1078 ( .A(n983), .B(G24), .ZN(n984) );
  NAND2_X1 U1079 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1080 ( .A(KEYINPUT58), .B(n986), .ZN(n987) );
  NOR2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1083 ( .A(n991), .B(KEYINPUT61), .ZN(n992) );
  XOR2_X1 U1084 ( .A(KEYINPUT126), .B(n992), .Z(n993) );
  NAND2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1088 ( .A1(G11), .A2(n999), .ZN(n1000) );
  XNOR2_X1 U1089 ( .A(n1000), .B(KEYINPUT127), .ZN(n1029) );
  XOR2_X1 U1090 ( .A(G2072), .B(n1001), .Z(n1003) );
  XOR2_X1 U1091 ( .A(G164), .B(G2078), .Z(n1002) );
  NOR2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1093 ( .A(KEYINPUT50), .B(n1004), .Z(n1023) );
  XNOR2_X1 U1094 ( .A(G160), .B(G2084), .ZN(n1007) );
  INV_X1 U1095 ( .A(n1005), .ZN(n1006) );
  NAND2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  NAND2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1016) );
  XOR2_X1 U1099 ( .A(G2090), .B(G162), .Z(n1012) );
  NOR2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(n1014), .B(KEYINPUT51), .ZN(n1015) );
  NOR2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1018) );
  NAND2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1104 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1105 ( .A(KEYINPUT122), .B(n1021), .Z(n1022) );
  NOR2_X1 U1106 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1107 ( .A(KEYINPUT52), .B(n1024), .ZN(n1026) );
  INV_X1 U1108 ( .A(KEYINPUT55), .ZN(n1025) );
  NAND2_X1 U1109 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1110 ( .A1(n1027), .A2(G29), .ZN(n1028) );
  NAND2_X1 U1111 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1030), .Z(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
  INV_X1 U1114 ( .A(G171), .ZN(G301) );
endmodule

