//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 0 1 1 0 1 1 1 0 1 1 0 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 0 0 0 0 1 0 1 1 1 1 0 0 1 0 1 0 1 1 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1245, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1309, new_n1310, new_n1311,
    new_n1312;
  XOR2_X1   g0000(.A(KEYINPUT65), .B(G50), .Z(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT64), .ZN(new_n204));
  INV_X1    g0004(.A(KEYINPUT64), .ZN(new_n205));
  OAI21_X1  g0005(.A(new_n205), .B1(G58), .B2(G68), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n201), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT0), .ZN(new_n217));
  INV_X1    g0017(.A(G50), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n207), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n220), .A2(new_n212), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G226), .ZN(new_n223));
  INV_X1    g0023(.A(G107), .ZN(new_n224));
  INV_X1    g0024(.A(G264), .ZN(new_n225));
  OAI22_X1  g0025(.A1(new_n218), .A2(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(G116), .B2(G270), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n228));
  INV_X1    g0028(.A(G77), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT66), .B(G244), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n227), .B(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  AOI22_X1  g0031(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT67), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n214), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n217), .B(new_n222), .C1(KEYINPUT1), .C2(new_n234), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n235), .B1(KEYINPUT1), .B2(new_n234), .ZN(G361));
  XOR2_X1   g0036(.A(G238), .B(G244), .Z(new_n237));
  XNOR2_X1  g0037(.A(G226), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G250), .B(G257), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT69), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n241), .B(new_n245), .Z(G358));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XOR2_X1   g0047(.A(G50), .B(G58), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n249), .B(new_n252), .Z(G351));
  INV_X1    g0053(.A(KEYINPUT74), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G97), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT73), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(KEYINPUT73), .B1(G33), .B2(G97), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT3), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G33), .ZN(new_n263));
  INV_X1    g0063(.A(G1698), .ZN(new_n264));
  NAND4_X1  g0064(.A1(new_n261), .A2(new_n263), .A3(G226), .A4(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n259), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT3), .B(G33), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT72), .ZN(new_n268));
  NAND4_X1  g0068(.A1(new_n267), .A2(new_n268), .A3(G232), .A4(G1698), .ZN(new_n269));
  NAND4_X1  g0069(.A1(new_n261), .A2(new_n263), .A3(G232), .A4(G1698), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT72), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n266), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(G1), .A3(G13), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n254), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n274), .ZN(new_n276));
  AND2_X1   g0076(.A1(new_n271), .A2(new_n269), .ZN(new_n277));
  OAI211_X1 g0077(.A(KEYINPUT74), .B(new_n276), .C1(new_n277), .C2(new_n266), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT13), .ZN(new_n280));
  INV_X1    g0080(.A(G41), .ZN(new_n281));
  INV_X1    g0081(.A(G45), .ZN(new_n282));
  AOI21_X1  g0082(.A(G1), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(new_n274), .A3(G274), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n274), .A2(G238), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT75), .ZN(new_n288));
  XNOR2_X1  g0088(.A(new_n287), .B(new_n288), .ZN(new_n289));
  AND3_X1   g0089(.A1(new_n279), .A2(new_n280), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n280), .B1(new_n279), .B2(new_n289), .ZN(new_n291));
  OAI21_X1  g0091(.A(G169), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT14), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n279), .A2(new_n289), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT13), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n279), .A2(new_n280), .A3(new_n289), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT14), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n297), .A2(new_n298), .A3(G169), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n295), .A2(G179), .A3(new_n296), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n293), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(G20), .A2(G33), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n302), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n212), .A2(G33), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n303), .B1(new_n229), .B2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n220), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  XOR2_X1   g0108(.A(new_n308), .B(KEYINPUT76), .Z(new_n309));
  OR2_X1    g0109(.A1(new_n309), .A2(KEYINPUT11), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(KEYINPUT11), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n211), .A2(G13), .A3(G20), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT12), .B1(new_n312), .B2(G68), .ZN(new_n313));
  OR3_X1    g0113(.A1(new_n312), .A2(KEYINPUT12), .A3(G68), .ZN(new_n314));
  INV_X1    g0114(.A(new_n312), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n315), .A2(new_n307), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n203), .B1(new_n211), .B2(G20), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n313), .A2(new_n314), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n310), .A2(new_n311), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n301), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(G222), .A2(G1698), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n264), .A2(G223), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n267), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n323), .B(new_n276), .C1(G77), .C2(new_n267), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n276), .A2(new_n283), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G226), .ZN(new_n326));
  AND3_X1   g0126(.A1(new_n324), .A2(new_n284), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G179), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n329), .B1(G169), .B2(new_n327), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n211), .A2(G20), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n316), .A2(G50), .A3(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(G50), .B2(new_n312), .ZN(new_n333));
  XNOR2_X1  g0133(.A(KEYINPUT8), .B(G58), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n304), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n335), .A2(new_n336), .B1(G150), .B2(new_n302), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n337), .A2(KEYINPUT70), .B1(G20), .B2(new_n208), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(KEYINPUT70), .B2(new_n337), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n333), .B1(new_n339), .B2(new_n307), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n330), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n267), .A2(G232), .A3(new_n264), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT71), .ZN(new_n343));
  XNOR2_X1  g0143(.A(new_n342), .B(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n261), .A2(new_n263), .ZN(new_n345));
  INV_X1    g0145(.A(G238), .ZN(new_n346));
  NOR3_X1   g0146(.A1(new_n345), .A2(new_n346), .A3(new_n264), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n347), .B1(G107), .B2(new_n345), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n274), .B1(new_n344), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n274), .A2(new_n285), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n284), .B1(new_n230), .B2(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n328), .ZN(new_n353));
  INV_X1    g0153(.A(new_n307), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n335), .A2(new_n302), .B1(G20), .B2(G77), .ZN(new_n355));
  XOR2_X1   g0155(.A(KEYINPUT15), .B(G87), .Z(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n336), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n354), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n316), .A2(G77), .A3(new_n331), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(G77), .B2(new_n312), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(G169), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(new_n349), .B2(new_n351), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n353), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n352), .A2(G190), .ZN(new_n366));
  OAI21_X1  g0166(.A(G200), .B1(new_n349), .B2(new_n351), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(new_n361), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(G200), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n327), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n371), .B1(G190), .B2(new_n327), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT9), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n340), .A2(new_n373), .ZN(new_n374));
  AOI211_X1 g0174(.A(KEYINPUT9), .B(new_n333), .C1(new_n339), .C2(new_n307), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n372), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT10), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT10), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n372), .B(new_n378), .C1(new_n374), .C2(new_n375), .ZN(new_n379));
  AOI211_X1 g0179(.A(new_n341), .B(new_n369), .C1(new_n377), .C2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n297), .A2(G200), .ZN(new_n381));
  INV_X1    g0181(.A(new_n319), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n295), .A2(G190), .A3(new_n296), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n334), .B1(new_n211), .B2(G20), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n385), .A2(new_n316), .B1(new_n315), .B2(new_n334), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT7), .B1(new_n345), .B2(new_n212), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT7), .ZN(new_n389));
  AOI211_X1 g0189(.A(new_n389), .B(G20), .C1(new_n261), .C2(new_n263), .ZN(new_n390));
  OAI21_X1  g0190(.A(G68), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(G159), .ZN(new_n392));
  NOR3_X1   g0192(.A1(new_n392), .A2(G20), .A3(G33), .ZN(new_n393));
  NAND2_X1  g0193(.A1(G58), .A2(G68), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n204), .A2(new_n206), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n393), .B1(new_n395), .B2(G20), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n391), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT16), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n354), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI211_X1 g0199(.A(new_n398), .B(new_n393), .C1(new_n395), .C2(G20), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT77), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(new_n262), .B2(G33), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n260), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(new_n263), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n404), .A2(new_n389), .A3(new_n212), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(G68), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n389), .B1(new_n404), .B2(new_n212), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n400), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n387), .B1(new_n399), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(G190), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n274), .A2(G232), .A3(new_n285), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n284), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G33), .A2(G87), .ZN(new_n413));
  OR2_X1    g0213(.A1(G223), .A2(G1698), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n223), .A2(G1698), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n413), .B1(new_n404), .B2(new_n416), .ZN(new_n417));
  AOI211_X1 g0217(.A(new_n410), .B(new_n412), .C1(new_n276), .C2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n276), .ZN(new_n419));
  INV_X1    g0219(.A(new_n412), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n370), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n409), .A2(KEYINPUT79), .A3(KEYINPUT17), .A4(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n389), .B1(new_n267), .B2(G20), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n345), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n203), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n395), .A2(G20), .ZN(new_n427));
  INV_X1    g0227(.A(new_n393), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n398), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n430), .A2(new_n408), .A3(new_n307), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n422), .A2(new_n431), .A3(KEYINPUT79), .A4(new_n386), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT17), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n423), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n419), .A2(new_n420), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(G169), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n419), .A2(G179), .A3(new_n420), .ZN(new_n438));
  AOI221_X4 g0238(.A(KEYINPUT18), .B1(new_n437), .B2(new_n438), .C1(new_n431), .C2(new_n386), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT18), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n431), .A2(new_n386), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n437), .A2(new_n438), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT78), .B1(new_n439), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n442), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT18), .B1(new_n409), .B2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT78), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n441), .A2(new_n440), .A3(new_n442), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n435), .B1(new_n444), .B2(new_n449), .ZN(new_n450));
  AND4_X1   g0250(.A1(new_n320), .A2(new_n380), .A3(new_n384), .A4(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n402), .A2(new_n403), .A3(new_n212), .A4(new_n263), .ZN(new_n452));
  NAND2_X1  g0252(.A1(KEYINPUT22), .A2(G87), .ZN(new_n453));
  OR2_X1    g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n224), .A2(G20), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT90), .B1(new_n455), .B2(KEYINPUT23), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT90), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT23), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n457), .A2(new_n458), .A3(new_n224), .A4(G20), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n212), .A2(G33), .A3(G116), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n456), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  OR2_X1    g0262(.A1(KEYINPUT88), .A2(KEYINPUT23), .ZN(new_n463));
  NAND2_X1  g0263(.A1(KEYINPUT88), .A2(KEYINPUT23), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(new_n455), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT89), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT89), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n463), .A2(new_n455), .A3(new_n467), .A4(new_n464), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n267), .A2(new_n212), .A3(G87), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT22), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n454), .A2(new_n462), .A3(new_n469), .A4(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(KEYINPUT24), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n461), .B1(new_n471), .B2(new_n470), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT24), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n475), .A2(new_n476), .A3(new_n454), .A4(new_n469), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n307), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n315), .A2(KEYINPUT25), .A3(new_n224), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(KEYINPUT91), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT25), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(new_n312), .B2(G107), .ZN(new_n483));
  OR2_X1    g0283(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n481), .A2(new_n483), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n211), .A2(G33), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n312), .A2(new_n486), .A3(new_n220), .A4(new_n306), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n484), .A2(new_n485), .B1(G107), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n479), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT93), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT92), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n211), .A2(G45), .ZN(new_n493));
  OR2_X1    g0293(.A1(KEYINPUT5), .A2(G41), .ZN(new_n494));
  NAND2_X1  g0294(.A1(KEYINPUT5), .A2(G41), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n496), .A2(new_n276), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n492), .B1(new_n497), .B2(G264), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n282), .A2(G1), .ZN(new_n499));
  INV_X1    g0299(.A(new_n495), .ZN(new_n500));
  NOR2_X1   g0300(.A1(KEYINPUT5), .A2(G41), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n502), .A2(new_n492), .A3(G264), .A4(new_n274), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n491), .B1(new_n498), .B2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(G257), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G1698), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n507), .B1(G250), .B2(G1698), .ZN(new_n508));
  INV_X1    g0308(.A(G294), .ZN(new_n509));
  OAI22_X1  g0309(.A1(new_n404), .A2(new_n508), .B1(new_n260), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n274), .A2(G274), .ZN(new_n511));
  OAI21_X1  g0311(.A(KEYINPUT82), .B1(new_n511), .B2(new_n502), .ZN(new_n512));
  INV_X1    g0312(.A(G274), .ZN(new_n513));
  INV_X1    g0313(.A(new_n220), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n513), .B1(new_n514), .B2(new_n273), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT82), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n496), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n276), .A2(new_n510), .B1(new_n512), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n502), .A2(new_n274), .ZN(new_n519));
  OAI21_X1  g0319(.A(KEYINPUT92), .B1(new_n519), .B2(new_n225), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n520), .A2(KEYINPUT93), .A3(new_n503), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n505), .A2(new_n518), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n503), .ZN(new_n523));
  AND2_X1   g0323(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n522), .A2(new_n370), .B1(new_n524), .B2(new_n410), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n490), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g0326(.A(new_n493), .B(KEYINPUT84), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n274), .A2(G250), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n527), .A2(new_n528), .B1(new_n515), .B2(new_n499), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n402), .A2(new_n403), .A3(G244), .A4(new_n263), .ZN(new_n530));
  INV_X1    g0330(.A(G116), .ZN(new_n531));
  OAI22_X1  g0331(.A1(new_n530), .A2(new_n264), .B1(new_n260), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n346), .A2(G1698), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n402), .A2(new_n403), .A3(new_n533), .A4(new_n263), .ZN(new_n534));
  OR2_X1    g0334(.A1(new_n534), .A2(KEYINPUT85), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(KEYINPUT85), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n532), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n328), .B(new_n529), .C1(new_n537), .C2(new_n274), .ZN(new_n538));
  INV_X1    g0338(.A(G97), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n304), .A2(new_n539), .ZN(new_n540));
  OAI22_X1  g0340(.A1(new_n452), .A2(new_n203), .B1(KEYINPUT19), .B2(new_n540), .ZN(new_n541));
  NOR3_X1   g0341(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n542));
  OAI21_X1  g0342(.A(KEYINPUT19), .B1(new_n257), .B2(new_n258), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n542), .B1(new_n543), .B2(new_n212), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n307), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n356), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n315), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n545), .B(new_n547), .C1(new_n546), .C2(new_n487), .ZN(new_n548));
  INV_X1    g0348(.A(new_n529), .ZN(new_n549));
  XNOR2_X1  g0349(.A(new_n534), .B(KEYINPUT85), .ZN(new_n550));
  INV_X1    g0350(.A(new_n532), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n549), .B1(new_n552), .B2(new_n276), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n538), .B(new_n548), .C1(new_n553), .C2(G169), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n488), .A2(G87), .ZN(new_n555));
  AND3_X1   g0355(.A1(new_n545), .A2(new_n547), .A3(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(G190), .B(new_n529), .C1(new_n537), .C2(new_n274), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n556), .B(new_n557), .C1(new_n553), .C2(new_n370), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n526), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n497), .A2(KEYINPUT83), .A3(G257), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT83), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(new_n519), .B2(new_n506), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n561), .A2(new_n563), .B1(new_n517), .B2(new_n512), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT4), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n530), .B2(G1698), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n267), .A2(G250), .A3(G1698), .ZN(new_n567));
  AND2_X1   g0367(.A1(KEYINPUT4), .A2(G244), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n261), .A2(new_n263), .A3(new_n568), .A4(new_n264), .ZN(new_n569));
  NAND2_X1  g0369(.A1(G33), .A2(G283), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(KEYINPUT80), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT80), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n572), .A2(G33), .A3(G283), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n566), .A2(new_n567), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n576), .A2(KEYINPUT81), .A3(new_n276), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT81), .B1(new_n576), .B2(new_n276), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n564), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(G200), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n302), .A2(G77), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT6), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n583), .A2(new_n539), .A3(G107), .ZN(new_n584));
  XNOR2_X1  g0384(.A(G97), .B(G107), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n584), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n582), .B1(new_n586), .B2(new_n212), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n224), .B1(new_n424), .B2(new_n425), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n307), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n315), .A2(new_n539), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(new_n487), .B2(new_n539), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n576), .A2(new_n276), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n564), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n593), .B1(new_n595), .B2(G190), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n328), .B(new_n564), .C1(new_n578), .C2(new_n579), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n564), .A2(new_n594), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n598), .A2(new_n363), .B1(new_n589), .B2(new_n592), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n581), .A2(new_n596), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n560), .A2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT20), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n212), .B1(new_n539), .B2(G33), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n603), .B1(new_n571), .B2(new_n573), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n306), .A2(new_n220), .B1(G20), .B2(new_n531), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n602), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n571), .A2(new_n573), .ZN(new_n608));
  OAI211_X1 g0408(.A(KEYINPUT20), .B(new_n605), .C1(new_n608), .C2(new_n603), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT86), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n312), .A2(G116), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n612), .B1(new_n488), .B2(G116), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n611), .B1(new_n610), .B2(new_n613), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n512), .A2(new_n517), .B1(new_n497), .B2(G270), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n225), .A2(G1698), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n618), .B1(G257), .B2(G1698), .ZN(new_n619));
  INV_X1    g0419(.A(G303), .ZN(new_n620));
  OAI22_X1  g0420(.A1(new_n404), .A2(new_n619), .B1(new_n620), .B2(new_n267), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n276), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n617), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(G200), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n616), .B(new_n624), .C1(new_n410), .C2(new_n623), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n511), .A2(new_n502), .A3(KEYINPUT82), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n516), .B1(new_n496), .B2(new_n515), .ZN(new_n627));
  INV_X1    g0427(.A(G270), .ZN(new_n628));
  OAI22_X1  g0428(.A1(new_n626), .A2(new_n627), .B1(new_n628), .B2(new_n519), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n621), .A2(new_n276), .ZN(new_n630));
  OAI21_X1  g0430(.A(G169), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n610), .A2(new_n613), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(KEYINPUT86), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n631), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT87), .ZN(new_n636));
  OAI21_X1  g0436(.A(KEYINPUT21), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n505), .A2(G179), .A3(new_n518), .A4(new_n521), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n518), .A2(new_n523), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(G169), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n354), .B1(new_n474), .B2(new_n477), .ZN(new_n642));
  INV_X1    g0442(.A(new_n489), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT21), .ZN(new_n645));
  OAI211_X1 g0445(.A(KEYINPUT87), .B(new_n645), .C1(new_n616), .C2(new_n631), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n633), .A2(new_n634), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n623), .A2(new_n328), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n637), .A2(new_n644), .A3(new_n646), .A4(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n601), .A2(new_n625), .A3(new_n651), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n451), .A2(new_n652), .ZN(G372));
  NOR2_X1   g0453(.A1(new_n439), .A2(new_n443), .ZN(new_n654));
  INV_X1    g0454(.A(new_n365), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n301), .A2(new_n319), .B1(new_n384), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n654), .B1(new_n656), .B2(new_n435), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n377), .A2(new_n379), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n341), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n560), .A2(new_n650), .A3(new_n600), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n599), .A2(new_n597), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n661), .A2(KEYINPUT26), .A3(new_n554), .A4(new_n558), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT26), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n599), .A2(new_n597), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n663), .B1(new_n559), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g0466(.A(new_n554), .B(KEYINPUT94), .Z(new_n667));
  NAND3_X1  g0467(.A1(new_n660), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n451), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n659), .A2(new_n669), .ZN(G369));
  NOR2_X1   g0470(.A1(new_n642), .A2(new_n643), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n211), .A2(new_n212), .A3(G13), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G213), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(G343), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  OR3_X1    g0478(.A1(new_n671), .A2(KEYINPUT95), .A3(new_n678), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n490), .A2(new_n525), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT95), .B1(new_n671), .B2(new_n678), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n679), .A2(new_n680), .A3(new_n644), .A4(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n637), .A2(new_n646), .A3(new_n649), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n678), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n677), .B(KEYINPUT96), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  OAI22_X1  g0486(.A1(new_n682), .A2(new_n684), .B1(new_n644), .B2(new_n686), .ZN(new_n687));
  XOR2_X1   g0487(.A(new_n687), .B(KEYINPUT97), .Z(new_n688));
  NOR2_X1   g0488(.A1(new_n616), .A2(new_n678), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n683), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n625), .ZN(new_n691));
  INV_X1    g0491(.A(G330), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n682), .B1(new_n644), .B2(new_n678), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n688), .A2(new_n695), .ZN(G399));
  INV_X1    g0496(.A(new_n215), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(G41), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n542), .A2(new_n531), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n699), .A2(G1), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n219), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n702), .B1(new_n703), .B2(new_n699), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT28), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT31), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n328), .B1(new_n629), .B2(new_n630), .ZN(new_n707));
  AND3_X1   g0507(.A1(new_n520), .A2(KEYINPUT93), .A3(new_n503), .ZN(new_n708));
  AOI21_X1  g0508(.A(KEYINPUT93), .B1(new_n520), .B2(new_n503), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n707), .B1(new_n710), .B2(new_n518), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT98), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n529), .B1(new_n537), .B2(new_n274), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n711), .A2(new_n712), .A3(new_n580), .A4(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(G179), .B1(new_n617), .B2(new_n622), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n522), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n561), .A2(new_n563), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n512), .A2(new_n517), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT81), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n594), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n719), .B1(new_n721), .B2(new_n577), .ZN(new_n722));
  OAI21_X1  g0522(.A(KEYINPUT98), .B1(new_n716), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n714), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT30), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n510), .A2(new_n276), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n648), .A2(new_n710), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n595), .A2(new_n553), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n725), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n710), .A2(new_n726), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n598), .A2(new_n713), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n730), .A2(KEYINPUT30), .A3(new_n648), .A4(new_n731), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n724), .A2(KEYINPUT99), .A3(new_n729), .A4(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(new_n677), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n732), .A2(new_n729), .ZN(new_n735));
  AOI21_X1  g0535(.A(KEYINPUT99), .B1(new_n735), .B2(new_n724), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n706), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n601), .A2(new_n651), .A3(new_n625), .A4(new_n685), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n732), .A2(new_n729), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n716), .A2(new_n722), .ZN(new_n741));
  OAI211_X1 g0541(.A(KEYINPUT31), .B(new_n686), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n692), .B1(new_n739), .B2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT29), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n744), .B1(new_n668), .B2(new_n678), .ZN(new_n745));
  AND3_X1   g0545(.A1(new_n668), .A2(new_n744), .A3(new_n685), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n743), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n705), .B1(new_n747), .B2(G1), .ZN(G364));
  AND2_X1   g0548(.A1(new_n212), .A2(G13), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n211), .B1(new_n749), .B2(G45), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n698), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n693), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(G330), .B1(new_n690), .B2(new_n625), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G13), .A2(G33), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n691), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n215), .A2(new_n267), .ZN(new_n760));
  INV_X1    g0560(.A(G355), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n760), .A2(new_n761), .B1(G116), .B2(new_n215), .ZN(new_n762));
  INV_X1    g0562(.A(new_n404), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n697), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n765), .B1(new_n282), .B2(new_n219), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n249), .A2(G45), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n762), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n514), .B1(new_n212), .B2(G169), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n769), .A2(KEYINPUT100), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(KEYINPUT100), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n758), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n752), .B1(new_n768), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n212), .A2(new_n328), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n776), .A2(G190), .A3(new_n370), .ZN(new_n777));
  INV_X1    g0577(.A(G322), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G190), .A2(G200), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G311), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n777), .A2(new_n778), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n212), .A2(G179), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(new_n779), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n267), .B(new_n782), .C1(G329), .C2(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n776), .A2(new_n410), .A3(G200), .ZN(new_n787));
  AND2_X1   g0587(.A1(new_n787), .A2(KEYINPUT102), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n787), .A2(KEYINPUT102), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(KEYINPUT33), .B(G317), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n410), .A2(G179), .A3(G200), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n212), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n783), .A2(G190), .A3(G200), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n796), .A2(G294), .B1(new_n798), .B2(G303), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n776), .A2(G200), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n410), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n783), .A2(new_n410), .A3(G200), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n801), .A2(G326), .B1(new_n803), .B2(G283), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n786), .A2(new_n793), .A3(new_n799), .A4(new_n804), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n790), .A2(new_n203), .B1(new_n539), .B2(new_n795), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n806), .B(KEYINPUT103), .Z(new_n807));
  XOR2_X1   g0607(.A(new_n777), .B(KEYINPUT101), .Z(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G58), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n784), .A2(new_n392), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT32), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n802), .A2(new_n224), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(G87), .B2(new_n798), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n267), .B1(new_n780), .B2(new_n229), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n815), .B1(G50), .B2(new_n801), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n810), .A2(new_n812), .A3(new_n814), .A4(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n805), .B1(new_n807), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n775), .B1(new_n818), .B2(new_n772), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n753), .A2(new_n755), .B1(new_n759), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(G396));
  INV_X1    g0621(.A(new_n752), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n772), .A2(new_n756), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n822), .B1(new_n823), .B2(new_n229), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n368), .B1(new_n361), .B2(new_n678), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n365), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n655), .A2(new_n678), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n780), .ZN(new_n830));
  AOI22_X1  g0630(.A1(G116), .A2(new_n830), .B1(new_n785), .B2(G311), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n831), .B(new_n345), .C1(new_n509), .C2(new_n777), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n801), .A2(G303), .B1(new_n798), .B2(G107), .ZN(new_n833));
  INV_X1    g0633(.A(G87), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n833), .B1(new_n834), .B2(new_n802), .C1(new_n539), .C2(new_n795), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n832), .B(new_n835), .C1(G283), .C2(new_n791), .ZN(new_n836));
  INV_X1    g0636(.A(G132), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n763), .B1(new_n837), .B2(new_n784), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n796), .A2(G58), .B1(new_n803), .B2(G68), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n218), .B2(new_n797), .ZN(new_n840));
  INV_X1    g0640(.A(G150), .ZN(new_n841));
  INV_X1    g0641(.A(G137), .ZN(new_n842));
  INV_X1    g0642(.A(new_n801), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n790), .A2(new_n841), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT104), .ZN(new_n845));
  INV_X1    g0645(.A(G143), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n845), .B1(new_n846), .B2(new_n808), .C1(new_n392), .C2(new_n780), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n838), .B(new_n840), .C1(new_n848), .C2(KEYINPUT34), .ZN(new_n849));
  OR2_X1    g0649(.A1(new_n848), .A2(KEYINPUT34), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n836), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n772), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n824), .B1(new_n829), .B2(new_n757), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n743), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n668), .A2(new_n685), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(new_n829), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n822), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n858), .A2(KEYINPUT105), .B1(new_n854), .B2(new_n856), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n858), .A2(KEYINPUT105), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n853), .B1(new_n860), .B2(new_n861), .ZN(G384));
  NAND2_X1  g0662(.A1(new_n855), .A2(new_n829), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n827), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n319), .A2(new_n677), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n320), .A2(new_n384), .A3(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n384), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n319), .B(new_n677), .C1(new_n867), .C2(new_n301), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n864), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n409), .A2(new_n422), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n441), .A2(new_n442), .ZN(new_n873));
  INV_X1    g0673(.A(new_n675), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n441), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n872), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  OR2_X1    g0676(.A1(new_n876), .A2(KEYINPUT37), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n408), .A2(new_n307), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n396), .B1(new_n406), .B2(new_n407), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n398), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n387), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n872), .B1(new_n445), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n881), .A2(new_n675), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT37), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n877), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT106), .ZN(new_n887));
  INV_X1    g0687(.A(new_n435), .ZN(new_n888));
  NOR3_X1   g0688(.A1(new_n439), .A2(new_n443), .A3(KEYINPUT78), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n447), .B1(new_n446), .B2(new_n448), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n887), .B1(new_n891), .B2(new_n883), .ZN(new_n892));
  INV_X1    g0692(.A(new_n883), .ZN(new_n893));
  NOR3_X1   g0693(.A1(new_n450), .A2(KEYINPUT106), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n886), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT38), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n891), .A2(new_n887), .A3(new_n883), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT106), .B1(new_n450), .B2(new_n893), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n885), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(KEYINPUT38), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n897), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n654), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n871), .A2(new_n902), .B1(new_n903), .B2(new_n675), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n441), .B(new_n874), .C1(new_n903), .C2(new_n435), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n876), .B(KEYINPUT37), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT38), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n901), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g0709(.A(KEYINPUT108), .B(KEYINPUT39), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n900), .A2(KEYINPUT38), .ZN(new_n912));
  AOI211_X1 g0712(.A(new_n896), .B(new_n885), .C1(new_n898), .C2(new_n899), .ZN(new_n913));
  OAI21_X1  g0713(.A(KEYINPUT39), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT107), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n902), .A2(KEYINPUT107), .A3(KEYINPUT39), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n911), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n301), .A2(new_n319), .A3(new_n678), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n904), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n451), .B1(new_n746), .B2(new_n745), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n659), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n922), .B(KEYINPUT109), .Z(new_n923));
  XNOR2_X1  g0723(.A(new_n920), .B(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT99), .ZN(new_n925));
  INV_X1    g0725(.A(new_n724), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n925), .B1(new_n926), .B2(new_n740), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n927), .A2(KEYINPUT31), .A3(new_n677), .A4(new_n733), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n737), .A2(new_n738), .A3(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n929), .A2(new_n829), .A3(new_n869), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n907), .B1(new_n900), .B2(KEYINPUT38), .ZN(new_n931));
  OAI21_X1  g0731(.A(KEYINPUT40), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT40), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n912), .B2(new_n913), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n932), .B1(new_n930), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n929), .A2(new_n451), .ZN(new_n937));
  OAI21_X1  g0737(.A(G330), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(new_n937), .B2(new_n936), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n924), .A2(new_n939), .B1(new_n211), .B2(new_n749), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(new_n924), .B2(new_n939), .ZN(new_n941));
  INV_X1    g0741(.A(new_n586), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n942), .A2(KEYINPUT35), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(KEYINPUT35), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n943), .A2(G116), .A3(new_n221), .A4(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT36), .Z(new_n946));
  NAND3_X1  g0746(.A1(new_n219), .A2(G77), .A3(new_n394), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n201), .A2(G68), .ZN(new_n948));
  AOI211_X1 g0748(.A(new_n211), .B(G13), .C1(new_n947), .C2(new_n948), .ZN(new_n949));
  OR3_X1    g0749(.A1(new_n941), .A2(new_n946), .A3(new_n949), .ZN(G367));
  AOI21_X1  g0750(.A(new_n774), .B1(new_n697), .B2(new_n356), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n245), .A2(new_n764), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n822), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT114), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n830), .A2(G283), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT46), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n797), .B2(new_n531), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n785), .A2(G317), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n955), .A2(new_n957), .A3(new_n958), .A4(new_n404), .ZN(new_n959));
  NOR3_X1   g0759(.A1(new_n797), .A2(new_n956), .A3(new_n531), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n959), .B(new_n960), .C1(new_n809), .C2(G303), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n791), .A2(G294), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n803), .A2(G97), .ZN(new_n963));
  AOI22_X1  g0763(.A1(G107), .A2(new_n796), .B1(new_n801), .B2(G311), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n961), .A2(new_n962), .A3(new_n963), .A4(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n790), .A2(new_n392), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n201), .A2(new_n780), .B1(new_n784), .B2(new_n842), .ZN(new_n967));
  INV_X1    g0767(.A(new_n777), .ZN(new_n968));
  AOI211_X1 g0768(.A(new_n345), .B(new_n967), .C1(G150), .C2(new_n968), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n796), .A2(G68), .B1(new_n803), .B2(G77), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n801), .A2(G143), .B1(new_n798), .B2(G58), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n965), .B1(new_n966), .B2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n974), .A2(KEYINPUT47), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT47), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n772), .B1(new_n973), .B2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n667), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n556), .A2(new_n678), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n559), .A2(new_n979), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n758), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n954), .B1(new_n975), .B2(new_n977), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n686), .A2(new_n593), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n600), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n661), .A2(new_n686), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OR3_X1    g0788(.A1(new_n688), .A2(KEYINPUT112), .A3(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(KEYINPUT112), .B1(new_n688), .B2(new_n988), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT44), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n688), .A2(new_n988), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT45), .Z(new_n995));
  NAND3_X1  g0795(.A1(new_n989), .A2(KEYINPUT44), .A3(new_n990), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n993), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n695), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT113), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n999), .A2(KEYINPUT113), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n682), .A2(new_n684), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n684), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1004), .B1(new_n694), .B2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n693), .B(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n747), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n993), .A2(new_n995), .A3(new_n695), .A4(new_n996), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1002), .A2(new_n1003), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n747), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n698), .B(KEYINPUT41), .Z(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n751), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n988), .B(KEYINPUT110), .Z(new_n1016));
  NOR2_X1   g0816(.A1(new_n695), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT111), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1018), .B(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1004), .B1(new_n986), .B2(new_n987), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT42), .Z(new_n1023));
  OR2_X1    g0823(.A1(new_n1016), .A2(new_n644), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n686), .B1(new_n1024), .B2(new_n664), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1021), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1020), .B(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n984), .B1(new_n1015), .B2(new_n1028), .ZN(G387));
  NOR2_X1   g0829(.A1(new_n1009), .A2(new_n699), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n747), .B2(new_n1007), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n694), .A2(new_n983), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n760), .A2(new_n701), .B1(G107), .B2(new_n215), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n241), .A2(new_n282), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n334), .A2(G50), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT50), .ZN(new_n1036));
  AOI211_X1 g0836(.A(G45), .B(new_n700), .C1(G68), .C2(G77), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n765), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1033), .B1(new_n1034), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n752), .B1(new_n1039), .B2(new_n774), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n843), .A2(new_n392), .B1(new_n546), .B2(new_n795), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n797), .A2(new_n229), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n791), .A2(new_n335), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n777), .A2(new_n218), .B1(new_n784), .B2(new_n841), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(G68), .B2(new_n830), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n404), .B1(new_n803), .B2(G97), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1043), .A2(new_n1044), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n796), .A2(G283), .B1(new_n798), .B2(G294), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n801), .A2(G322), .B1(new_n830), .B2(G303), .ZN(new_n1050));
  INV_X1    g0850(.A(G317), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1050), .B1(new_n790), .B2(new_n781), .C1(new_n808), .C2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT48), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1049), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT115), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1055), .A2(KEYINPUT49), .A3(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n763), .B1(G326), .B2(new_n785), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1057), .B(new_n1058), .C1(new_n531), .C2(new_n802), .ZN(new_n1059));
  AOI21_X1  g0859(.A(KEYINPUT49), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1048), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1040), .B1(new_n1061), .B2(new_n772), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n1007), .A2(new_n751), .B1(new_n1032), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1031), .A2(new_n1063), .ZN(G393));
  NAND2_X1  g0864(.A1(new_n999), .A2(new_n1010), .ZN(new_n1065));
  AND3_X1   g0865(.A1(new_n1065), .A2(KEYINPUT117), .A3(new_n1008), .ZN(new_n1066));
  AOI21_X1  g0866(.A(KEYINPUT117), .B1(new_n1065), .B2(new_n1008), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1011), .B(new_n698), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1065), .A2(new_n750), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n843), .A2(new_n841), .B1(new_n392), .B2(new_n777), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT51), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n780), .A2(new_n334), .B1(new_n784), .B2(new_n846), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n203), .A2(new_n797), .B1(new_n802), .B2(new_n834), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n795), .A2(new_n229), .ZN(new_n1074));
  NOR4_X1   g0874(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .A4(new_n404), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1071), .B(new_n1075), .C1(new_n201), .C2(new_n790), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT116), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n843), .A2(new_n1051), .B1(new_n781), .B2(new_n777), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT52), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n813), .B1(G116), .B2(new_n796), .ZN(new_n1081));
  INV_X1    g0881(.A(G283), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1081), .B1(new_n1082), .B2(new_n797), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n345), .B1(new_n784), .B2(new_n778), .C1(new_n509), .C2(new_n780), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1080), .B(new_n1085), .C1(new_n620), .C2(new_n790), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1078), .A2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n772), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n765), .A2(new_n252), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n773), .B1(new_n539), .B2(new_n215), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1089), .B(new_n752), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n1016), .B2(new_n758), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1069), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1068), .A2(new_n1094), .ZN(G390));
  OR2_X1    g0895(.A1(new_n909), .A2(new_n910), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n870), .A2(new_n919), .ZN(new_n1097));
  AOI21_X1  g0897(.A(KEYINPUT107), .B1(new_n902), .B2(KEYINPUT39), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT39), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n915), .B(new_n1099), .C1(new_n897), .C2(new_n901), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1096), .B(new_n1097), .C1(new_n1098), .C2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n668), .A2(new_n678), .A3(new_n826), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n827), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n869), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n909), .A2(new_n919), .A3(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n743), .A2(new_n829), .A3(new_n869), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1101), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n929), .A2(new_n451), .A3(G330), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1108), .A2(new_n921), .A3(new_n659), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(KEYINPUT118), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT118), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1108), .A2(new_n921), .A3(new_n659), .A4(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n869), .B1(new_n743), .B2(new_n829), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n929), .A2(G330), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n869), .ZN(new_n1116));
  NOR3_X1   g0916(.A1(new_n1115), .A2(new_n1116), .A3(new_n828), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n864), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1116), .B1(new_n1115), .B2(new_n828), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1106), .A2(new_n827), .A3(new_n1119), .A4(new_n1102), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1113), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1105), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(new_n918), .B2(new_n1097), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1117), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1107), .B(new_n1121), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(KEYINPUT119), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n1117), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT119), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1128), .A2(new_n1129), .A3(new_n1107), .A4(new_n1121), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1126), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1128), .A2(new_n1107), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1121), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n699), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1128), .A2(new_n751), .A3(new_n1107), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n823), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n752), .B1(new_n1137), .B2(new_n335), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(KEYINPUT54), .B(G143), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n796), .A2(G159), .B1(new_n830), .B2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1141), .B1(new_n790), .B2(new_n842), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT120), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n797), .A2(new_n841), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT53), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n968), .A2(G132), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n345), .B1(new_n785), .B2(G125), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n201), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(G128), .A2(new_n801), .B1(new_n1148), .B2(new_n803), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .A4(new_n1149), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n790), .A2(new_n224), .B1(new_n539), .B2(new_n780), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT121), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n345), .B1(new_n777), .B2(new_n531), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(G294), .B2(new_n785), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n203), .A2(new_n802), .B1(new_n797), .B2(new_n834), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n1074), .B(new_n1156), .C1(G283), .C2(new_n801), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1153), .A2(new_n1155), .A3(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n1143), .A2(new_n1150), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1138), .B1(new_n1160), .B2(new_n772), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1096), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1161), .B1(new_n1162), .B2(new_n757), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1135), .A2(new_n1136), .A3(new_n1163), .ZN(G378));
  AOI21_X1  g0964(.A(new_n1113), .B1(new_n1126), .B2(new_n1130), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n341), .B1(new_n377), .B2(new_n379), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n340), .A2(new_n675), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT55), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1166), .B(new_n1168), .ZN(new_n1169));
  XOR2_X1   g0969(.A(KEYINPUT122), .B(KEYINPUT56), .Z(new_n1170));
  XOR2_X1   g0970(.A(new_n1169), .B(new_n1170), .Z(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n935), .A2(G330), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1173), .B(new_n904), .C1(new_n918), .C2(new_n919), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n919), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1162), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1173), .B1(new_n1177), .B2(new_n904), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1172), .B1(new_n1175), .B2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n920), .A2(G330), .A3(new_n935), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1180), .A2(new_n1174), .A3(new_n1171), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1179), .A2(KEYINPUT57), .A3(new_n1181), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n1165), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT57), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1184), .B1(new_n1165), .B2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1183), .A2(new_n698), .A3(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n752), .B1(new_n1137), .B2(new_n1148), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n803), .A2(G58), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n843), .B2(new_n531), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1042), .B(new_n1190), .C1(G68), .C2(new_n796), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n404), .A2(new_n281), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n777), .A2(new_n224), .B1(new_n784), .B2(new_n1082), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1192), .B(new_n1193), .C1(new_n356), .C2(new_n830), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1191), .B(new_n1194), .C1(new_n539), .C2(new_n790), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT58), .ZN(new_n1196));
  AOI21_X1  g0996(.A(G50), .B1(new_n260), .B2(new_n281), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1195), .A2(new_n1196), .B1(new_n1192), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(G128), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n777), .A2(new_n1199), .B1(new_n780), .B2(new_n842), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(G150), .B2(new_n796), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n801), .A2(G125), .B1(new_n798), .B2(new_n1140), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1201), .B(new_n1202), .C1(new_n790), .C2(new_n837), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1203), .A2(KEYINPUT59), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(KEYINPUT59), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n803), .A2(G159), .ZN(new_n1206));
  AOI211_X1 g1006(.A(G33), .B(G41), .C1(new_n785), .C2(G124), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1198), .B1(new_n1196), .B2(new_n1195), .C1(new_n1204), .C2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1188), .B1(new_n1209), .B2(new_n772), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n1171), .B2(new_n757), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT123), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1185), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1212), .B1(new_n1213), .B2(new_n751), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1187), .A2(new_n1214), .ZN(G375));
  NAND2_X1  g1015(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1116), .A2(new_n756), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n752), .B1(new_n1137), .B2(G68), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n791), .A2(G116), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n780), .A2(new_n224), .B1(new_n784), .B2(new_n620), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n267), .B(new_n1220), .C1(G283), .C2(new_n968), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n796), .A2(new_n356), .B1(new_n803), .B2(G77), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n801), .A2(G294), .B1(new_n798), .B2(G97), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1219), .A2(new_n1221), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n808), .A2(new_n842), .B1(new_n837), .B2(new_n843), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n791), .B2(new_n1140), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n1226), .A2(KEYINPUT124), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1189), .B1(new_n392), .B2(new_n797), .C1(new_n218), .C2(new_n795), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n780), .A2(new_n841), .B1(new_n784), .B2(new_n1199), .ZN(new_n1229));
  NOR3_X1   g1029(.A1(new_n1228), .A2(new_n404), .A3(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n1226), .B2(KEYINPUT124), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1224), .B1(new_n1227), .B2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1218), .B1(new_n1232), .B2(new_n772), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1216), .A2(new_n751), .B1(new_n1217), .B2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1133), .A2(new_n1014), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1113), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1216), .A2(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1234), .B1(new_n1235), .B2(new_n1237), .ZN(G381));
  NOR2_X1   g1038(.A1(G393), .A2(G396), .ZN(new_n1239));
  INV_X1    g1039(.A(G384), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NOR4_X1   g1041(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1241), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(G375), .A2(G378), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(G407));
  OAI21_X1  g1044(.A(new_n1243), .B1(new_n1242), .B2(new_n676), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(G213), .ZN(G409));
  INV_X1    g1046(.A(KEYINPUT126), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1131), .A2(new_n1236), .ZN(new_n1248));
  AOI21_X1  g1048(.A(KEYINPUT57), .B1(new_n1248), .B2(new_n1213), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n698), .B1(new_n1165), .B2(new_n1182), .ZN(new_n1250));
  OAI211_X1 g1050(.A(G378), .B(new_n1214), .C1(new_n1249), .C2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(KEYINPUT125), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT125), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1187), .A2(new_n1253), .A3(G378), .A4(new_n1214), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1213), .A2(new_n751), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1256), .A2(new_n1211), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1248), .A2(new_n1213), .A3(new_n1014), .ZN(new_n1258));
  AOI21_X1  g1058(.A(G378), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1255), .A2(new_n1260), .ZN(new_n1261));
  AND2_X1   g1061(.A1(new_n1133), .A2(KEYINPUT60), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n699), .B1(new_n1262), .B2(new_n1237), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1263), .B1(new_n1237), .B2(new_n1262), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n1234), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1240), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1264), .A2(G384), .A3(new_n1234), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n676), .A2(G213), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1261), .A2(KEYINPUT63), .A3(new_n1269), .A4(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1270), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(G2897), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1268), .B(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1259), .B1(new_n1252), .B2(new_n1254), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1274), .B1(new_n1275), .B2(new_n1272), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT61), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1271), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  OR2_X1    g1078(.A1(new_n1015), .A2(new_n1028), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n820), .B1(new_n1031), .B2(new_n1063), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1239), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(G390), .A2(new_n1281), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1068), .B(new_n1094), .C1(new_n1239), .C2(new_n1280), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1279), .A2(new_n984), .A3(new_n1282), .A4(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(G387), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1284), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  NOR3_X1   g1088(.A1(new_n1275), .A2(new_n1268), .A3(new_n1272), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1288), .B1(new_n1289), .B2(KEYINPUT63), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1247), .B1(new_n1278), .B2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1261), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT63), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1287), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1261), .A2(new_n1270), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT61), .B1(new_n1295), .B2(new_n1274), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1294), .A2(new_n1296), .A3(KEYINPUT126), .A4(new_n1271), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1291), .A2(new_n1297), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1289), .A2(KEYINPUT62), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT62), .ZN(new_n1300));
  NOR4_X1   g1100(.A1(new_n1275), .A2(new_n1300), .A3(new_n1268), .A4(new_n1272), .ZN(new_n1301));
  OAI211_X1 g1101(.A(new_n1296), .B(KEYINPUT127), .C1(new_n1299), .C2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1287), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1301), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1292), .A2(new_n1300), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(KEYINPUT127), .B1(new_n1306), .B2(new_n1296), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1298), .B1(new_n1303), .B2(new_n1307), .ZN(G405));
  INV_X1    g1108(.A(G378), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(G375), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1255), .A2(new_n1310), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(new_n1311), .B(new_n1268), .ZN(new_n1312));
  XNOR2_X1  g1112(.A(new_n1312), .B(new_n1288), .ZN(G402));
endmodule


