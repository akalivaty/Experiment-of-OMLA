//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 1 1 0 1 1 0 1 0 0 1 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 0 0 0 1 1 0 0 0 1 0 1 0 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985;
  INV_X1    g000(.A(G119), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G116), .ZN(new_n188));
  INV_X1    g002(.A(G116), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G119), .ZN(new_n190));
  INV_X1    g004(.A(G113), .ZN(new_n191));
  AND2_X1   g005(.A1(new_n191), .A2(KEYINPUT2), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n191), .A2(KEYINPUT2), .ZN(new_n193));
  OAI211_X1 g007(.A(new_n188), .B(new_n190), .C1(new_n192), .C2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n188), .A2(new_n190), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT2), .B(G113), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT67), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n194), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n195), .A2(new_n196), .A3(KEYINPUT67), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT4), .ZN(new_n203));
  INV_X1    g017(.A(G107), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(G104), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n206));
  INV_X1    g020(.A(G104), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(G107), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n204), .A2(KEYINPUT3), .A3(G104), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n205), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G101), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n203), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI211_X1 g026(.A(KEYINPUT78), .B(new_n205), .C1(new_n208), .C2(new_n209), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT78), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n208), .A2(new_n209), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n207), .A2(G107), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n213), .A2(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n212), .B1(new_n218), .B2(G101), .ZN(new_n219));
  AND3_X1   g033(.A1(new_n204), .A2(KEYINPUT3), .A3(G104), .ZN(new_n220));
  AOI21_X1  g034(.A(KEYINPUT3), .B1(new_n204), .B2(G104), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n216), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT78), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n210), .A2(new_n214), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n223), .A2(KEYINPUT4), .A3(new_n224), .A4(G101), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n202), .B1(new_n219), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n204), .A2(G104), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n228), .B1(new_n216), .B2(KEYINPUT79), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT79), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n205), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(G101), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n210), .A2(new_n211), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT5), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n235), .B(G113), .C1(KEYINPUT5), .C2(new_n188), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(new_n194), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  XOR2_X1   g053(.A(G110), .B(G122), .Z(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n227), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n223), .A2(G101), .A3(new_n224), .ZN(new_n243));
  INV_X1    g057(.A(new_n212), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n201), .B1(new_n245), .B2(new_n225), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n240), .B1(new_n246), .B2(new_n238), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n242), .A2(new_n247), .A3(KEYINPUT6), .ZN(new_n248));
  XNOR2_X1  g062(.A(G143), .B(G146), .ZN(new_n249));
  INV_X1    g063(.A(G128), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n250), .A2(KEYINPUT1), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G125), .ZN(new_n253));
  INV_X1    g067(.A(G146), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n250), .A2(new_n254), .A3(G143), .ZN(new_n255));
  INV_X1    g069(.A(G143), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n256), .B(G146), .C1(new_n250), .C2(KEYINPUT1), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n252), .A2(new_n253), .A3(new_n255), .A4(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n254), .A2(G143), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n256), .A2(G146), .ZN(new_n260));
  NAND2_X1  g074(.A1(KEYINPUT0), .A2(G128), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n261), .ZN(new_n263));
  NOR2_X1   g077(.A1(KEYINPUT0), .A2(G128), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n262), .B(G125), .C1(new_n265), .C2(new_n249), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n258), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G953), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G224), .ZN(new_n269));
  XOR2_X1   g083(.A(new_n267), .B(new_n269), .Z(new_n270));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n271), .B(new_n240), .C1(new_n246), .C2(new_n238), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n248), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT80), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n248), .A2(KEYINPUT80), .A3(new_n270), .A4(new_n272), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(G210), .B1(G237), .B2(G902), .ZN(new_n278));
  XOR2_X1   g092(.A(new_n278), .B(KEYINPUT85), .Z(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NOR3_X1   g094(.A1(new_n246), .A2(new_n238), .A3(new_n240), .ZN(new_n281));
  XNOR2_X1  g095(.A(KEYINPUT81), .B(KEYINPUT8), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n240), .B(new_n282), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n232), .A2(new_n233), .B1(new_n236), .B2(new_n194), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n283), .B1(new_n238), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n269), .A2(KEYINPUT7), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT82), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n266), .B1(new_n258), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT83), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n286), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n267), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n289), .B1(new_n286), .B2(KEYINPUT82), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n285), .A2(new_n290), .A3(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n291), .A2(KEYINPUT83), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n281), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(KEYINPUT84), .B1(new_n296), .B2(G902), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT84), .ZN(new_n298));
  INV_X1    g112(.A(G902), .ZN(new_n299));
  INV_X1    g113(.A(new_n295), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n242), .A2(new_n300), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n298), .B(new_n299), .C1(new_n301), .C2(new_n294), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n297), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n277), .A2(new_n280), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT87), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n277), .A2(new_n303), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n306), .A2(KEYINPUT86), .A3(new_n279), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT86), .ZN(new_n308));
  AOI22_X1  g122(.A1(new_n275), .A2(new_n276), .B1(new_n297), .B2(new_n302), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n308), .B1(new_n309), .B2(new_n280), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT87), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n309), .A2(new_n311), .A3(new_n280), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n305), .A2(new_n307), .A3(new_n310), .A4(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(G214), .B1(G237), .B2(G902), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT92), .ZN(new_n315));
  XNOR2_X1  g129(.A(G113), .B(G122), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(new_n207), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT91), .ZN(new_n318));
  INV_X1    g132(.A(G140), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G125), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n253), .A2(G140), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n318), .B1(new_n322), .B2(KEYINPUT19), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n322), .A2(KEYINPUT19), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT90), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n320), .A2(new_n321), .A3(KEYINPUT90), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n324), .B1(new_n328), .B2(KEYINPUT19), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n254), .B(new_n323), .C1(new_n329), .C2(new_n318), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n320), .A2(new_n321), .A3(new_n331), .A4(KEYINPUT16), .ZN(new_n332));
  AND3_X1   g146(.A1(new_n320), .A2(new_n321), .A3(KEYINPUT16), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT75), .B1(new_n320), .B2(KEYINPUT16), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G146), .ZN(new_n336));
  NOR2_X1   g150(.A1(G237), .A2(G953), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n337), .A2(KEYINPUT88), .A3(new_n256), .A4(G214), .ZN(new_n338));
  XOR2_X1   g152(.A(KEYINPUT88), .B(G143), .Z(new_n339));
  AND2_X1   g153(.A1(new_n337), .A2(G214), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n338), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G131), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI211_X1 g157(.A(G131), .B(new_n338), .C1(new_n339), .C2(new_n340), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n330), .A2(new_n336), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n328), .A2(G146), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n347), .B1(G146), .B2(new_n322), .ZN(new_n348));
  NAND2_X1  g162(.A1(KEYINPUT18), .A2(G131), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n350), .B(new_n338), .C1(new_n339), .C2(new_n340), .ZN(new_n351));
  OR2_X1    g165(.A1(new_n351), .A2(KEYINPUT89), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n341), .A2(new_n349), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n351), .A2(KEYINPUT89), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n348), .A2(new_n352), .A3(new_n353), .A4(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n317), .B1(new_n346), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT17), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n343), .A2(new_n357), .A3(new_n344), .ZN(new_n358));
  OR2_X1    g172(.A1(new_n344), .A2(new_n357), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n254), .B(new_n332), .C1(new_n333), .C2(new_n334), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n358), .A2(new_n359), .A3(new_n336), .A4(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n355), .A2(new_n361), .A3(new_n317), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n315), .B1(new_n356), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT20), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G475), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n367), .B(new_n299), .C1(new_n356), .C2(new_n363), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n346), .A2(new_n355), .ZN(new_n370));
  INV_X1    g184(.A(new_n317), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(G475), .B1(new_n372), .B2(new_n362), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n373), .A2(new_n365), .A3(new_n299), .A4(new_n364), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n369), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n317), .B1(new_n355), .B2(new_n361), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n299), .B1(new_n363), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G475), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n268), .A2(G952), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n380), .B1(G234), .B2(G237), .ZN(new_n381));
  XOR2_X1   g195(.A(KEYINPUT21), .B(G898), .Z(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(G234), .A2(G237), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(G902), .A3(G953), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n381), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G122), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G116), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n189), .A2(G122), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT93), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(G116), .B(G122), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT93), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G107), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n393), .A2(new_n395), .A3(new_n204), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(KEYINPUT94), .B1(new_n250), .B2(G143), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT94), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(new_n256), .A3(G128), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n250), .A2(G143), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G134), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n403), .A2(G134), .A3(new_n404), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT13), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n404), .A2(new_n409), .A3(G134), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n407), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n403), .A2(new_n409), .A3(G134), .A4(new_n404), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n399), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n189), .A2(KEYINPUT14), .A3(G122), .ZN(new_n414));
  OAI211_X1 g228(.A(G107), .B(new_n414), .C1(new_n391), .C2(KEYINPUT14), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n407), .A2(new_n398), .A3(new_n408), .A4(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  XOR2_X1   g231(.A(KEYINPUT9), .B(G234), .Z(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G217), .ZN(new_n420));
  NOR3_X1   g234(.A1(new_n419), .A2(new_n420), .A3(G953), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n417), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n413), .A2(new_n416), .A3(new_n421), .ZN(new_n424));
  AOI21_X1  g238(.A(G902), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT15), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(G478), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n425), .A2(KEYINPUT95), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n425), .A2(KEYINPUT95), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n427), .ZN(new_n431));
  INV_X1    g245(.A(new_n424), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n421), .B1(new_n413), .B2(new_n416), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n299), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT95), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n431), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n428), .B1(new_n430), .B2(new_n436), .ZN(new_n437));
  NOR3_X1   g251(.A1(new_n379), .A2(new_n387), .A3(new_n437), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n313), .A2(new_n314), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G469), .ZN(new_n440));
  NAND2_X1  g254(.A1(KEYINPUT11), .A2(G134), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  AND2_X1   g256(.A1(KEYINPUT65), .A2(G137), .ZN(new_n443));
  NOR2_X1   g257(.A1(KEYINPUT65), .A2(G137), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NOR2_X1   g259(.A1(KEYINPUT11), .A2(G134), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n446), .B1(G137), .B2(new_n441), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n445), .A2(new_n447), .A3(new_n342), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n342), .B1(new_n445), .B2(new_n447), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n252), .A2(new_n255), .A3(new_n257), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n452), .A2(new_n232), .A3(new_n233), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n452), .B1(new_n232), .B2(new_n233), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n451), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT12), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n455), .B(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n262), .B1(new_n265), .B2(new_n249), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n458), .B1(new_n219), .B2(new_n226), .ZN(new_n459));
  OR2_X1    g273(.A1(new_n453), .A2(KEYINPUT10), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n453), .A2(KEYINPUT10), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n459), .A2(new_n460), .A3(new_n450), .A4(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(G110), .B(G140), .ZN(new_n463));
  INV_X1    g277(.A(G227), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(G953), .ZN(new_n465));
  XOR2_X1   g279(.A(new_n463), .B(new_n465), .Z(new_n466));
  AND3_X1   g280(.A1(new_n457), .A2(new_n462), .A3(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n451), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n466), .B1(new_n469), .B2(new_n462), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n440), .B(new_n299), .C1(new_n467), .C2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(G469), .A2(G902), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n469), .A2(new_n462), .A3(new_n466), .ZN(new_n473));
  AND2_X1   g287(.A1(new_n457), .A2(new_n462), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n473), .B1(new_n474), .B2(new_n466), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n471), .B(new_n472), .C1(new_n440), .C2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(G221), .B1(new_n419), .B2(G902), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT32), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n458), .B1(new_n448), .B2(new_n449), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n443), .A2(new_n444), .A3(G134), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT66), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n483), .B1(new_n406), .B2(G137), .ZN(new_n484));
  INV_X1    g298(.A(G137), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n485), .A2(KEYINPUT66), .A3(G134), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(G131), .B1(new_n482), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n445), .A2(new_n447), .A3(new_n342), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n452), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n481), .A2(new_n490), .A3(new_n201), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(KEYINPUT68), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT68), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n481), .A2(new_n490), .A3(new_n201), .A4(new_n493), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT64), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n458), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n262), .B(KEYINPUT64), .C1(new_n265), .C2(new_n249), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n490), .B1(new_n499), .B2(new_n450), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT30), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n481), .A2(new_n490), .A3(KEYINPUT30), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(new_n202), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT31), .ZN(new_n505));
  XOR2_X1   g319(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n506));
  NAND2_X1  g320(.A1(new_n337), .A2(G210), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n506), .B(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT26), .B(G101), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n495), .A2(new_n504), .A3(new_n505), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(KEYINPUT70), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n495), .A2(new_n504), .A3(new_n510), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT31), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n491), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n516), .A2(KEYINPUT28), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n500), .A2(new_n202), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(new_n492), .A3(new_n494), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n517), .B1(new_n519), .B2(KEYINPUT28), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT71), .B1(new_n520), .B2(new_n510), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT71), .ZN(new_n522));
  INV_X1    g336(.A(new_n510), .ZN(new_n523));
  AND2_X1   g337(.A1(new_n519), .A2(KEYINPUT28), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n522), .B(new_n523), .C1(new_n524), .C2(new_n517), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n513), .A2(KEYINPUT70), .A3(KEYINPUT31), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n515), .A2(new_n521), .A3(new_n525), .A4(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(G472), .A2(G902), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n527), .A2(KEYINPUT72), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(KEYINPUT72), .B1(new_n527), .B2(new_n528), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n480), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n527), .A2(KEYINPUT32), .A3(new_n528), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n495), .A2(new_n504), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT73), .B1(new_n534), .B2(new_n510), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT29), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n520), .A2(new_n510), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT73), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n533), .A2(new_n538), .A3(new_n523), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n535), .A2(new_n536), .A3(new_n537), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n481), .A2(new_n490), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n202), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n492), .A2(new_n542), .A3(new_n494), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n517), .B1(new_n543), .B2(KEYINPUT28), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n523), .A2(new_n536), .ZN(new_n545));
  AOI21_X1  g359(.A(G902), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n540), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(G472), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n531), .A2(new_n532), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n336), .A2(new_n360), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT74), .B1(new_n187), .B2(G128), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(KEYINPUT23), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT23), .ZN(new_n553));
  OAI211_X1 g367(.A(KEYINPUT74), .B(new_n553), .C1(new_n187), .C2(G128), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n552), .B(new_n554), .C1(G119), .C2(new_n250), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(G110), .ZN(new_n556));
  XOR2_X1   g370(.A(G119), .B(G128), .Z(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT24), .B(G110), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n550), .B(new_n556), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n322), .A2(G146), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n560), .B1(new_n335), .B2(G146), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT76), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n557), .A2(new_n558), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n563), .B1(new_n555), .B2(G110), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n562), .B1(new_n561), .B2(new_n564), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n559), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(KEYINPUT77), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT77), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n559), .B(new_n569), .C1(new_n565), .C2(new_n566), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n268), .A2(G221), .A3(G234), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(KEYINPUT22), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(G137), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n567), .A2(new_n575), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n576), .A2(new_n299), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT25), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n420), .B1(G234), .B2(new_n299), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n574), .B1(new_n568), .B2(new_n570), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n582), .A2(new_n577), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT25), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(new_n584), .A3(new_n299), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n580), .A2(new_n581), .A3(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n581), .A2(G902), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n439), .A2(new_n479), .A3(new_n549), .A4(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(KEYINPUT96), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(G101), .ZN(G3));
  NAND2_X1  g406(.A1(new_n527), .A2(new_n299), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(G472), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n594), .B1(new_n529), .B2(new_n530), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n586), .A2(new_n588), .ZN(new_n596));
  NOR3_X1   g410(.A1(new_n595), .A2(new_n478), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT33), .B1(new_n432), .B2(new_n433), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT33), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n423), .A2(new_n599), .A3(new_n424), .ZN(new_n600));
  AOI21_X1  g414(.A(G902), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT98), .ZN(new_n602));
  XOR2_X1   g416(.A(KEYINPUT97), .B(G478), .Z(new_n603));
  OAI21_X1  g417(.A(new_n602), .B1(new_n425), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n603), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n434), .A2(KEYINPUT98), .A3(new_n605), .ZN(new_n606));
  AOI22_X1  g420(.A1(G478), .A2(new_n601), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n607), .B1(new_n375), .B2(new_n378), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n609), .A2(new_n387), .ZN(new_n610));
  INV_X1    g424(.A(new_n314), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n306), .A2(new_n279), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n611), .B1(new_n612), .B2(new_n304), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n597), .A2(new_n610), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(KEYINPUT34), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(new_n207), .ZN(G6));
  INV_X1    g430(.A(new_n387), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n277), .A2(new_n280), .A3(new_n303), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n280), .B1(new_n277), .B2(new_n303), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n314), .B(new_n437), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n373), .A2(KEYINPUT20), .A3(new_n299), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n368), .A2(new_n365), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n621), .A2(new_n378), .A3(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n597), .A2(new_n617), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(KEYINPUT35), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(new_n204), .ZN(G9));
  INV_X1    g441(.A(new_n595), .ZN(new_n628));
  OR2_X1    g442(.A1(new_n575), .A2(KEYINPUT36), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(KEYINPUT99), .ZN(new_n630));
  XOR2_X1   g444(.A(new_n630), .B(new_n571), .Z(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n587), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n586), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n633), .A2(new_n478), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n439), .A2(new_n628), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G110), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT100), .B(KEYINPUT37), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G12));
  INV_X1    g452(.A(new_n381), .ZN(new_n639));
  INV_X1    g453(.A(G900), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n386), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  OR2_X1    g457(.A1(new_n623), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n437), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n549), .A2(new_n613), .A3(new_n634), .A4(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G128), .ZN(G30));
  AND4_X1   g462(.A1(new_n305), .A2(new_n307), .A3(new_n310), .A4(new_n312), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(KEYINPUT38), .ZN(new_n650));
  XOR2_X1   g464(.A(new_n642), .B(KEYINPUT101), .Z(new_n651));
  XOR2_X1   g465(.A(new_n651), .B(KEYINPUT39), .Z(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n478), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n650), .B1(KEYINPUT40), .B2(new_n655), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n531), .A2(new_n532), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n534), .A2(new_n523), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n299), .B1(new_n543), .B2(new_n510), .ZN(new_n659));
  OAI21_X1  g473(.A(G472), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n437), .B1(new_n655), .B2(KEYINPUT40), .ZN(new_n662));
  AOI22_X1  g476(.A1(new_n369), .A2(new_n374), .B1(G475), .B2(new_n377), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n586), .A2(new_n632), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n656), .A2(new_n314), .A3(new_n661), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G143), .ZN(G45));
  AOI21_X1  g481(.A(KEYINPUT102), .B1(new_n608), .B2(new_n642), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT102), .ZN(new_n669));
  NOR4_X1   g483(.A1(new_n663), .A2(new_n669), .A3(new_n607), .A4(new_n643), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n549), .A2(new_n613), .A3(new_n671), .A4(new_n634), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G146), .ZN(G48));
  OAI21_X1  g487(.A(new_n314), .B1(new_n618), .B2(new_n619), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n299), .B1(new_n467), .B2(new_n470), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(G469), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n676), .A2(new_n477), .A3(new_n471), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n549), .A2(new_n589), .A3(new_n610), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT41), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G113), .ZN(G15));
  NOR2_X1   g495(.A1(new_n677), .A2(new_n387), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n549), .A2(new_n624), .A3(new_n589), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G116), .ZN(G18));
  NOR3_X1   g498(.A1(new_n674), .A2(new_n633), .A3(new_n677), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n549), .A3(new_n438), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G119), .ZN(G21));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n594), .A2(new_n688), .ZN(new_n689));
  OR2_X1    g503(.A1(new_n544), .A2(new_n510), .ZN(new_n690));
  AND2_X1   g504(.A1(new_n690), .A2(new_n514), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT103), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n511), .B1(new_n691), .B2(new_n692), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n528), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n593), .A2(KEYINPUT104), .A3(G472), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n689), .A2(new_n589), .A3(new_n695), .A4(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n682), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g513(.A(KEYINPUT105), .B1(new_n620), .B2(new_n663), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n613), .A2(new_n701), .A3(new_n437), .A4(new_n379), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G122), .ZN(G24));
  AND3_X1   g519(.A1(new_n689), .A2(new_n695), .A3(new_n696), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n706), .A2(new_n685), .A3(new_n671), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(KEYINPUT106), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(new_n253), .ZN(G27));
  NAND2_X1  g523(.A1(new_n532), .A2(KEYINPUT107), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n527), .A2(new_n528), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n480), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n527), .A2(new_n713), .A3(KEYINPUT32), .A4(new_n528), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n710), .A2(new_n712), .A3(new_n548), .A4(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT108), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n715), .A2(new_n716), .A3(new_n589), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n716), .B1(new_n715), .B2(new_n589), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n671), .A2(new_n649), .A3(new_n479), .A4(new_n314), .ZN(new_n720));
  OAI21_X1  g534(.A(KEYINPUT42), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT42), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n549), .A2(new_n722), .A3(new_n589), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n307), .A2(new_n310), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n305), .A2(new_n312), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n724), .A2(new_n725), .A3(new_n479), .A4(new_n314), .ZN(new_n726));
  OR2_X1    g540(.A1(new_n668), .A2(new_n670), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n723), .A2(new_n728), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n721), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G131), .ZN(G33));
  AND3_X1   g545(.A1(new_n549), .A2(new_n589), .A3(new_n646), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n313), .A2(new_n478), .A3(new_n611), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G134), .ZN(G36));
  NOR2_X1   g549(.A1(new_n313), .A2(new_n611), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n475), .B(KEYINPUT45), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(G469), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(KEYINPUT46), .A3(new_n472), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT46), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n740), .B(G469), .C1(new_n737), .C2(G902), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n739), .A2(new_n471), .A3(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n477), .A3(new_n652), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT44), .ZN(new_n744));
  INV_X1    g558(.A(new_n607), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n663), .A2(new_n745), .ZN(new_n746));
  XOR2_X1   g560(.A(new_n746), .B(KEYINPUT43), .Z(new_n747));
  NAND3_X1  g561(.A1(new_n747), .A2(new_n595), .A3(new_n664), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n743), .B1(new_n744), .B2(new_n748), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n748), .A2(new_n744), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n736), .B(new_n749), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G137), .ZN(G39));
  NAND2_X1  g569(.A1(new_n742), .A2(new_n477), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(KEYINPUT110), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT110), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n742), .A2(new_n758), .A3(new_n477), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT47), .ZN(new_n763));
  AOI22_X1  g577(.A1(new_n757), .A2(new_n759), .B1(KEYINPUT111), .B2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n736), .ZN(new_n765));
  NOR4_X1   g579(.A1(new_n762), .A2(new_n764), .A3(new_n727), .A4(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n549), .A2(new_n589), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G140), .ZN(G42));
  INV_X1    g583(.A(new_n746), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n676), .A2(new_n471), .ZN(new_n771));
  OAI211_X1 g585(.A(new_n770), .B(new_n314), .C1(KEYINPUT49), .C2(new_n771), .ZN(new_n772));
  AOI211_X1 g586(.A(new_n596), .B(new_n772), .C1(KEYINPUT49), .C2(new_n771), .ZN(new_n773));
  INV_X1    g587(.A(new_n661), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n773), .A2(new_n477), .A3(new_n774), .A4(new_n650), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n747), .A2(new_n381), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n776), .A2(new_n589), .A3(new_n706), .ZN(new_n777));
  INV_X1    g591(.A(new_n677), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(new_n613), .A3(new_n778), .ZN(new_n779));
  XOR2_X1   g593(.A(new_n779), .B(KEYINPUT121), .Z(new_n780));
  OAI22_X1  g594(.A1(new_n762), .A2(new_n764), .B1(new_n477), .B2(new_n771), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(new_n736), .A3(new_n777), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n736), .A2(new_n778), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n774), .A2(new_n784), .A3(new_n589), .A4(new_n381), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n785), .A2(new_n379), .A3(new_n745), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n782), .A2(new_n787), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n784), .A2(new_n776), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n593), .A2(KEYINPUT104), .A3(G472), .ZN(new_n790));
  AOI21_X1  g604(.A(KEYINPUT104), .B1(new_n593), .B2(G472), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n792), .A2(new_n664), .A3(new_n695), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n789), .A2(new_n793), .ZN(new_n794));
  XOR2_X1   g608(.A(new_n794), .B(KEYINPUT120), .Z(new_n795));
  NAND4_X1  g609(.A1(new_n777), .A2(new_n611), .A3(new_n650), .A4(new_n778), .ZN(new_n796));
  XOR2_X1   g610(.A(new_n796), .B(KEYINPUT50), .Z(new_n797));
  NAND3_X1  g611(.A1(new_n788), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT51), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n380), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n719), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n789), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(KEYINPUT48), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n785), .A2(new_n609), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n788), .A2(KEYINPUT51), .A3(new_n795), .A4(new_n797), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n800), .A2(new_n803), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n700), .A2(new_n702), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n792), .A2(new_n589), .A3(new_n682), .A4(new_n695), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n686), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n683), .A2(new_n679), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n597), .A2(new_n314), .A3(new_n313), .A4(new_n610), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n590), .A2(new_n635), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n437), .A2(KEYINPUT112), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT112), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n815), .B(new_n428), .C1(new_n430), .C2(new_n436), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n817), .A2(new_n379), .A3(new_n387), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n313), .A2(new_n314), .A3(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT113), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n313), .A2(KEYINPUT113), .A3(new_n818), .A4(new_n314), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n821), .A2(new_n597), .A3(new_n822), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n549), .A2(new_n634), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n644), .B1(new_n814), .B2(new_n816), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n824), .A2(new_n736), .A3(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n811), .A2(new_n813), .A3(new_n823), .A4(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n733), .A2(new_n664), .A3(new_n706), .A4(new_n671), .ZN(new_n828));
  AOI22_X1  g642(.A1(new_n828), .A2(KEYINPUT114), .B1(new_n732), .B2(new_n733), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT114), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n728), .A2(new_n830), .A3(new_n793), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n829), .A2(new_n721), .A3(new_n729), .A4(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(KEYINPUT115), .B1(new_n827), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n715), .A2(new_n716), .A3(new_n589), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n715), .A2(new_n589), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT108), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n720), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n729), .B(new_n831), .C1(new_n837), .C2(new_n722), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n828), .A2(KEYINPUT114), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n734), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n823), .A2(new_n590), .A3(new_n635), .A4(new_n812), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n704), .A2(new_n679), .A3(new_n683), .A4(new_n686), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n824), .A2(new_n736), .A3(new_n825), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT115), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n841), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n707), .A2(new_n647), .A3(new_n672), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT116), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n633), .A2(new_n849), .A3(new_n642), .ZN(new_n850));
  OAI21_X1  g664(.A(KEYINPUT116), .B1(new_n664), .B2(new_n643), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n478), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n661), .A2(new_n703), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT52), .B1(new_n848), .B2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n848), .A2(KEYINPUT52), .A3(new_n853), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n833), .A2(new_n847), .A3(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n858), .B(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(KEYINPUT54), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n858), .A2(new_n859), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT117), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n865));
  INV_X1    g679(.A(new_n856), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT53), .B1(new_n866), .B2(new_n854), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n841), .A2(new_n845), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT118), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n827), .A2(new_n832), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT118), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n870), .A2(new_n871), .A3(KEYINPUT53), .A4(new_n857), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n858), .A2(KEYINPUT117), .A3(new_n859), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n864), .A2(new_n865), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n861), .A2(new_n875), .A3(KEYINPUT119), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n858), .A2(KEYINPUT117), .A3(new_n859), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT117), .B1(new_n858), .B2(new_n859), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n869), .A2(new_n872), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT119), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n880), .A2(new_n881), .A3(new_n865), .ZN(new_n882));
  AOI211_X1 g696(.A(new_n780), .B(new_n806), .C1(new_n876), .C2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(G952), .A2(G953), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n775), .B1(new_n883), .B2(new_n884), .ZN(G75));
  NAND3_X1  g699(.A1(new_n864), .A2(new_n873), .A3(new_n874), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(G902), .A3(new_n279), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT56), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n248), .A2(new_n272), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(new_n270), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT55), .Z(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n887), .A2(new_n888), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n892), .B1(new_n887), .B2(new_n888), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n268), .A2(G952), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(G51));
  OR2_X1    g710(.A1(new_n467), .A2(new_n470), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n886), .A2(KEYINPUT54), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n875), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n472), .A2(KEYINPUT57), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n472), .A2(KEYINPUT57), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n897), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n880), .A2(new_n299), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n904), .A2(G469), .A3(new_n737), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n895), .B1(new_n903), .B2(new_n905), .ZN(G54));
  NAND3_X1  g720(.A1(new_n904), .A2(KEYINPUT58), .A3(G475), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n356), .A2(new_n363), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n895), .ZN(new_n910));
  INV_X1    g724(.A(new_n908), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n904), .A2(KEYINPUT58), .A3(G475), .A4(new_n911), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n909), .A2(new_n910), .A3(new_n912), .ZN(G60));
  NAND2_X1  g727(.A1(new_n598), .A2(new_n600), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n876), .A2(new_n882), .ZN(new_n916));
  NAND2_X1  g730(.A1(G478), .A2(G902), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT59), .Z(new_n918));
  OAI21_X1  g732(.A(new_n915), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n918), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n899), .A2(new_n914), .A3(new_n920), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n919), .A2(new_n910), .A3(new_n921), .ZN(G63));
  NAND2_X1  g736(.A1(G217), .A2(G902), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT60), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n886), .A2(new_n631), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n910), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n583), .B1(new_n886), .B2(new_n925), .ZN(new_n928));
  OAI211_X1 g742(.A(KEYINPUT122), .B(KEYINPUT61), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n583), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n931), .B1(new_n880), .B2(new_n924), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n932), .A2(new_n910), .A3(new_n926), .ZN(new_n933));
  AOI21_X1  g747(.A(KEYINPUT61), .B1(new_n933), .B2(KEYINPUT122), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n930), .A2(new_n934), .ZN(G66));
  INV_X1    g749(.A(G224), .ZN(new_n936));
  OAI21_X1  g750(.A(G953), .B1(new_n383), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n842), .A2(new_n843), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n937), .B1(new_n938), .B2(G953), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n889), .B1(G898), .B2(new_n268), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(G69));
  NAND2_X1  g755(.A1(new_n640), .A2(G953), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n502), .A2(new_n503), .ZN(new_n943));
  MUX2_X1   g757(.A(new_n324), .B(new_n329), .S(KEYINPUT91), .Z(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(KEYINPUT126), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n946), .A2(new_n464), .A3(G953), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n945), .A2(new_n942), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n549), .A2(new_n589), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n609), .B1(new_n379), .B2(new_n817), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n949), .A2(new_n654), .A3(new_n736), .A4(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n754), .A2(new_n951), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT124), .Z(new_n953));
  XOR2_X1   g767(.A(new_n848), .B(KEYINPUT123), .Z(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n666), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT62), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n953), .A2(new_n768), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n268), .ZN(new_n959));
  AOI22_X1  g773(.A1(new_n766), .A2(new_n767), .B1(new_n733), .B2(new_n732), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n801), .A2(new_n703), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n730), .B1(new_n743), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n960), .A2(new_n754), .A3(new_n954), .A4(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT125), .ZN(new_n965));
  OR2_X1    g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n964), .A2(new_n965), .ZN(new_n967));
  AOI21_X1  g781(.A(G953), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AOI22_X1  g782(.A1(new_n948), .A2(new_n959), .B1(new_n968), .B2(new_n945), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n942), .B(new_n947), .C1(new_n969), .C2(KEYINPUT126), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT126), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n947), .A2(new_n942), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n959), .A2(new_n948), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n968), .A2(new_n945), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n971), .B(new_n972), .C1(new_n973), .C2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n970), .A2(new_n975), .ZN(G72));
  NAND3_X1  g790(.A1(new_n966), .A2(new_n938), .A3(new_n967), .ZN(new_n977));
  NAND2_X1  g791(.A1(G472), .A2(G902), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT63), .Z(new_n979));
  AOI211_X1 g793(.A(new_n510), .B(new_n533), .C1(new_n977), .C2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n938), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n979), .B1(new_n958), .B2(new_n981), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n982), .A2(new_n658), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n535), .A2(new_n513), .A3(new_n539), .ZN(new_n984));
  AND3_X1   g798(.A1(new_n860), .A2(new_n979), .A3(new_n984), .ZN(new_n985));
  NOR4_X1   g799(.A1(new_n980), .A2(new_n983), .A3(new_n895), .A4(new_n985), .ZN(G57));
endmodule


