//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 0 0 0 0 0 1 0 1 0 0 1 0 0 1 0 1 0 1 1 1 1 1 1 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n208));
  NAND3_X1  g0008(.A1(new_n207), .A2(new_n208), .A3(KEYINPUT64), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n211));
  NAND3_X1  g0011(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  AOI21_X1  g0012(.A(KEYINPUT64), .B1(new_n207), .B2(new_n208), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n206), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT1), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n206), .A2(G13), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT0), .ZN(new_n218));
  INV_X1    g0018(.A(new_n201), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(new_n217), .A2(new_n218), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n225), .B1(new_n218), .B2(new_n217), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n215), .A2(new_n226), .ZN(G361));
  XOR2_X1   g0027(.A(G238), .B(G244), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT65), .B(KEYINPUT66), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n231), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(G97), .B(G107), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(KEYINPUT14), .ZN(new_n245));
  NOR2_X1   g0045(.A1(new_n245), .A2(KEYINPUT74), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT13), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT3), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G33), .ZN(new_n252));
  NAND4_X1  g0052(.A1(new_n250), .A2(new_n252), .A3(G232), .A4(G1698), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT71), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT3), .B(G33), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT71), .ZN(new_n256));
  NAND4_X1  g0056(.A1(new_n255), .A2(new_n256), .A3(G232), .A4(G1698), .ZN(new_n257));
  NAND2_X1  g0057(.A1(G33), .A2(G97), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n255), .A2(G226), .A3(new_n259), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n254), .A2(new_n257), .A3(new_n258), .A4(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n222), .B1(G33), .B2(G41), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT72), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n261), .A2(KEYINPUT72), .A3(new_n262), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G41), .ZN(new_n268));
  INV_X1    g0068(.A(G45), .ZN(new_n269));
  AOI21_X1  g0069(.A(G1), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G274), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n262), .A2(new_n270), .ZN(new_n273));
  OR2_X1    g0073(.A1(new_n273), .A2(KEYINPUT73), .ZN(new_n274));
  INV_X1    g0074(.A(G238), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n275), .B1(new_n273), .B2(KEYINPUT73), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n272), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n248), .B1(new_n267), .B2(new_n277), .ZN(new_n278));
  AND3_X1   g0078(.A1(new_n261), .A2(KEYINPUT72), .A3(new_n262), .ZN(new_n279));
  AOI21_X1  g0079(.A(KEYINPUT72), .B1(new_n261), .B2(new_n262), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n248), .B(new_n277), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  OAI211_X1 g0082(.A(G169), .B(new_n247), .C1(new_n278), .C2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n277), .B1(new_n279), .B2(new_n280), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT13), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(G179), .A3(new_n281), .ZN(new_n286));
  INV_X1    g0086(.A(G169), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n287), .B1(new_n285), .B2(new_n281), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT74), .B(KEYINPUT14), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n283), .B(new_n286), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G1), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(G13), .A3(G20), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G68), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT12), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(G20), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n223), .A2(G33), .ZN(new_n298));
  INV_X1    g0098(.A(G77), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n223), .A2(new_n249), .ZN(new_n300));
  OAI221_X1 g0100(.A(new_n297), .B1(new_n298), .B2(new_n299), .C1(new_n202), .C2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n222), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n301), .A2(KEYINPUT11), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n303), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n305), .B1(G1), .B2(new_n223), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n296), .B(new_n304), .C1(new_n294), .C2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(KEYINPUT11), .B1(new_n301), .B2(new_n303), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(G200), .B1(new_n278), .B2(new_n282), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n285), .A2(G190), .A3(new_n281), .ZN(new_n312));
  AND2_X1   g0112(.A1(new_n312), .A2(new_n309), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n290), .A2(new_n310), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n273), .ZN(new_n316));
  XNOR2_X1  g0116(.A(KEYINPUT67), .B(G226), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n271), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n250), .A2(new_n252), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n319), .A2(new_n259), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n320), .A2(G223), .B1(G77), .B2(new_n319), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n255), .A2(KEYINPUT68), .A3(G222), .A4(new_n259), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT68), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n255), .A2(new_n259), .ZN(new_n324));
  INV_X1    g0124(.A(G222), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n323), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n321), .A2(new_n322), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n318), .B1(new_n327), .B2(new_n262), .ZN(new_n328));
  INV_X1    g0128(.A(G200), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT70), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n330), .B(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n292), .A2(G50), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n303), .B1(new_n291), .B2(G20), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n333), .B1(new_n334), .B2(G50), .ZN(new_n335));
  XNOR2_X1  g0135(.A(KEYINPUT8), .B(G58), .ZN(new_n336));
  INV_X1    g0136(.A(G150), .ZN(new_n337));
  OAI22_X1  g0137(.A1(new_n336), .A2(new_n298), .B1(new_n337), .B2(new_n300), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n338), .B1(G20), .B2(new_n203), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n335), .B1(new_n339), .B2(new_n305), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT9), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n340), .B(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n342), .B1(G190), .B2(new_n328), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n332), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT10), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT10), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n332), .A2(new_n343), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G179), .ZN(new_n349));
  AND2_X1   g0149(.A1(new_n328), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n340), .B1(new_n328), .B2(G169), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT18), .ZN(new_n355));
  INV_X1    g0155(.A(new_n336), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n306), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n336), .A2(new_n292), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  XOR2_X1   g0159(.A(new_n359), .B(KEYINPUT78), .Z(new_n360));
  INV_X1    g0160(.A(KEYINPUT7), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(new_n255), .B2(G20), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n319), .A2(KEYINPUT7), .A3(new_n223), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(G68), .ZN(new_n365));
  INV_X1    g0165(.A(G58), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n366), .A2(new_n294), .ZN(new_n367));
  OAI21_X1  g0167(.A(G20), .B1(new_n367), .B2(new_n201), .ZN(new_n368));
  NOR2_X1   g0168(.A1(G20), .A2(G33), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n369), .A2(KEYINPUT75), .A3(G159), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(KEYINPUT75), .B1(new_n369), .B2(G159), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n368), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n365), .A2(KEYINPUT16), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT76), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n373), .B1(new_n364), .B2(G68), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT76), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(new_n378), .A3(KEYINPUT16), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n305), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  OAI211_X1 g0180(.A(KEYINPUT77), .B(new_n361), .C1(new_n255), .C2(G20), .ZN(new_n381));
  OAI211_X1 g0181(.A(G68), .B(new_n381), .C1(new_n364), .C2(KEYINPUT77), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n374), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT16), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n360), .B1(new_n380), .B2(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n250), .A2(new_n252), .A3(G223), .A4(new_n259), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT79), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT79), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n255), .A2(new_n389), .A3(G223), .A4(new_n259), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n255), .A2(G226), .A3(G1698), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G33), .A2(G87), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n388), .A2(new_n390), .A3(new_n391), .A4(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n262), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n272), .B1(new_n273), .B2(G232), .ZN(new_n395));
  AND3_X1   g0195(.A1(new_n394), .A2(G179), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n287), .B1(new_n394), .B2(new_n395), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n355), .B1(new_n386), .B2(new_n398), .ZN(new_n399));
  XNOR2_X1  g0199(.A(new_n359), .B(KEYINPUT78), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n378), .B1(new_n377), .B2(KEYINPUT16), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n294), .B1(new_n362), .B2(new_n363), .ZN(new_n402));
  NOR4_X1   g0202(.A1(new_n402), .A2(new_n373), .A3(KEYINPUT76), .A4(new_n384), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n303), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(KEYINPUT16), .B1(new_n382), .B2(new_n374), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n400), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OR2_X1    g0206(.A1(new_n396), .A2(new_n397), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n406), .A2(new_n407), .A3(KEYINPUT18), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n385), .B(new_n303), .C1(new_n403), .C2(new_n401), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n329), .B1(new_n394), .B2(new_n395), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n394), .A2(new_n395), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n410), .B1(new_n412), .B2(G190), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n409), .A2(new_n400), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT17), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT17), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n386), .A2(new_n416), .A3(new_n413), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n399), .A2(new_n408), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n272), .B1(new_n273), .B2(G244), .ZN(new_n420));
  INV_X1    g0220(.A(G107), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n319), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(G232), .A2(G1698), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n423), .B1(new_n275), .B2(G1698), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n422), .B(new_n262), .C1(new_n319), .C2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n420), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(G190), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g0228(.A(new_n428), .B(KEYINPUT69), .ZN(new_n429));
  OAI22_X1  g0229(.A1(new_n336), .A2(new_n300), .B1(new_n223), .B2(new_n299), .ZN(new_n430));
  XNOR2_X1  g0230(.A(KEYINPUT15), .B(G87), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n431), .A2(new_n298), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n303), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n334), .A2(G77), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n433), .B(new_n434), .C1(G77), .C2(new_n292), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n435), .B1(G200), .B2(new_n426), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n429), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n426), .A2(new_n287), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n420), .A2(new_n425), .A3(new_n349), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(new_n435), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  NOR4_X1   g0241(.A1(new_n315), .A2(new_n354), .A3(new_n419), .A4(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(KEYINPUT25), .B1(new_n293), .B2(new_n421), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n293), .A2(KEYINPUT25), .A3(new_n421), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n291), .A2(G33), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n292), .A2(new_n446), .A3(new_n222), .A4(new_n302), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n444), .A2(new_n445), .B1(new_n448), .B2(G107), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(G87), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(KEYINPUT85), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n255), .A2(new_n223), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT22), .ZN(new_n454));
  OR2_X1    g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n454), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G33), .A2(G116), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(G20), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT23), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n459), .B1(new_n223), .B2(G107), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n421), .A2(KEYINPUT23), .A3(G20), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n458), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n455), .A2(new_n456), .A3(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT24), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n305), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n455), .A2(KEYINPUT24), .A3(new_n456), .A4(new_n462), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n450), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  XNOR2_X1  g0267(.A(KEYINPUT5), .B(G41), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n269), .A2(G1), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n468), .A2(G274), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n262), .B1(new_n469), .B2(new_n468), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n471), .B1(new_n472), .B2(G264), .ZN(new_n473));
  NOR2_X1   g0273(.A1(G250), .A2(G1698), .ZN(new_n474));
  INV_X1    g0274(.A(G257), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n474), .B1(new_n475), .B2(G1698), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n255), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G294), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n479), .A2(KEYINPUT86), .A3(new_n262), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT86), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n476), .A2(new_n255), .B1(G33), .B2(G294), .ZN(new_n482));
  OAI211_X1 g0282(.A(G1), .B(G13), .C1(new_n249), .C2(new_n268), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n473), .A2(new_n480), .A3(new_n484), .A4(new_n427), .ZN(new_n485));
  AND2_X1   g0285(.A1(new_n472), .A2(G264), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n482), .A2(new_n483), .ZN(new_n487));
  NOR3_X1   g0287(.A1(new_n486), .A2(new_n487), .A3(new_n471), .ZN(new_n488));
  OAI22_X1  g0288(.A1(new_n485), .A2(KEYINPUT87), .B1(new_n488), .B2(G200), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n485), .A2(KEYINPUT87), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n467), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI211_X1 g0291(.A(G107), .B(new_n381), .C1(new_n364), .C2(KEYINPUT77), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n421), .A2(KEYINPUT6), .A3(G97), .ZN(new_n493));
  INV_X1    g0293(.A(new_n242), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n493), .B1(new_n494), .B2(KEYINPUT6), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n495), .A2(G20), .B1(G77), .B2(new_n369), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n305), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n447), .A2(G97), .ZN(new_n498));
  INV_X1    g0298(.A(G97), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n292), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g0301(.A(new_n501), .B(KEYINPUT80), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n250), .A2(new_n252), .A3(G244), .A4(new_n259), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT4), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n255), .A2(KEYINPUT4), .A3(G244), .A4(new_n259), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G283), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT81), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT81), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n510), .A2(G33), .A3(G283), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n255), .A2(G250), .A3(G1698), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n506), .A2(new_n507), .A3(new_n512), .A4(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n262), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n472), .A2(G257), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n515), .A2(new_n470), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G200), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n503), .B(new_n518), .C1(new_n427), .C2(new_n517), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n287), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n514), .A2(new_n262), .B1(G257), .B2(new_n472), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n521), .A2(new_n349), .A3(new_n470), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n520), .B(new_n522), .C1(new_n497), .C2(new_n502), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n491), .A2(new_n519), .A3(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT20), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n223), .B1(new_n499), .B2(G33), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n526), .B1(new_n509), .B2(new_n511), .ZN(new_n527));
  INV_X1    g0327(.A(G116), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n302), .A2(new_n222), .B1(G20), .B2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n525), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n509), .A2(new_n511), .ZN(new_n532));
  OAI211_X1 g0332(.A(KEYINPUT20), .B(new_n529), .C1(new_n532), .C2(new_n526), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n292), .A2(G116), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n535), .B1(new_n448), .B2(G116), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n468), .A2(new_n469), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n538), .A2(G270), .A3(new_n483), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT83), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n472), .A2(KEYINPUT83), .A3(G270), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n471), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(G303), .ZN(new_n544));
  OAI21_X1  g0344(.A(KEYINPUT84), .B1(new_n255), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n255), .A2(G264), .A3(G1698), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT84), .ZN(new_n548));
  OAI22_X1  g0348(.A1(new_n546), .A2(new_n548), .B1(new_n324), .B2(new_n475), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n262), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  AND4_X1   g0350(.A1(G179), .A2(new_n537), .A3(new_n543), .A4(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n543), .A2(new_n550), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n537), .B1(new_n553), .B2(G200), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n543), .A2(new_n550), .A3(G190), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n287), .B1(new_n534), .B2(new_n536), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n553), .A2(KEYINPUT21), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n553), .A2(new_n557), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT21), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AND4_X1   g0361(.A1(new_n552), .A2(new_n556), .A3(new_n558), .A4(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n473), .A2(new_n480), .A3(new_n484), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G169), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n488), .A2(G179), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n467), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n469), .A2(G274), .ZN(new_n567));
  OAI21_X1  g0367(.A(G250), .B1(new_n269), .B2(G1), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n567), .B1(new_n262), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n255), .A2(G238), .A3(new_n259), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n250), .A2(new_n252), .A3(G244), .A4(G1698), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n570), .A2(new_n457), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n569), .B1(new_n572), .B2(new_n262), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n349), .ZN(new_n574));
  INV_X1    g0374(.A(new_n431), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n575), .A2(new_n292), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n255), .A2(new_n223), .A3(G68), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT19), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n223), .B1(new_n258), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n451), .A2(new_n499), .A3(new_n421), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n578), .B1(new_n298), .B2(new_n499), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n577), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n576), .B1(new_n583), .B2(new_n303), .ZN(new_n584));
  XNOR2_X1  g0384(.A(new_n431), .B(KEYINPUT82), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n448), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n574), .B(new_n587), .C1(G169), .C2(new_n573), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n573), .A2(G190), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n447), .A2(new_n451), .ZN(new_n590));
  AOI211_X1 g0390(.A(new_n590), .B(new_n576), .C1(new_n583), .C2(new_n303), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n589), .B(new_n591), .C1(new_n329), .C2(new_n573), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n566), .A2(new_n593), .ZN(new_n594));
  AND4_X1   g0394(.A1(new_n442), .A2(new_n524), .A3(new_n562), .A4(new_n594), .ZN(G372));
  INV_X1    g0395(.A(KEYINPUT90), .ZN(new_n596));
  AOI211_X1 g0396(.A(new_n355), .B(new_n398), .C1(new_n409), .C2(new_n400), .ZN(new_n597));
  AOI21_X1  g0397(.A(KEYINPUT18), .B1(new_n406), .B2(new_n407), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n399), .A2(KEYINPUT90), .A3(new_n408), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n311), .A2(new_n309), .A3(new_n312), .ZN(new_n602));
  INV_X1    g0402(.A(new_n440), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n290), .A2(new_n310), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n604), .A2(KEYINPUT91), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n415), .A2(new_n417), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n604), .B2(KEYINPUT91), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n601), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n352), .B1(new_n608), .B2(new_n348), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n517), .A2(G179), .ZN(new_n610));
  AOI21_X1  g0410(.A(G169), .B1(new_n521), .B2(new_n470), .ZN(new_n611));
  NOR3_X1   g0411(.A1(new_n503), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT26), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n588), .A2(new_n592), .A3(KEYINPUT88), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT88), .B1(new_n588), .B2(new_n592), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n612), .B(new_n613), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(KEYINPUT26), .B1(new_n523), .B2(new_n593), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n616), .A2(new_n588), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(KEYINPUT89), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT89), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n616), .A2(new_n620), .A3(new_n588), .A4(new_n617), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n553), .A2(KEYINPUT21), .A3(new_n557), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT21), .B1(new_n553), .B2(new_n557), .ZN(new_n623));
  NOR3_X1   g0423(.A1(new_n622), .A2(new_n623), .A3(new_n551), .ZN(new_n624));
  INV_X1    g0424(.A(new_n467), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n565), .A2(new_n564), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT88), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n593), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n588), .A2(new_n592), .A3(KEYINPUT88), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n624), .A2(new_n627), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n524), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n619), .A2(new_n621), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n442), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n609), .A2(new_n634), .ZN(G369));
  INV_X1    g0435(.A(G13), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n636), .A2(G20), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n291), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(G213), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(G343), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n537), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n562), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(new_n624), .B2(new_n644), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n646), .A2(G330), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n625), .A2(KEYINPUT92), .A3(new_n643), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT92), .ZN(new_n649));
  INV_X1    g0449(.A(new_n643), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n649), .B1(new_n467), .B2(new_n650), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n648), .A2(new_n627), .A3(new_n651), .A4(new_n491), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n566), .A2(new_n643), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n647), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n552), .A2(new_n561), .A3(new_n558), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n650), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n652), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n627), .A2(new_n643), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n655), .A2(new_n660), .ZN(G399));
  INV_X1    g0461(.A(new_n216), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(G41), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n580), .A2(G116), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G1), .A3(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n220), .B2(new_n664), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT28), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT31), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n488), .A2(new_n521), .A3(new_n573), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n553), .A2(new_n349), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT30), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g0474(.A(new_n573), .B(KEYINPUT93), .Z(new_n675));
  NOR2_X1   g0475(.A1(new_n488), .A2(G179), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n675), .A2(new_n517), .A3(new_n553), .A4(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n670), .A2(new_n671), .A3(KEYINPUT30), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n674), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n669), .B1(new_n679), .B2(new_n643), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n524), .A2(new_n562), .A3(new_n594), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n680), .B1(new_n681), .B2(new_n643), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n679), .A2(new_n669), .A3(new_n643), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(G330), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT95), .ZN(new_n687));
  INV_X1    g0487(.A(new_n588), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n688), .B1(new_n631), .B2(new_n524), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n613), .B1(new_n523), .B2(new_n593), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT94), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OAI211_X1 g0492(.A(new_n612), .B(KEYINPUT26), .C1(new_n614), .C2(new_n615), .ZN(new_n693));
  OAI211_X1 g0493(.A(KEYINPUT94), .B(new_n613), .C1(new_n523), .C2(new_n593), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n689), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n687), .B1(new_n696), .B2(new_n650), .ZN(new_n697));
  AOI211_X1 g0497(.A(KEYINPUT95), .B(new_n643), .C1(new_n689), .C2(new_n695), .ZN(new_n698));
  OAI21_X1  g0498(.A(KEYINPUT29), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n633), .A2(new_n650), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT29), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n686), .B1(new_n699), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n668), .B1(new_n703), .B2(G1), .ZN(G364));
  AOI21_X1  g0504(.A(new_n291), .B1(new_n637), .B2(G45), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n663), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n647), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(G330), .B2(new_n646), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n662), .A2(new_n319), .ZN(new_n710));
  NAND2_X1  g0510(.A1(G355), .A2(KEYINPUT96), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(G355), .A2(KEYINPUT96), .ZN(new_n713));
  OAI22_X1  g0513(.A1(new_n712), .A2(new_n713), .B1(G116), .B2(new_n216), .ZN(new_n714));
  OR2_X1    g0514(.A1(new_n240), .A2(new_n269), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n662), .A2(new_n255), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n717), .B1(new_n269), .B2(new_n221), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n714), .B1(new_n715), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(G13), .A2(G33), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(G20), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n222), .B1(G20), .B2(new_n287), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n707), .B1(new_n719), .B2(new_n725), .ZN(new_n726));
  NOR4_X1   g0526(.A1(new_n223), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  OR2_X1    g0528(.A1(new_n728), .A2(KEYINPUT99), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(KEYINPUT99), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G159), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n223), .A2(new_n349), .A3(new_n329), .ZN(new_n734));
  OR2_X1    g0534(.A1(new_n734), .A2(KEYINPUT98), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(KEYINPUT98), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n735), .A2(new_n427), .A3(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AOI22_X1  g0538(.A1(new_n733), .A2(KEYINPUT32), .B1(G68), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n735), .A2(G190), .A3(new_n736), .ZN(new_n740));
  OAI221_X1 g0540(.A(new_n739), .B1(KEYINPUT32), .B2(new_n733), .C1(new_n202), .C2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n329), .A2(G179), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n742), .A2(G20), .A3(new_n427), .ZN(new_n743));
  OR2_X1    g0543(.A1(new_n743), .A2(KEYINPUT100), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(KEYINPUT100), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G107), .ZN(new_n748));
  OR3_X1    g0548(.A1(new_n223), .A2(new_n349), .A3(KEYINPUT97), .ZN(new_n749));
  OAI21_X1  g0549(.A(KEYINPUT97), .B1(new_n223), .B2(new_n349), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n427), .A2(G200), .ZN(new_n751));
  AND3_X1   g0551(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G58), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n742), .A2(G20), .A3(G190), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n255), .B1(new_n754), .B2(new_n451), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n427), .A2(G179), .A3(G200), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n223), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n755), .B1(G97), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G190), .A2(G200), .ZN(new_n760));
  AND3_X1   g0560(.A1(new_n749), .A2(new_n750), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G77), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n748), .A2(new_n753), .A3(new_n759), .A4(new_n762), .ZN(new_n763));
  AOI22_X1  g0563(.A1(new_n732), .A2(G329), .B1(G283), .B2(new_n747), .ZN(new_n764));
  INV_X1    g0564(.A(G322), .ZN(new_n765));
  INV_X1    g0565(.A(new_n752), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(G294), .ZN(new_n768));
  OAI221_X1 g0568(.A(new_n319), .B1(new_n754), .B2(new_n544), .C1(new_n757), .C2(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n769), .B1(G311), .B2(new_n761), .ZN(new_n770));
  INV_X1    g0570(.A(G326), .ZN(new_n771));
  XOR2_X1   g0571(.A(KEYINPUT33), .B(G317), .Z(new_n772));
  OAI221_X1 g0572(.A(new_n770), .B1(new_n771), .B2(new_n740), .C1(new_n737), .C2(new_n772), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n741), .A2(new_n763), .B1(new_n767), .B2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n726), .B1(new_n774), .B2(new_n723), .ZN(new_n775));
  INV_X1    g0575(.A(new_n722), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n775), .B1(new_n646), .B2(new_n776), .ZN(new_n777));
  AND2_X1   g0577(.A1(new_n709), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(G396));
  NAND2_X1  g0579(.A1(new_n435), .A2(new_n643), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n437), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(new_n440), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n603), .A2(new_n650), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n700), .B(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n686), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n707), .B1(new_n786), .B2(new_n686), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT103), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n790), .B1(new_n789), .B2(new_n788), .ZN(new_n791));
  INV_X1    g0591(.A(new_n754), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n319), .B1(new_n792), .B2(G50), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n793), .B1(new_n366), .B2(new_n757), .C1(new_n746), .C2(new_n294), .ZN(new_n794));
  AOI22_X1  g0594(.A1(G143), .A2(new_n752), .B1(new_n761), .B2(G159), .ZN(new_n795));
  INV_X1    g0595(.A(G137), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n795), .B1(new_n796), .B2(new_n740), .C1(new_n337), .C2(new_n737), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT34), .Z(new_n798));
  AOI211_X1 g0598(.A(new_n794), .B(new_n798), .C1(G132), .C2(new_n732), .ZN(new_n799));
  INV_X1    g0599(.A(G311), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n731), .A2(new_n800), .B1(new_n768), .B2(new_n766), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n319), .B1(new_n754), .B2(new_n421), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n746), .A2(new_n451), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n802), .B(new_n803), .C1(G97), .C2(new_n758), .ZN(new_n804));
  INV_X1    g0604(.A(G283), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n804), .B1(new_n805), .B2(new_n737), .C1(new_n544), .C2(new_n740), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n801), .B(new_n806), .C1(G116), .C2(new_n761), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n723), .B1(new_n799), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n723), .A2(new_n720), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT101), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n808), .B(new_n707), .C1(G77), .C2(new_n810), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n811), .A2(KEYINPUT102), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(KEYINPUT102), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n812), .B(new_n813), .C1(new_n721), .C2(new_n785), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n791), .A2(new_n814), .ZN(G384));
  OAI21_X1  g0615(.A(G77), .B1(new_n366), .B2(new_n294), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n220), .A2(new_n816), .B1(G50), .B2(new_n294), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n817), .A2(G1), .A3(new_n636), .ZN(new_n818));
  OAI211_X1 g0618(.A(G116), .B(new_n224), .C1(new_n495), .C2(KEYINPUT35), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(KEYINPUT35), .B2(new_n495), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n818), .B1(new_n820), .B2(KEYINPUT36), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(KEYINPUT36), .B2(new_n820), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n633), .A2(new_n650), .A3(new_n785), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n783), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n286), .B1(new_n288), .B2(new_n289), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n287), .B(new_n246), .C1(new_n285), .C2(new_n281), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n310), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(new_n650), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n310), .A2(new_n643), .ZN(new_n830));
  AOI21_X1  g0630(.A(KEYINPUT104), .B1(new_n314), .B2(new_n830), .ZN(new_n831));
  AND4_X1   g0631(.A1(KEYINPUT104), .A2(new_n827), .A3(new_n602), .A4(new_n830), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n829), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n824), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT38), .ZN(new_n835));
  INV_X1    g0635(.A(new_n641), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n303), .B1(new_n377), .B2(KEYINPUT16), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(new_n376), .B2(new_n379), .ZN(new_n838));
  INV_X1    g0638(.A(new_n359), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n407), .A2(new_n836), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n414), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(KEYINPUT37), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n406), .A2(new_n407), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n641), .B(KEYINPUT105), .Z(new_n844));
  NAND2_X1  g0644(.A1(new_n406), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT37), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n843), .A2(new_n845), .A3(new_n846), .A4(new_n414), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n842), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n836), .B1(new_n838), .B2(new_n839), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n399), .A2(new_n408), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n850), .B1(new_n851), .B2(new_n606), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n835), .B1(new_n849), .B2(new_n852), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n848), .B(KEYINPUT38), .C1(new_n418), .C2(new_n850), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n834), .A2(new_n856), .B1(new_n601), .B2(new_n844), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n827), .A2(new_n643), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n855), .A2(KEYINPUT39), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT39), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n599), .A2(new_n606), .A3(new_n600), .ZN(new_n862));
  INV_X1    g0662(.A(new_n845), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n843), .A2(new_n845), .A3(new_n414), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(KEYINPUT37), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n862), .A2(new_n863), .B1(new_n847), .B2(new_n865), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n861), .B(new_n854), .C1(new_n866), .C2(KEYINPUT38), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n859), .B1(new_n860), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n857), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n699), .A2(new_n442), .A3(new_n702), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n609), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n869), .B(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n682), .A2(new_n683), .A3(new_n785), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n833), .A2(new_n855), .A3(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT40), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n854), .B1(new_n866), .B2(KEYINPUT38), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n878), .A2(new_n833), .A3(KEYINPUT40), .A4(new_n874), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n877), .A2(G330), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n442), .A2(new_n686), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n862), .A2(new_n863), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n865), .A2(new_n847), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n835), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n876), .B1(new_n884), .B2(new_n854), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n827), .A2(new_n602), .A3(new_n830), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT104), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n314), .A2(KEYINPUT104), .A3(new_n830), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n828), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n890), .A2(new_n873), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n885), .A2(new_n891), .B1(new_n875), .B2(new_n876), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n442), .A2(new_n682), .A3(new_n683), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n880), .A2(new_n881), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n872), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(new_n291), .B2(new_n637), .ZN(new_n896));
  OAI22_X1  g0696(.A1(new_n896), .A2(KEYINPUT106), .B1(new_n872), .B2(new_n894), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n896), .A2(KEYINPUT106), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n822), .B1(new_n897), .B2(new_n898), .ZN(G367));
  INV_X1    g0699(.A(new_n723), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n747), .A2(G97), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n544), .B2(new_n766), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n255), .B1(new_n758), .B2(G107), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT112), .B1(new_n754), .B2(new_n528), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n903), .B1(KEYINPUT46), .B2(new_n904), .ZN(new_n905));
  OAI22_X1  g0705(.A1(new_n768), .A2(new_n737), .B1(new_n740), .B2(new_n800), .ZN(new_n906));
  NOR3_X1   g0706(.A1(new_n902), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(G317), .ZN(new_n908));
  INV_X1    g0708(.A(new_n761), .ZN(new_n909));
  OAI22_X1  g0709(.A1(new_n731), .A2(new_n908), .B1(new_n805), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(KEYINPUT46), .B2(new_n904), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n907), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n747), .A2(G77), .ZN(new_n913));
  OAI221_X1 g0713(.A(new_n913), .B1(new_n796), .B2(new_n731), .C1(new_n337), .C2(new_n766), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n757), .A2(new_n294), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n319), .B1(new_n792), .B2(G58), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n916), .B(new_n917), .C1(new_n909), .C2(new_n202), .ZN(new_n918));
  INV_X1    g0718(.A(new_n740), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n918), .B1(G143), .B2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(G159), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n920), .B1(new_n921), .B2(new_n737), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n912), .B1(new_n914), .B2(new_n922), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n923), .B(KEYINPUT113), .Z(new_n924));
  AOI21_X1  g0724(.A(new_n900), .B1(new_n924), .B2(KEYINPUT47), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(KEYINPUT47), .B2(new_n924), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n236), .A2(new_n716), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n725), .B1(new_n662), .B2(new_n575), .ZN(new_n928));
  AOI211_X1 g0728(.A(new_n663), .B(new_n706), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n650), .A2(new_n591), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n614), .B2(new_n615), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n930), .A2(new_n588), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n926), .B(new_n929), .C1(new_n776), .C2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n660), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n519), .B(new_n523), .C1(new_n503), .C2(new_n650), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n936), .A2(KEYINPUT108), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(KEYINPUT108), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n937), .A2(new_n938), .B1(new_n612), .B2(new_n643), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n935), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT44), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n940), .B(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n939), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n943), .A2(KEYINPUT45), .A3(new_n660), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT45), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n935), .B2(new_n939), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n942), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n655), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n942), .A2(new_n947), .A3(new_n655), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n652), .A2(new_n653), .A3(new_n657), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n953), .B(KEYINPUT110), .Z(new_n954));
  INV_X1    g0754(.A(new_n658), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n647), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n954), .A2(new_n647), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(KEYINPUT111), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT111), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n954), .A2(new_n959), .A3(new_n647), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n956), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n703), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n703), .B1(new_n952), .B2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n663), .B(KEYINPUT41), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n706), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n937), .A2(new_n938), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n523), .B1(new_n966), .B2(new_n627), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT109), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n643), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n968), .B2(new_n967), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n966), .A2(new_n955), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT42), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n933), .ZN(new_n974));
  XOR2_X1   g0774(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n655), .A2(new_n939), .ZN(new_n979));
  INV_X1    g0779(.A(new_n973), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT43), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n976), .B1(new_n981), .B2(new_n974), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n978), .B(new_n979), .C1(new_n980), .C2(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n980), .A2(new_n982), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n984), .A2(new_n977), .B1(new_n655), .B2(new_n939), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n934), .B1(new_n965), .B2(new_n986), .ZN(G387));
  OR3_X1    g0787(.A1(new_n961), .A2(new_n703), .A3(KEYINPUT116), .ZN(new_n988));
  OAI21_X1  g0788(.A(KEYINPUT116), .B1(new_n961), .B2(new_n703), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n988), .A2(new_n663), .A3(new_n962), .A4(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n654), .A2(new_n776), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n717), .B1(new_n231), .B2(G45), .ZN(new_n992));
  INV_X1    g0792(.A(new_n665), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n992), .B1(new_n993), .B2(new_n710), .ZN(new_n994));
  AOI21_X1  g0794(.A(G45), .B1(G68), .B2(G77), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n356), .A2(new_n202), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n665), .B(new_n995), .C1(new_n996), .C2(KEYINPUT50), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(KEYINPUT50), .B2(new_n996), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n994), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(new_n421), .B2(new_n662), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n707), .B1(new_n1000), .B2(new_n725), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n792), .A2(G77), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n901), .A2(new_n255), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(new_n356), .B2(new_n738), .ZN(new_n1004));
  AND2_X1   g0804(.A1(new_n585), .A2(new_n758), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(G50), .B2(new_n752), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n732), .A2(G150), .B1(G68), .B2(new_n761), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n919), .A2(G159), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1004), .A2(new_n1006), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n255), .B1(new_n747), .B2(G116), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n758), .A2(G283), .B1(new_n792), .B2(G294), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(G303), .A2(new_n761), .B1(new_n752), .B2(G317), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1012), .B1(new_n800), .B2(new_n737), .C1(new_n765), .C2(new_n740), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(KEYINPUT114), .B(KEYINPUT48), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1011), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT115), .Z(new_n1017));
  INV_X1    g0817(.A(KEYINPUT49), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1010), .B1(new_n771), .B2(new_n731), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1019));
  AND2_X1   g0819(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1009), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n991), .B(new_n1001), .C1(new_n1021), .C2(new_n723), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(new_n961), .B2(new_n706), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n990), .A2(new_n1023), .ZN(G393));
  NOR2_X1   g0824(.A1(new_n243), .A2(new_n717), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n724), .B1(new_n499), .B2(new_n216), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n707), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n761), .A2(new_n356), .B1(G77), .B2(new_n758), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n202), .B2(new_n737), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT117), .Z(new_n1030));
  AOI22_X1  g0830(.A1(new_n919), .A2(G150), .B1(new_n752), .B2(G159), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1030), .B1(KEYINPUT51), .B2(new_n1031), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n319), .B(new_n803), .C1(G68), .C2(new_n792), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1031), .A2(KEYINPUT51), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n732), .A2(G143), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n919), .A2(G317), .B1(new_n752), .B2(G311), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT52), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n732), .A2(G322), .B1(G294), .B2(new_n761), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n738), .A2(G303), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n319), .B1(new_n754), .B2(new_n805), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(G116), .B2(new_n758), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1039), .A2(new_n748), .A3(new_n1040), .A4(new_n1042), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n1032), .A2(new_n1036), .B1(new_n1038), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT118), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n900), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1027), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n943), .B2(new_n776), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n952), .B2(new_n705), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n663), .B1(new_n952), .B2(new_n962), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n952), .A2(new_n962), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1050), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(G390));
  NAND2_X1  g0855(.A1(new_n888), .A2(new_n889), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n1056), .A2(new_n829), .B1(new_n823), .B2(new_n783), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n860), .B(new_n867), .C1(new_n1057), .C2(new_n858), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n695), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n656), .A2(new_n566), .B1(new_n615), .B2(new_n614), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n491), .A2(new_n519), .A3(new_n523), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n588), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n650), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(KEYINPUT95), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n696), .A2(new_n687), .A3(new_n650), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1064), .A2(new_n1065), .A3(new_n783), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1066), .A2(new_n782), .A3(new_n833), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n858), .B1(new_n884), .B2(new_n854), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n833), .A2(G330), .A3(new_n874), .ZN(new_n1070));
  AND3_X1   g0870(.A1(new_n1058), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1070), .B1(new_n1058), .B2(new_n1069), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n891), .A2(G330), .B1(new_n1066), .B2(new_n782), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n682), .A2(G330), .A3(new_n683), .A4(new_n785), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1056), .A2(new_n829), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT119), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n890), .A2(KEYINPUT119), .A3(new_n1074), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1070), .A2(new_n1075), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n1073), .A2(new_n1079), .B1(new_n1080), .B2(new_n824), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n870), .A2(new_n609), .A3(new_n881), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n1071), .A2(new_n1072), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1070), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n858), .B1(new_n824), .B2(new_n833), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n860), .A2(new_n867), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1084), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1066), .A2(new_n782), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1091));
  AOI21_X1  g0891(.A(KEYINPUT119), .B1(new_n890), .B2(new_n1074), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1070), .B(new_n1090), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1080), .A2(new_n824), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1058), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1082), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1089), .A2(new_n1095), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1083), .A2(new_n1098), .A3(new_n663), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n707), .B1(new_n810), .B2(new_n356), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1087), .A2(new_n721), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n319), .B1(new_n754), .B2(new_n451), .C1(new_n757), .C2(new_n299), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n740), .A2(new_n805), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1102), .B(new_n1103), .C1(G68), .C2(new_n747), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n499), .A2(new_n909), .B1(new_n766), .B2(new_n528), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(G294), .B2(new_n732), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1104), .B(new_n1106), .C1(new_n421), .C2(new_n737), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n754), .A2(new_n337), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT53), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1109), .B(new_n255), .C1(new_n921), .C2(new_n757), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(G128), .B2(new_n919), .ZN(new_n1111));
  XOR2_X1   g0911(.A(KEYINPUT54), .B(G143), .Z(new_n1112));
  NAND2_X1  g0912(.A1(new_n761), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n737), .B2(new_n796), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT120), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n747), .A2(G50), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n732), .A2(G125), .B1(G132), .B2(new_n752), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1111), .A2(new_n1116), .A3(new_n1117), .A4(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1107), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1100), .B(new_n1101), .C1(new_n723), .C2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1122), .B1(new_n1123), .B2(new_n706), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1099), .A2(new_n1124), .ZN(G378));
  INV_X1    g0925(.A(new_n869), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n352), .B1(new_n345), .B2(new_n347), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n340), .A2(new_n836), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  OR3_X1    g0932(.A1(new_n1129), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1132), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(new_n892), .B2(G330), .ZN(new_n1136));
  AND4_X1   g0936(.A1(G330), .A2(new_n877), .A3(new_n879), .A4(new_n1135), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1126), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT122), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n892), .A2(G330), .A3(new_n1135), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1135), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n880), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1140), .A2(new_n1142), .A3(new_n869), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1138), .A2(new_n1139), .A3(new_n1143), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1140), .A2(new_n1142), .A3(KEYINPUT122), .A4(new_n869), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1098), .A2(new_n1097), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT57), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1148), .B1(new_n1098), .B2(new_n1097), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1138), .A2(new_n1143), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n664), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1144), .A2(new_n1145), .A3(new_n706), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n707), .B1(new_n810), .B2(G50), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n746), .A2(new_n366), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n585), .A2(new_n761), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1157), .B(new_n1158), .C1(new_n805), .C2(new_n731), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n740), .A2(new_n528), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n737), .A2(new_n499), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n752), .A2(G107), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n255), .A2(G41), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1162), .A2(new_n916), .A3(new_n1002), .A4(new_n1163), .ZN(new_n1164));
  NOR4_X1   g0964(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .A4(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(KEYINPUT58), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1163), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1167), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1168));
  AND2_X1   g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n758), .A2(G150), .B1(new_n792), .B2(new_n1112), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n909), .B2(new_n796), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(G125), .A2(new_n919), .B1(new_n738), .B2(G132), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1171), .B(new_n1173), .C1(G128), .C2(new_n752), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n747), .A2(G159), .ZN(new_n1177));
  AOI211_X1 g0977(.A(G33), .B(G41), .C1(new_n732), .C2(G124), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1169), .B1(KEYINPUT58), .B2(new_n1165), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1155), .B1(new_n1181), .B2(new_n723), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n1135), .B2(new_n721), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT121), .Z(new_n1184));
  NAND2_X1  g0984(.A1(new_n1154), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1153), .A2(new_n1186), .ZN(G375));
  NAND2_X1  g0987(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1188), .A2(new_n1189), .A3(new_n964), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n731), .A2(new_n544), .B1(new_n421), .B2(new_n909), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n1005), .B(new_n1191), .C1(G283), .C2(new_n752), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n255), .B1(new_n792), .B2(G97), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n913), .B(new_n1193), .C1(new_n768), .C2(new_n740), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G116), .B2(new_n738), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n732), .A2(G128), .B1(G137), .B2(new_n752), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n319), .B1(new_n792), .B2(G159), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(G132), .A2(new_n919), .B1(new_n738), .B2(new_n1112), .ZN(new_n1198));
  AND4_X1   g0998(.A1(new_n1157), .A2(new_n1196), .A3(new_n1197), .A4(new_n1198), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n761), .A2(G150), .B1(G50), .B2(new_n758), .ZN(new_n1200));
  XOR2_X1   g1000(.A(new_n1200), .B(KEYINPUT124), .Z(new_n1201));
  AOI22_X1  g1001(.A1(new_n1192), .A2(new_n1195), .B1(new_n1199), .B2(new_n1201), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n707), .B1(G68), .B2(new_n810), .C1(new_n1202), .C2(new_n900), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n890), .B2(new_n720), .ZN(new_n1204));
  XOR2_X1   g1004(.A(new_n705), .B(KEYINPUT123), .Z(new_n1205));
  AOI21_X1  g1005(.A(new_n1204), .B1(new_n1095), .B2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1190), .A2(new_n1206), .ZN(G381));
  AOI21_X1  g1007(.A(new_n1185), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1208));
  INV_X1    g1008(.A(G378), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n1054), .B(new_n934), .C1(new_n965), .C2(new_n986), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(G393), .A2(G396), .ZN(new_n1212));
  INV_X1    g1012(.A(G384), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  OR4_X1    g1014(.A1(G381), .A2(new_n1210), .A3(new_n1211), .A4(new_n1214), .ZN(G407));
  OAI211_X1 g1015(.A(G407), .B(G213), .C1(G343), .C2(new_n1210), .ZN(G409));
  NAND2_X1  g1016(.A1(G390), .A2(G387), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n778), .B1(new_n990), .B2(new_n1023), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1212), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT126), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n1217), .A2(new_n1211), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n1217), .A2(new_n1211), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1223));
  OAI21_X1  g1023(.A(KEYINPUT126), .B1(new_n1212), .B2(new_n1218), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1221), .B1(new_n1222), .B2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1209), .B1(new_n1153), .B2(new_n1186), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT60), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1189), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1081), .A2(KEYINPUT60), .A3(new_n1082), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1229), .A2(new_n663), .A3(new_n1188), .A4(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1231), .A2(G384), .A3(new_n1206), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(G384), .B1(new_n1231), .B2(new_n1206), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(G213), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1237), .A2(G343), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1144), .A2(new_n1146), .A3(new_n964), .A4(new_n1145), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1151), .A2(new_n1205), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1242), .A2(new_n1099), .A3(new_n1124), .A4(new_n1184), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1239), .B1(new_n1241), .B2(new_n1243), .ZN(new_n1244));
  NOR3_X1   g1044(.A1(new_n1227), .A2(new_n1236), .A3(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1226), .B1(new_n1245), .B2(KEYINPUT63), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1099), .A2(new_n1124), .A3(new_n1184), .ZN(new_n1247));
  AND2_X1   g1047(.A1(new_n1151), .A2(new_n1205), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1238), .B1(new_n1249), .B2(new_n1240), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1250), .B(new_n1235), .C1(new_n1208), .C2(new_n1209), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT63), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT125), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  OAI211_X1 g1055(.A(G2897), .B(new_n1238), .C1(new_n1233), .C2(new_n1234), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1234), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1238), .A2(G2897), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1257), .A2(new_n1232), .A3(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1256), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1250), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1262));
  AOI21_X1  g1062(.A(KEYINPUT61), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1251), .A2(KEYINPUT125), .A3(new_n1252), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1246), .A2(new_n1255), .A3(new_n1263), .A4(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT127), .ZN(new_n1266));
  AND3_X1   g1066(.A1(new_n1251), .A2(new_n1266), .A3(KEYINPUT62), .ZN(new_n1267));
  AOI21_X1  g1067(.A(KEYINPUT62), .B1(new_n1251), .B2(new_n1266), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT61), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1244), .B1(G375), .B2(G378), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1269), .B1(new_n1270), .B2(new_n1260), .ZN(new_n1271));
  NOR3_X1   g1071(.A1(new_n1267), .A2(new_n1268), .A3(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1226), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1265), .B1(new_n1272), .B2(new_n1273), .ZN(G405));
  NAND2_X1  g1074(.A1(G375), .A2(G378), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1210), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1235), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1275), .A2(new_n1210), .A3(new_n1236), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1279), .B(new_n1273), .ZN(G402));
endmodule


