//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 0 1 0 0 1 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 1 0 1 1 0 0 0 1 0 1 0 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0 1 1 1 0 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n446, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n546, new_n547, new_n548, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n615, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT66), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT67), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT68), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT69), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT70), .Z(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT71), .Z(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n456), .A2(G567), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n459), .A2(KEYINPUT72), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(KEYINPUT72), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n454), .A2(G2106), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  OR2_X1    g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n467), .A2(G137), .B1(G101), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n471), .B1(new_n465), .B2(new_n466), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(KEYINPUT73), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT73), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(G113), .A3(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g052(.A(G2105), .B1(new_n472), .B2(new_n477), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n470), .A2(new_n478), .ZN(G160));
  XNOR2_X1  g054(.A(KEYINPUT3), .B(G2104), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  OAI21_X1  g056(.A(KEYINPUT74), .B1(new_n481), .B2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT74), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n467), .A2(new_n483), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n468), .B1(new_n465), .B2(new_n466), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  XOR2_X1   g063(.A(new_n488), .B(KEYINPUT75), .Z(new_n489));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n491));
  AND3_X1   g066(.A1(new_n486), .A2(new_n489), .A3(new_n491), .ZN(G162));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(G2105), .B1(KEYINPUT76), .B2(G114), .ZN(new_n494));
  AND2_X1   g069(.A1(KEYINPUT76), .A2(G114), .ZN(new_n495));
  OAI211_X1 g070(.A(G2104), .B(new_n493), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  AND2_X1   g071(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n497));
  NOR2_X1   g072(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n498));
  OAI211_X1 g073(.A(G126), .B(G2105), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(G138), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(G2105), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n502), .B1(new_n497), .B2(new_n498), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT4), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n502), .B(new_n505), .C1(new_n498), .C2(new_n497), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n500), .B1(new_n504), .B2(new_n506), .ZN(G164));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT5), .B(G543), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(new_n513), .A3(G88), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n515), .B1(new_n510), .B2(new_n511), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G50), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  OAI211_X1 g093(.A(new_n514), .B(new_n517), .C1(new_n518), .C2(new_n509), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n512), .A2(new_n513), .ZN(new_n523));
  XOR2_X1   g098(.A(KEYINPUT77), .B(G89), .Z(new_n524));
  OAI21_X1  g099(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT78), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(G63), .A2(G651), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n516), .A2(G51), .B1(new_n513), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n529), .B1(new_n525), .B2(new_n526), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n527), .A2(new_n530), .ZN(G168));
  XNOR2_X1  g106(.A(KEYINPUT79), .B(G52), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n516), .A2(new_n532), .ZN(new_n533));
  XOR2_X1   g108(.A(KEYINPUT80), .B(G90), .Z(new_n534));
  AOI22_X1  g109(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  OAI221_X1 g110(.A(new_n533), .B1(new_n523), .B2(new_n534), .C1(new_n535), .C2(new_n509), .ZN(G301));
  INV_X1    g111(.A(G301), .ZN(G171));
  NAND2_X1  g112(.A1(new_n516), .A2(G43), .ZN(new_n538));
  INV_X1    g113(.A(G81), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n539), .B2(new_n523), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n509), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND4_X1  g122(.A1(G319), .A2(G483), .A3(G661), .A4(new_n547), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT81), .ZN(G188));
  NAND2_X1  g124(.A1(new_n512), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G53), .ZN(new_n551));
  OAI21_X1  g126(.A(KEYINPUT9), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT9), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n516), .A2(new_n553), .A3(G53), .ZN(new_n554));
  AND2_X1   g129(.A1(new_n512), .A2(new_n513), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n552), .A2(new_n554), .B1(G91), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(G78), .A2(G543), .ZN(new_n557));
  AND2_X1   g132(.A1(KEYINPUT5), .A2(G543), .ZN(new_n558));
  NOR2_X1   g133(.A1(KEYINPUT5), .A2(G543), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n557), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT82), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI211_X1 g139(.A(KEYINPUT82), .B(new_n557), .C1(new_n560), .C2(new_n561), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n564), .A2(G651), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n556), .A2(new_n566), .ZN(G299));
  INV_X1    g142(.A(G168), .ZN(G286));
  INV_X1    g143(.A(G74), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n509), .B1(new_n560), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n570), .B1(G87), .B2(new_n555), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n516), .A2(KEYINPUT83), .A3(G49), .ZN(new_n572));
  INV_X1    g147(.A(new_n511), .ZN(new_n573));
  NOR2_X1   g148(.A1(KEYINPUT6), .A2(G651), .ZN(new_n574));
  OAI211_X1 g149(.A(G49), .B(G543), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT83), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n572), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n571), .A2(new_n578), .ZN(G288));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G61), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n560), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(G651), .B1(G48), .B2(new_n516), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n512), .A2(new_n513), .A3(G86), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n584), .A2(KEYINPUT84), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(KEYINPUT84), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n583), .A2(new_n585), .A3(new_n586), .ZN(G305));
  NAND2_X1  g162(.A1(new_n516), .A2(G47), .ZN(new_n588));
  INV_X1    g163(.A(G85), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n589), .B2(new_n523), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n591), .A2(new_n509), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  INV_X1    g170(.A(G54), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT86), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n596), .B1(new_n550), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n598), .B1(new_n597), .B2(new_n550), .ZN(new_n599));
  XNOR2_X1  g174(.A(KEYINPUT85), .B(KEYINPUT10), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n555), .A2(G92), .A3(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n600), .ZN(new_n602));
  INV_X1    g177(.A(G92), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n523), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n513), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n606), .A2(new_n509), .ZN(new_n607));
  AND3_X1   g182(.A1(new_n599), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n595), .B1(new_n608), .B2(G868), .ZN(G284));
  OAI21_X1  g184(.A(new_n595), .B1(new_n608), .B2(G868), .ZN(G321));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(G299), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(new_n611), .B2(G168), .ZN(G297));
  OAI21_X1  g188(.A(new_n612), .B1(new_n611), .B2(G168), .ZN(G280));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n608), .B1(new_n615), .B2(G860), .ZN(G148));
  NAND2_X1  g191(.A1(new_n608), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G868), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(G868), .B2(new_n543), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g195(.A1(new_n485), .A2(G135), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  INV_X1    g197(.A(G111), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G2105), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n624), .B1(G123), .B2(new_n487), .ZN(new_n625));
  AND2_X1   g200(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n480), .A2(new_n469), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  AOI22_X1  g206(.A1(G2096), .A2(new_n627), .B1(new_n631), .B2(G2100), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(G2100), .ZN(new_n633));
  OAI211_X1 g208(.A(new_n632), .B(new_n633), .C1(G2096), .C2(new_n627), .ZN(G156));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2435), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT88), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2427), .B(G2430), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(KEYINPUT14), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT89), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT87), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n642), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(G14), .A3(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(G401));
  XNOR2_X1  g228(.A(G2084), .B(G2090), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2072), .B(G2078), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT90), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n654), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(KEYINPUT91), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n656), .B(KEYINPUT17), .Z(new_n662));
  INV_X1    g237(.A(new_n657), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n660), .B(new_n661), .C1(new_n662), .C2(new_n663), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n654), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n656), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT18), .Z(new_n667));
  NOR2_X1   g242(.A1(new_n654), .A2(new_n657), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n664), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G2096), .B(G2100), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G227));
  XNOR2_X1  g247(.A(G1956), .B(G2474), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1961), .B(G1966), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n675), .A2(KEYINPUT92), .ZN(new_n676));
  XOR2_X1   g251(.A(G1971), .B(G1976), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(KEYINPUT92), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n676), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT20), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n673), .A2(new_n674), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(new_n678), .B2(new_n675), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT93), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n678), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n683), .B(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n681), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT94), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n687), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1991), .B(G1996), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1981), .B(G1986), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(G229));
  INV_X1    g269(.A(KEYINPUT95), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n695), .A2(G29), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(G29), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n626), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT31), .B(G11), .Z(new_n701));
  INV_X1    g276(.A(G28), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n702), .A2(KEYINPUT30), .ZN(new_n703));
  AOI21_X1  g278(.A(G29), .B1(new_n702), .B2(KEYINPUT30), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n701), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n700), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(G5), .A2(G16), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT101), .Z(new_n708));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(G301), .B2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G1961), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(G160), .A2(G29), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT24), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n714), .A2(G34), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(G34), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n698), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G2084), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR3_X1   g295(.A1(new_n706), .A2(new_n712), .A3(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(G4), .A2(G16), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT99), .Z(new_n723));
  INV_X1    g298(.A(new_n608), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(new_n709), .ZN(new_n725));
  INV_X1    g300(.A(G1348), .ZN(new_n726));
  INV_X1    g301(.A(G1956), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n709), .A2(G20), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT23), .Z(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G299), .B2(G16), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n725), .A2(new_n726), .B1(new_n727), .B2(new_n730), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n721), .B(new_n731), .C1(new_n727), .C2(new_n730), .ZN(new_n732));
  NOR2_X1   g307(.A1(G16), .A2(G19), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n543), .B2(G16), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(G1341), .Z(new_n735));
  INV_X1    g310(.A(G32), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n736), .A2(G29), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n469), .A2(G105), .ZN(new_n738));
  NAND3_X1  g313(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT26), .ZN(new_n740));
  AOI211_X1 g315(.A(new_n738), .B(new_n740), .C1(G129), .C2(new_n487), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n482), .A2(new_n484), .ZN(new_n742));
  INV_X1    g317(.A(G141), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n737), .B1(new_n744), .B2(G29), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT27), .B(G1996), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n699), .A2(G27), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G164), .B2(new_n699), .ZN(new_n749));
  INV_X1    g324(.A(G2078), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n735), .A2(new_n747), .A3(new_n751), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n732), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT25), .Z(new_n755));
  AOI22_X1  g330(.A1(new_n480), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n755), .B1(new_n756), .B2(new_n468), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n485), .B2(G139), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT100), .ZN(new_n759));
  MUX2_X1   g334(.A(G33), .B(new_n759), .S(G29), .Z(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G2072), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n725), .A2(new_n726), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n709), .A2(G21), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G168), .B2(new_n709), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n762), .B1(new_n764), .B2(G1966), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n698), .A2(G26), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT28), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n485), .A2(G140), .ZN(new_n768));
  OAI21_X1  g343(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n769));
  INV_X1    g344(.A(G116), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n769), .B1(new_n770), .B2(G2105), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G128), .B2(new_n487), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n767), .B1(new_n773), .B2(G29), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G2067), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n765), .B(new_n775), .C1(G1966), .C2(new_n764), .ZN(new_n776));
  NOR3_X1   g351(.A1(new_n753), .A2(new_n761), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(G162), .A2(new_n699), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G35), .B2(new_n699), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n779), .A2(KEYINPUT29), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(KEYINPUT29), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(G2090), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n780), .A2(G2090), .A3(new_n781), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n718), .A2(new_n719), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n710), .A2(new_n711), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n786), .B(new_n787), .C1(new_n745), .C2(new_n746), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT102), .Z(new_n789));
  NAND3_X1  g364(.A1(new_n784), .A2(new_n785), .A3(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n777), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n709), .A2(G23), .ZN(new_n793));
  INV_X1    g368(.A(G288), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(new_n709), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT33), .ZN(new_n796));
  INV_X1    g371(.A(G1976), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  MUX2_X1   g373(.A(G6), .B(G305), .S(G16), .Z(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT32), .B(G1981), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  NOR2_X1   g377(.A1(G16), .A2(G22), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G166), .B2(G16), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT97), .B(G1971), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n801), .A2(new_n802), .A3(new_n806), .ZN(new_n807));
  OR3_X1    g382(.A1(new_n798), .A2(KEYINPUT34), .A3(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(KEYINPUT34), .B1(new_n798), .B2(new_n807), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n485), .A2(G131), .ZN(new_n810));
  OAI21_X1  g385(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n811));
  INV_X1    g386(.A(G107), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n811), .B1(new_n812), .B2(G2105), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(G119), .B2(new_n487), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n816), .A2(new_n698), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(G25), .B2(new_n698), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT35), .B(G1991), .Z(new_n819));
  AND2_X1   g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n818), .A2(new_n819), .ZN(new_n821));
  INV_X1    g396(.A(G24), .ZN(new_n822));
  OR3_X1    g397(.A1(new_n822), .A2(KEYINPUT96), .A3(G16), .ZN(new_n823));
  OAI21_X1  g398(.A(KEYINPUT96), .B1(new_n822), .B2(G16), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n823), .B(new_n824), .C1(new_n593), .C2(new_n709), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G1986), .ZN(new_n826));
  NOR3_X1   g401(.A1(new_n820), .A2(new_n821), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n808), .A2(new_n809), .A3(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT98), .B(KEYINPUT36), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n808), .A2(new_n809), .A3(new_n827), .A4(new_n829), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n792), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT103), .ZN(G311));
  INV_X1    g409(.A(new_n833), .ZN(G150));
  NAND2_X1  g410(.A1(new_n608), .A2(G559), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT38), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n516), .A2(G55), .ZN(new_n838));
  INV_X1    g413(.A(G93), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n838), .B1(new_n839), .B2(new_n523), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n841), .A2(new_n509), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n543), .A2(new_n843), .ZN(new_n844));
  OAI22_X1  g419(.A1(new_n542), .A2(new_n540), .B1(new_n840), .B2(new_n842), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n837), .B(new_n847), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n848), .A2(KEYINPUT39), .ZN(new_n849));
  INV_X1    g424(.A(G860), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(KEYINPUT39), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n843), .A2(new_n850), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT37), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n854), .ZN(G145));
  XOR2_X1   g430(.A(G160), .B(KEYINPUT104), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n627), .B(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(G162), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n773), .B(new_n744), .Z(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(G164), .Z(new_n861));
  INV_X1    g436(.A(new_n759), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n487), .A2(G130), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n468), .A2(G118), .ZN(new_n865));
  OAI21_X1  g440(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n867), .B1(new_n485), .B2(G142), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(new_n629), .Z(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n816), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n860), .B(G164), .ZN(new_n871));
  INV_X1    g446(.A(new_n758), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AND3_X1   g448(.A1(new_n863), .A2(new_n870), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n870), .B1(new_n863), .B2(new_n873), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n859), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n863), .A2(new_n873), .ZN(new_n877));
  INV_X1    g452(.A(new_n870), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n863), .A2(new_n870), .A3(new_n873), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(new_n858), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(G37), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n876), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g459(.A(new_n611), .B1(new_n840), .B2(new_n842), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n847), .B(new_n617), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT105), .ZN(new_n887));
  NAND2_X1  g462(.A1(G299), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n556), .A2(new_n566), .A3(KEYINPUT105), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n608), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n888), .A2(new_n608), .A3(new_n890), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n886), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT41), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n892), .A2(KEYINPUT41), .A3(new_n893), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n896), .B1(new_n886), .B2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n794), .B(G305), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n593), .B(G303), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n902), .B(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT42), .ZN(new_n905));
  OR3_X1    g480(.A1(new_n901), .A2(new_n905), .A3(KEYINPUT106), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n901), .B1(new_n905), .B2(KEYINPUT106), .ZN(new_n907));
  AOI22_X1  g482(.A1(new_n906), .A2(new_n907), .B1(KEYINPUT106), .B2(new_n905), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n885), .B1(new_n908), .B2(new_n611), .ZN(G295));
  OAI21_X1  g484(.A(new_n885), .B1(new_n908), .B2(new_n611), .ZN(G331));
  INV_X1    g485(.A(KEYINPUT109), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT107), .ZN(new_n913));
  OAI21_X1  g488(.A(G301), .B1(new_n527), .B2(new_n530), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NOR3_X1   g490(.A1(new_n527), .A2(new_n530), .A3(G301), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n846), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(G168), .A2(G171), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n918), .A2(new_n845), .A3(new_n844), .A4(new_n914), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n913), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n919), .A2(new_n913), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n898), .B(new_n899), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n917), .A2(new_n919), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n895), .A2(new_n923), .A3(KEYINPUT108), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n917), .A2(new_n919), .A3(new_n892), .A4(new_n893), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT108), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n922), .A2(new_n904), .A3(new_n924), .A4(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n882), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n925), .B(KEYINPUT108), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n904), .B1(new_n930), .B2(new_n922), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n912), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n904), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n900), .A2(new_n923), .ZN(new_n935));
  NOR3_X1   g510(.A1(new_n920), .A2(new_n921), .A3(new_n894), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AND4_X1   g512(.A1(KEYINPUT43), .A2(new_n937), .A3(new_n882), .A4(new_n928), .ZN(new_n938));
  OAI21_X1  g513(.A(KEYINPUT44), .B1(new_n933), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n928), .A2(new_n882), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n930), .A2(new_n922), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n934), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n912), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n937), .A2(new_n912), .A3(new_n882), .A4(new_n928), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n940), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n911), .B1(new_n939), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n941), .A2(KEYINPUT43), .A3(new_n937), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n940), .B1(new_n949), .B2(new_n932), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT43), .B1(new_n929), .B2(new_n931), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT44), .B1(new_n951), .B2(new_n945), .ZN(new_n952));
  NOR3_X1   g527(.A1(new_n950), .A2(new_n952), .A3(KEYINPUT109), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n948), .A2(new_n953), .ZN(G397));
  NAND2_X1  g529(.A1(new_n773), .A2(G2067), .ZN(new_n955));
  INV_X1    g530(.A(G2067), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n768), .A2(new_n956), .A3(new_n772), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(G1996), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n744), .B(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  XOR2_X1   g536(.A(new_n815), .B(new_n819), .Z(new_n962));
  NOR2_X1   g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n593), .B(G1986), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G1384), .ZN(new_n966));
  INV_X1    g541(.A(new_n506), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n505), .B1(new_n480), .B2(new_n502), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n966), .B1(new_n969), .B2(new_n500), .ZN(new_n970));
  XNOR2_X1  g545(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n470), .A2(new_n478), .A3(G40), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n965), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n470), .A2(new_n478), .A3(G40), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT50), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n978), .B(new_n966), .C1(new_n969), .C2(new_n500), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n976), .A2(new_n719), .A3(new_n977), .A4(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT116), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n973), .B1(new_n970), .B2(KEYINPUT50), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT116), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n982), .A2(new_n983), .A3(new_n719), .A4(new_n979), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G1966), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n504), .A2(new_n506), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n496), .A2(new_n499), .ZN(new_n988));
  AOI21_X1  g563(.A(G1384), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OAI211_X1 g564(.A(KEYINPUT115), .B(new_n977), .C1(new_n989), .C2(KEYINPUT45), .ZN(new_n990));
  INV_X1    g565(.A(new_n971), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n994), .B1(G164), .B2(G1384), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT115), .B1(new_n995), .B2(new_n977), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n986), .B1(new_n993), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n985), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n998), .A2(G8), .A3(G286), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT120), .ZN(new_n1000));
  INV_X1    g575(.A(G8), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1001), .B1(new_n985), .B2(new_n997), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT120), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1002), .A2(new_n1003), .A3(G286), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1000), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n985), .A2(G168), .A3(new_n997), .ZN(new_n1006));
  AND2_X1   g581(.A1(KEYINPUT121), .A2(G8), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT51), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1006), .A2(KEYINPUT51), .A3(new_n1007), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT62), .ZN(new_n1013));
  AND3_X1   g588(.A1(new_n1005), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT123), .ZN(new_n1015));
  NAND3_X1  g590(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G1971), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n989), .A2(KEYINPUT45), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n977), .B1(new_n989), .B2(new_n991), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1021), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n982), .A2(new_n783), .A3(new_n979), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(new_n1026), .A3(KEYINPUT114), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n1027), .A2(G8), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT114), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1020), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1001), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n1020), .ZN(new_n1033));
  XNOR2_X1  g608(.A(KEYINPUT112), .B(G1981), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n583), .A2(new_n585), .A3(new_n586), .A4(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n582), .A2(G651), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n516), .A2(G48), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(new_n1038), .A3(new_n584), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(G1981), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT113), .B1(new_n1036), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT49), .ZN(new_n1042));
  OR2_X1    g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  AOI211_X1 g618(.A(KEYINPUT113), .B(KEYINPUT49), .C1(new_n1036), .C2(new_n1040), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1001), .B1(new_n989), .B2(new_n977), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1043), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT52), .B1(G288), .B2(new_n797), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n571), .A2(new_n578), .A3(G1976), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1048), .A2(new_n1046), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT111), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1048), .A2(new_n1046), .A3(KEYINPUT111), .A4(new_n1049), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT52), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1033), .A2(new_n1047), .A3(new_n1054), .A4(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1015), .B1(new_n1031), .B2(new_n1057), .ZN(new_n1058));
  AOI211_X1 g633(.A(new_n1001), .B(new_n1019), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1046), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1056), .B1(new_n1061), .B2(new_n1044), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n1059), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1027), .A2(G8), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1019), .B1(new_n1064), .B2(new_n1029), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1063), .A2(KEYINPUT123), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n982), .A2(new_n979), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n972), .A2(new_n750), .A3(new_n1022), .A4(new_n977), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1067), .A2(new_n711), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n977), .B1(new_n989), .B2(KEYINPUT45), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT115), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1069), .A2(G2078), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1073), .A2(new_n992), .A3(new_n990), .A4(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(G301), .B1(new_n1070), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1058), .A2(new_n1066), .A3(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT126), .B1(new_n1014), .B2(new_n1077), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1031), .A2(new_n1057), .A3(new_n1015), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT123), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1005), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT126), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .A4(new_n1076), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1005), .A2(new_n1012), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT62), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1078), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1047), .A2(new_n797), .A3(new_n794), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1036), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1046), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1047), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1090), .B1(new_n1033), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1020), .B1(new_n1032), .B2(KEYINPUT117), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1093), .B1(KEYINPUT117), .B2(new_n1032), .ZN(new_n1094));
  AND2_X1   g669(.A1(new_n1002), .A2(G168), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1063), .A2(new_n1094), .A3(new_n1095), .A4(KEYINPUT63), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1063), .A2(new_n1095), .A3(new_n1065), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT63), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1092), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1067), .A2(new_n711), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1075), .A2(new_n1101), .A3(new_n1102), .A4(G301), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT124), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT124), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1070), .A2(new_n1105), .A3(G301), .A4(new_n1075), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n972), .A2(new_n977), .A3(new_n1022), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n750), .A2(KEYINPUT53), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1101), .B(new_n1102), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1108), .B1(new_n1111), .B2(G171), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1107), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT125), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT125), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1107), .A2(new_n1112), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1108), .A2(KEYINPUT122), .ZN(new_n1118));
  OR2_X1    g693(.A1(new_n1108), .A2(KEYINPUT122), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1111), .A2(G171), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1118), .B(new_n1119), .C1(new_n1120), .C2(new_n1076), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1117), .A2(new_n1081), .A3(new_n1085), .A4(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1067), .A2(new_n727), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n1124));
  XNOR2_X1  g699(.A(G299), .B(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g700(.A(KEYINPUT56), .B(G2072), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n1126), .B(KEYINPUT118), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1123), .B(new_n1125), .C1(new_n1109), .C2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n977), .B1(new_n989), .B2(new_n978), .ZN(new_n1130));
  INV_X1    g705(.A(new_n979), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n989), .A2(new_n977), .ZN(new_n1133));
  OAI22_X1  g708(.A1(new_n1132), .A2(G1348), .B1(G2067), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1129), .A2(new_n608), .A3(new_n1134), .ZN(new_n1135));
  OAI22_X1  g710(.A1(new_n1132), .A2(G1956), .B1(new_n1109), .B2(new_n1128), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1125), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT60), .ZN(new_n1140));
  OR3_X1    g715(.A1(new_n1134), .A2(new_n1140), .A3(new_n608), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n608), .B1(new_n1134), .B2(new_n1140), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1141), .A2(new_n1142), .B1(new_n1140), .B2(new_n1134), .ZN(new_n1143));
  XOR2_X1   g718(.A(KEYINPUT58), .B(G1341), .Z(new_n1144));
  NAND2_X1  g719(.A1(new_n1133), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1145), .B1(new_n1109), .B2(G1996), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n543), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1147), .B(KEYINPUT59), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT61), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1138), .A2(new_n1129), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1149), .B1(new_n1138), .B2(new_n1129), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1148), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT119), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1143), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1148), .B(KEYINPUT119), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1139), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1100), .B1(new_n1122), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n975), .B1(new_n1087), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(new_n958), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n974), .B1(new_n1159), .B2(new_n744), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n974), .A2(new_n959), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n1161), .A2(KEYINPUT46), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1161), .A2(KEYINPUT46), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1160), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1164), .B(KEYINPUT47), .ZN(new_n1165));
  INV_X1    g740(.A(new_n974), .ZN(new_n1166));
  NOR3_X1   g741(.A1(new_n1166), .A2(G1986), .A3(G290), .ZN(new_n1167));
  XOR2_X1   g742(.A(new_n1167), .B(KEYINPUT48), .Z(new_n1168));
  OAI21_X1  g743(.A(new_n1168), .B1(new_n963), .B2(new_n1166), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n816), .A2(new_n819), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n957), .B1(new_n961), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(new_n974), .ZN(new_n1172));
  AND3_X1   g747(.A1(new_n1165), .A2(new_n1169), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1158), .A2(new_n1173), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g749(.A1(G227), .A2(new_n463), .ZN(new_n1176));
  NAND2_X1  g750(.A1(new_n652), .A2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g751(.A1(G229), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g752(.A1(new_n883), .A2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g753(.A1(new_n944), .A2(new_n946), .ZN(new_n1180));
  NOR2_X1   g754(.A1(new_n1179), .A2(new_n1180), .ZN(G308));
  OR2_X1    g755(.A1(new_n1179), .A2(new_n1180), .ZN(G225));
endmodule


