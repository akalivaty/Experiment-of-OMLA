//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 1 1 1 0 0 0 1 0 0 0 0 0 0 0 1 1 1 1 0 1 1 1 0 1 0 1 1 1 1 0 1 0 0 1 0 1 1 1 0 1 0 1 0 0 1 0 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n780, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n873, new_n874, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984, new_n985;
  AOI21_X1  g000(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(G197gat), .A2(G204gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G197gat), .A2(G204gat), .ZN(new_n205));
  AOI21_X1  g004(.A(new_n202), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G211gat), .B(G218gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  OR3_X1    g007(.A1(new_n206), .A2(new_n208), .A3(KEYINPUT77), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n208), .B1(new_n206), .B2(KEYINPUT77), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G226gat), .A2(G233gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  OR2_X1    g013(.A1(KEYINPUT69), .A2(G183gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(KEYINPUT69), .A2(G183gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n215), .A2(KEYINPUT27), .A3(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(G190gat), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT70), .B1(new_n220), .B2(KEYINPUT28), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT70), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT28), .ZN(new_n223));
  AND2_X1   g022(.A1(KEYINPUT69), .A2(G183gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(KEYINPUT69), .A2(G183gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n218), .B1(new_n226), .B2(KEYINPUT27), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n222), .B(new_n223), .C1(new_n227), .C2(G190gat), .ZN(new_n228));
  XNOR2_X1  g027(.A(KEYINPUT27), .B(G183gat), .ZN(new_n229));
  INV_X1    g028(.A(G190gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n229), .A2(KEYINPUT28), .A3(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n221), .A2(new_n228), .A3(new_n231), .ZN(new_n232));
  OR4_X1    g031(.A1(KEYINPUT71), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n233));
  INV_X1    g032(.A(G169gat), .ZN(new_n234));
  INV_X1    g033(.A(G176gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT71), .B1(new_n236), .B2(KEYINPUT26), .ZN(new_n237));
  NAND2_X1  g036(.A1(G169gat), .A2(G176gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(KEYINPUT66), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n240), .A2(G169gat), .A3(G176gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n236), .A2(KEYINPUT26), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n233), .A2(new_n237), .A3(new_n242), .A4(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(G183gat), .A2(G190gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n232), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n234), .A2(new_n235), .A3(KEYINPUT23), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT23), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(G169gat), .A2(G176gat), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n254), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n251), .A2(new_n242), .A3(new_n253), .A4(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT64), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OR2_X1    g061(.A1(G183gat), .A2(G190gat), .ZN(new_n263));
  AND3_X1   g062(.A1(new_n259), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  OR2_X1    g063(.A1(new_n260), .A2(new_n261), .ZN(new_n265));
  AOI22_X1  g064(.A1(new_n256), .A2(new_n257), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AOI22_X1  g065(.A1(new_n239), .A2(new_n241), .B1(new_n236), .B2(new_n252), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n267), .A2(KEYINPUT67), .A3(new_n255), .A4(new_n251), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT25), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n260), .B1(new_n258), .B2(new_n270), .ZN(new_n271));
  NAND4_X1  g070(.A1(KEYINPUT68), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n271), .B(new_n272), .C1(G190gat), .C2(new_n226), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT25), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n274), .B1(new_n254), .B2(KEYINPUT23), .ZN(new_n275));
  AND3_X1   g074(.A1(new_n273), .A2(new_n267), .A3(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n248), .B1(new_n269), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT29), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n214), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n256), .A2(new_n257), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n280), .A2(new_n268), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(new_n274), .ZN(new_n283));
  INV_X1    g082(.A(new_n276), .ZN(new_n284));
  AOI22_X1  g083(.A1(new_n283), .A2(new_n284), .B1(new_n232), .B2(new_n247), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n285), .A2(new_n213), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n212), .B1(new_n279), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n213), .B1(new_n285), .B2(KEYINPUT29), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n277), .A2(new_n214), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n288), .A2(new_n211), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G8gat), .B(G36gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(G64gat), .B(G92gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT38), .B1(new_n291), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT78), .ZN(new_n297));
  AND3_X1   g096(.A1(new_n288), .A2(new_n211), .A3(new_n289), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n211), .B1(new_n288), .B2(new_n289), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n287), .A2(KEYINPUT78), .A3(new_n290), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(KEYINPUT37), .A3(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT37), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n295), .B1(new_n291), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n296), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n303), .B1(new_n298), .B2(new_n299), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT38), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n287), .A2(KEYINPUT37), .A3(new_n290), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n294), .B(KEYINPUT79), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n306), .A2(new_n307), .A3(new_n308), .A4(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G225gat), .A2(G233gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n311), .B(KEYINPUT81), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G148gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G141gat), .ZN(new_n315));
  INV_X1    g114(.A(G141gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(G148gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT80), .ZN(new_n319));
  INV_X1    g118(.A(G155gat), .ZN(new_n320));
  INV_X1    g119(.A(G162gat), .ZN(new_n321));
  OAI21_X1  g120(.A(KEYINPUT2), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n318), .A2(new_n319), .A3(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G155gat), .B(G162gat), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT80), .B1(new_n315), .B2(new_n317), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n324), .B1(new_n327), .B2(new_n322), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT3), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(G120gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(G113gat), .ZN(new_n331));
  INV_X1    g130(.A(G113gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(G120gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT1), .ZN(new_n335));
  INV_X1    g134(.A(G134gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(G127gat), .ZN(new_n337));
  INV_X1    g136(.A(G127gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(G134gat), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n334), .A2(new_n335), .A3(new_n337), .A4(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n337), .A2(new_n339), .ZN(new_n341));
  XNOR2_X1  g140(.A(G113gat), .B(G120gat), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n341), .B1(new_n342), .B2(KEYINPUT1), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n323), .A2(new_n325), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT3), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n327), .A2(new_n324), .A3(new_n322), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n329), .A2(new_n344), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT4), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n326), .A2(new_n328), .ZN(new_n351));
  AND2_X1   g150(.A1(new_n340), .A2(new_n343), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n345), .A2(new_n347), .ZN(new_n354));
  NOR3_X1   g153(.A1(new_n354), .A2(KEYINPUT4), .A3(new_n344), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n313), .B(new_n349), .C1(new_n353), .C2(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n354), .B(new_n344), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(new_n312), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT5), .ZN(new_n360));
  XNOR2_X1  g159(.A(G1gat), .B(G29gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(G85gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT0), .B(G57gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n362), .B(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT5), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n356), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n360), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n364), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n365), .B1(new_n356), .B2(new_n358), .ZN(new_n369));
  AND2_X1   g168(.A1(new_n348), .A2(new_n344), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT4), .B1(new_n354), .B2(new_n344), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n352), .A2(new_n350), .A3(new_n345), .A4(new_n347), .ZN(new_n372));
  AOI22_X1  g171(.A1(new_n370), .A2(new_n329), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT5), .B1(new_n373), .B2(new_n313), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n368), .B1(new_n369), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT6), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n367), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n369), .A2(new_n374), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n378), .A2(KEYINPUT6), .A3(new_n364), .ZN(new_n379));
  AND2_X1   g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n310), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n305), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n371), .A2(new_n372), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n313), .B1(new_n383), .B2(new_n349), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n385), .B(KEYINPUT39), .C1(new_n312), .C2(new_n357), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT39), .ZN(new_n387));
  AOI211_X1 g186(.A(KEYINPUT86), .B(new_n364), .C1(new_n384), .C2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT86), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n383), .A2(new_n349), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n390), .A2(new_n387), .A3(new_n312), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n389), .B1(new_n391), .B2(new_n368), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n386), .B1(new_n388), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT87), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT40), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n396), .B(new_n386), .C1(new_n388), .C2(new_n392), .ZN(new_n399));
  AOI22_X1  g198(.A1(new_n378), .A2(new_n364), .B1(new_n394), .B2(new_n395), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT30), .B1(new_n291), .B2(new_n295), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT30), .ZN(new_n403));
  AOI211_X1 g202(.A(new_n403), .B(new_n294), .C1(new_n287), .C2(new_n290), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n300), .A2(new_n301), .A3(new_n309), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n401), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AND2_X1   g206(.A1(G228gat), .A2(G233gat), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n348), .A2(new_n278), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(new_n211), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT29), .B1(new_n345), .B2(new_n347), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT82), .ZN(new_n413));
  INV_X1    g212(.A(new_n205), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n414), .A2(new_n203), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n208), .B(new_n413), .C1(new_n202), .C2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT82), .B1(new_n206), .B2(new_n207), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n206), .A2(new_n207), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n412), .A2(new_n419), .B1(new_n354), .B2(KEYINPUT3), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n411), .B1(new_n420), .B2(KEYINPUT83), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n412), .A2(new_n419), .ZN(new_n422));
  AND3_X1   g221(.A1(new_n422), .A2(KEYINPUT83), .A3(new_n329), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n409), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(G22gat), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n209), .A2(new_n278), .A3(new_n210), .ZN(new_n426));
  AND2_X1   g225(.A1(new_n426), .A2(new_n346), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n408), .B(new_n411), .C1(new_n427), .C2(new_n351), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n424), .A2(new_n425), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT84), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n424), .A2(new_n428), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(G22gat), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT84), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n424), .A2(new_n433), .A3(new_n428), .A4(new_n425), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n430), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  XOR2_X1   g234(.A(KEYINPUT31), .B(G50gat), .Z(new_n436));
  XNOR2_X1  g235(.A(G78gat), .B(G106gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n436), .B(new_n437), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n425), .A2(KEYINPUT85), .ZN(new_n439));
  OR2_X1    g238(.A1(new_n431), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n438), .B1(new_n431), .B2(new_n439), .ZN(new_n441));
  AOI22_X1  g240(.A1(new_n435), .A2(new_n438), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NOR3_X1   g241(.A1(new_n382), .A2(new_n407), .A3(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n295), .B1(new_n298), .B2(new_n299), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n403), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n377), .A2(new_n379), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n291), .A2(KEYINPUT30), .A3(new_n295), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n406), .A2(new_n445), .A3(new_n446), .A4(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n442), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT36), .ZN(new_n450));
  NAND2_X1  g249(.A1(G227gat), .A2(G233gat), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n231), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n223), .B1(new_n227), .B2(G190gat), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n453), .B1(new_n454), .B2(KEYINPUT70), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n246), .B1(new_n455), .B2(new_n228), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n276), .B1(new_n282), .B2(new_n274), .ZN(new_n457));
  NOR3_X1   g256(.A1(new_n456), .A2(new_n457), .A3(new_n344), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n283), .A2(new_n284), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n352), .B1(new_n459), .B2(new_n248), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n452), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT32), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT33), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  XOR2_X1   g263(.A(G15gat), .B(G43gat), .Z(new_n465));
  XNOR2_X1  g264(.A(new_n465), .B(KEYINPUT72), .ZN(new_n466));
  XNOR2_X1  g265(.A(G71gat), .B(G99gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n467), .B(KEYINPUT73), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n466), .B(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n462), .A2(new_n464), .A3(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n344), .B1(new_n456), .B2(new_n457), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n248), .B(new_n352), .C1(new_n269), .C2(new_n276), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n451), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n469), .B1(new_n473), .B2(KEYINPUT33), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT32), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n470), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n471), .A2(new_n472), .A3(new_n451), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT34), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT75), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT34), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n471), .A2(new_n472), .A3(new_n482), .A4(new_n451), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n480), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n481), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT74), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n478), .A2(new_n487), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n471), .A2(new_n472), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n489), .A2(KEYINPUT75), .A3(new_n482), .A4(new_n451), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n490), .A2(new_n485), .A3(new_n480), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n470), .A2(new_n491), .A3(KEYINPUT74), .A4(new_n477), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n450), .B1(new_n488), .B2(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(KEYINPUT76), .B(KEYINPUT36), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n484), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n470), .A2(new_n496), .A3(new_n477), .A4(new_n485), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n474), .A2(new_n476), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n471), .A2(new_n472), .ZN(new_n499));
  AOI221_X4 g298(.A(new_n475), .B1(KEYINPUT33), .B2(new_n469), .C1(new_n499), .C2(new_n452), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n491), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n495), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n449), .B1(new_n493), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT35), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n442), .B1(new_n488), .B2(new_n492), .ZN(new_n505));
  INV_X1    g304(.A(new_n448), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n435), .A2(new_n438), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n440), .A2(new_n441), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(new_n504), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n497), .A2(new_n501), .ZN(new_n512));
  NOR3_X1   g311(.A1(new_n511), .A2(new_n448), .A3(new_n512), .ZN(new_n513));
  OAI22_X1  g312(.A1(new_n443), .A2(new_n503), .B1(new_n507), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(G15gat), .B(G22gat), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT16), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n516), .B1(new_n517), .B2(G1gat), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n518), .B1(G1gat), .B2(new_n516), .ZN(new_n519));
  INV_X1    g318(.A(G8gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  AND2_X1   g320(.A1(G71gat), .A2(G78gat), .ZN(new_n522));
  NOR2_X1   g321(.A1(G71gat), .A2(G78gat), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  XOR2_X1   g323(.A(G57gat), .B(G64gat), .Z(new_n525));
  INV_X1    g324(.A(KEYINPUT93), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n525), .B1(KEYINPUT9), .B2(new_n522), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI221_X1 g328(.A(new_n525), .B1(KEYINPUT9), .B2(new_n522), .C1(new_n524), .C2(new_n526), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT21), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n521), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(KEYINPUT95), .ZN(new_n535));
  NAND2_X1  g334(.A1(G231gat), .A2(G233gat), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n536), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n531), .A2(KEYINPUT21), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  XOR2_X1   g340(.A(KEYINPUT94), .B(KEYINPUT19), .Z(new_n542));
  XNOR2_X1  g341(.A(G183gat), .B(G211gat), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n542), .B(new_n543), .Z(new_n544));
  XOR2_X1   g343(.A(G127gat), .B(G155gat), .Z(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT20), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n544), .B(new_n546), .ZN(new_n547));
  OAI211_X1 g346(.A(new_n537), .B(new_n538), .C1(KEYINPUT21), .C2(new_n531), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n541), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n547), .B1(new_n541), .B2(new_n548), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  XOR2_X1   g350(.A(G134gat), .B(G162gat), .Z(new_n552));
  NAND2_X1  g351(.A1(G99gat), .A2(G106gat), .ZN(new_n553));
  INV_X1    g352(.A(G85gat), .ZN(new_n554));
  INV_X1    g353(.A(G92gat), .ZN(new_n555));
  AOI22_X1  g354(.A1(KEYINPUT8), .A2(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT7), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n557), .B1(new_n554), .B2(new_n555), .ZN(new_n558));
  NAND3_X1  g357(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n556), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(KEYINPUT96), .ZN(new_n561));
  XOR2_X1   g360(.A(G99gat), .B(G106gat), .Z(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n560), .A2(KEYINPUT96), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n560), .A2(KEYINPUT96), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n565), .A2(new_n562), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(G43gat), .B(G50gat), .Z(new_n569));
  INV_X1    g368(.A(KEYINPUT15), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT14), .ZN(new_n572));
  INV_X1    g371(.A(G29gat), .ZN(new_n573));
  INV_X1    g372(.A(G36gat), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n575), .A2(KEYINPUT89), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G29gat), .A2(G36gat), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n578), .B1(new_n576), .B2(KEYINPUT89), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n571), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT90), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n571), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n575), .A2(new_n576), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n570), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n583), .A2(new_n584), .A3(new_n578), .A4(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n580), .A2(new_n581), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT91), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n590), .B1(new_n587), .B2(new_n588), .ZN(new_n591));
  OR2_X1    g390(.A1(new_n580), .A2(new_n581), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n592), .A2(KEYINPUT91), .A3(new_n582), .A4(new_n586), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(KEYINPUT92), .B(KEYINPUT17), .Z(new_n595));
  AOI221_X4 g394(.A(new_n568), .B1(KEYINPUT17), .B2(new_n589), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n568), .ZN(new_n597));
  NAND2_X1  g396(.A1(G232gat), .A2(G233gat), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT41), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n552), .B1(new_n596), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n599), .A2(KEYINPUT41), .ZN(new_n603));
  XNOR2_X1  g402(.A(G190gat), .B(G218gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n594), .A2(new_n595), .ZN(new_n606));
  INV_X1    g405(.A(new_n567), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n562), .B1(new_n565), .B2(new_n566), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n589), .A2(KEYINPUT17), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n606), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n552), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n611), .A2(new_n612), .A3(new_n600), .A4(new_n597), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n602), .A2(new_n605), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n605), .B1(new_n602), .B2(new_n613), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n551), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(G113gat), .B(G141gat), .Z(new_n619));
  XNOR2_X1  g418(.A(KEYINPUT88), .B(G197gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(KEYINPUT11), .B(G169gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n623), .B(KEYINPUT12), .Z(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n606), .A2(new_n521), .A3(new_n610), .ZN(new_n626));
  NAND2_X1  g425(.A1(G229gat), .A2(G233gat), .ZN(new_n627));
  INV_X1    g426(.A(new_n521), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n594), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n626), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT18), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n627), .B(KEYINPUT13), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n591), .A2(new_n521), .A3(new_n593), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n633), .B1(new_n629), .B2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n626), .A2(KEYINPUT18), .A3(new_n627), .A4(new_n629), .ZN(new_n637));
  AND4_X1   g436(.A1(new_n625), .A2(new_n632), .A3(new_n636), .A4(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n635), .B1(new_n630), .B2(new_n631), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n625), .B1(new_n639), .B2(new_n637), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G120gat), .B(G148gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(G176gat), .B(G204gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(G230gat), .ZN(new_n645));
  INV_X1    g444(.A(G233gat), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n531), .B1(new_n607), .B2(new_n608), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT97), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n564), .A2(new_n532), .A3(new_n567), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n609), .A2(KEYINPUT97), .A3(new_n532), .ZN(new_n653));
  AOI21_X1  g452(.A(KEYINPUT10), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT10), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n649), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n648), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n652), .A2(new_n647), .A3(new_n653), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n644), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n644), .B1(new_n660), .B2(KEYINPUT98), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT98), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n662), .A2(new_n657), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n641), .A2(new_n667), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n515), .A2(new_n618), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n380), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(G1gat), .ZN(G1324gat));
  NAND3_X1  g470(.A1(new_n406), .A2(new_n445), .A3(new_n447), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT42), .B1(new_n674), .B2(new_n520), .ZN(new_n675));
  NAND2_X1  g474(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n517), .A2(new_n520), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n674), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  MUX2_X1   g477(.A(KEYINPUT42), .B(new_n675), .S(new_n678), .Z(G1325gat));
  INV_X1    g478(.A(new_n512), .ZN(new_n680));
  AOI21_X1  g479(.A(G15gat), .B1(new_n669), .B2(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n478), .A2(new_n487), .ZN(new_n682));
  AOI22_X1  g481(.A1(new_n477), .A2(new_n470), .B1(new_n491), .B2(KEYINPUT74), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT36), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n512), .A2(new_n494), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n687), .A2(G15gat), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n681), .B1(new_n669), .B2(new_n688), .ZN(G1326gat));
  NAND2_X1  g488(.A1(new_n669), .A2(new_n442), .ZN(new_n690));
  XNOR2_X1  g489(.A(KEYINPUT43), .B(G22gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1327gat));
  NOR2_X1   g491(.A1(new_n668), .A2(new_n551), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n617), .A2(KEYINPUT44), .ZN(new_n695));
  AND3_X1   g494(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n672), .A2(new_n696), .ZN(new_n697));
  OAI211_X1 g496(.A(new_n697), .B(new_n510), .C1(new_n305), .C2(new_n381), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n698), .A2(new_n449), .A3(new_n686), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n510), .B1(new_n682), .B2(new_n683), .ZN(new_n700));
  OAI21_X1  g499(.A(KEYINPUT35), .B1(new_n700), .B2(new_n448), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n680), .A2(new_n506), .A3(new_n504), .A4(new_n510), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT99), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n699), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n704), .B1(new_n699), .B2(new_n703), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n695), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n708), .B1(new_n514), .B2(new_n616), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n694), .B1(new_n707), .B2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(G29gat), .B1(new_n712), .B2(new_n446), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n515), .A2(new_n617), .A3(new_n694), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n714), .A2(new_n573), .A3(new_n380), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT45), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n713), .A2(new_n716), .ZN(G1328gat));
  INV_X1    g516(.A(new_n672), .ZN(new_n718));
  OAI21_X1  g517(.A(G36gat), .B1(new_n712), .B2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n714), .A2(new_n574), .A3(new_n672), .ZN(new_n720));
  XOR2_X1   g519(.A(KEYINPUT100), .B(KEYINPUT46), .Z(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n719), .A2(new_n722), .ZN(G1329gat));
  INV_X1    g522(.A(KEYINPUT104), .ZN(new_n724));
  XNOR2_X1  g523(.A(KEYINPUT101), .B(KEYINPUT47), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n512), .A2(G43gat), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n514), .A2(new_n616), .A3(new_n693), .A4(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n695), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n514), .A2(KEYINPUT99), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n699), .A2(new_n703), .A3(new_n704), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n687), .B(new_n693), .C1(new_n732), .C2(new_n709), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(G43gat), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n728), .B1(new_n734), .B2(KEYINPUT102), .ZN(new_n735));
  INV_X1    g534(.A(G43gat), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n736), .B1(new_n711), .B2(new_n687), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT102), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n725), .B1(new_n735), .B2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT103), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n727), .A2(KEYINPUT47), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n741), .B1(new_n737), .B2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n742), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n734), .A2(new_n744), .A3(KEYINPUT103), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n724), .B1(new_n740), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT103), .B1(new_n734), .B2(new_n744), .ZN(new_n748));
  AOI211_X1 g547(.A(new_n741), .B(new_n742), .C1(new_n733), .C2(G43gat), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AND3_X1   g549(.A1(new_n733), .A2(new_n738), .A3(G43gat), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n738), .B1(new_n733), .B2(G43gat), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n751), .A2(new_n752), .A3(new_n728), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n750), .B(KEYINPUT104), .C1(new_n753), .C2(new_n725), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n747), .A2(new_n754), .ZN(G1330gat));
  OAI21_X1  g554(.A(G50gat), .B1(new_n712), .B2(new_n510), .ZN(new_n756));
  INV_X1    g555(.A(G50gat), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n714), .A2(new_n757), .A3(new_n442), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(KEYINPUT48), .B1(new_n758), .B2(KEYINPUT105), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(G1331gat));
  NAND2_X1  g560(.A1(new_n730), .A2(new_n731), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n618), .A2(new_n641), .A3(new_n667), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n380), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g566(.A1(new_n764), .A2(new_n718), .ZN(new_n768));
  NOR2_X1   g567(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n769));
  AND2_X1   g568(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n771), .B1(new_n768), .B2(new_n769), .ZN(G1333gat));
  NAND3_X1  g571(.A1(new_n765), .A2(G71gat), .A3(new_n687), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n773), .A2(KEYINPUT106), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n773), .A2(KEYINPUT106), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n764), .A2(new_n512), .ZN(new_n776));
  OAI22_X1  g575(.A1(new_n774), .A2(new_n775), .B1(G71gat), .B2(new_n776), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g577(.A1(new_n764), .A2(new_n510), .ZN(new_n779));
  XNOR2_X1  g578(.A(KEYINPUT107), .B(G78gat), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n779), .B(new_n780), .ZN(G1335gat));
  INV_X1    g580(.A(new_n551), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n638), .A2(new_n640), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n514), .A2(new_n782), .A3(new_n616), .A4(new_n783), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT51), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n666), .B1(new_n785), .B2(KEYINPUT108), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n786), .B1(KEYINPUT108), .B2(new_n785), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n787), .A2(new_n554), .A3(new_n380), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n707), .A2(new_n710), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n641), .A2(new_n551), .A3(new_n667), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(G85gat), .B1(new_n791), .B2(new_n446), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n788), .A2(new_n792), .ZN(G1336gat));
  INV_X1    g592(.A(new_n791), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n555), .B1(new_n794), .B2(new_n672), .ZN(new_n795));
  NOR4_X1   g594(.A1(new_n785), .A2(G92gat), .A3(new_n718), .A4(new_n667), .ZN(new_n796));
  OAI21_X1  g595(.A(KEYINPUT52), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT110), .B1(new_n794), .B2(new_n672), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT110), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n791), .A2(new_n799), .A3(new_n718), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n798), .A2(new_n555), .A3(new_n800), .ZN(new_n801));
  XNOR2_X1  g600(.A(KEYINPUT109), .B(KEYINPUT52), .ZN(new_n802));
  OR2_X1    g601(.A1(new_n796), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n797), .B1(new_n801), .B2(new_n803), .ZN(G1337gat));
  INV_X1    g603(.A(G99gat), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n787), .A2(new_n805), .A3(new_n680), .ZN(new_n806));
  OAI21_X1  g605(.A(G99gat), .B1(new_n791), .B2(new_n686), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(G1338gat));
  NOR4_X1   g607(.A1(new_n785), .A2(G106gat), .A3(new_n510), .A4(new_n667), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n809), .A2(KEYINPUT53), .ZN(new_n810));
  OAI21_X1  g609(.A(KEYINPUT111), .B1(new_n791), .B2(new_n510), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(G106gat), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n791), .A2(KEYINPUT111), .A3(new_n510), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n810), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(G106gat), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n815), .B1(new_n794), .B2(new_n442), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT53), .B1(new_n816), .B2(new_n809), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n814), .A2(new_n817), .ZN(G1339gat));
  NAND4_X1  g617(.A1(new_n551), .A2(new_n783), .A3(new_n617), .A4(new_n667), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821));
  INV_X1    g620(.A(new_n656), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n652), .A2(new_n653), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n647), .B(new_n822), .C1(new_n823), .C2(KEYINPUT10), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n824), .A2(KEYINPUT54), .A3(new_n657), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n826), .B(new_n648), .C1(new_n654), .C2(new_n656), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n644), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n821), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n827), .A2(new_n644), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n824), .A2(KEYINPUT54), .A3(new_n657), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n830), .A2(KEYINPUT55), .A3(new_n831), .ZN(new_n832));
  AND4_X1   g631(.A1(new_n616), .A2(new_n829), .A3(new_n665), .A4(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n639), .A2(new_n625), .A3(new_n637), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n627), .B1(new_n626), .B2(new_n629), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n629), .A2(new_n634), .A3(new_n633), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n623), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n833), .A2(new_n839), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n666), .A2(new_n834), .A3(new_n837), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n830), .A2(KEYINPUT55), .A3(new_n831), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT55), .B1(new_n830), .B2(new_n831), .ZN(new_n843));
  INV_X1    g642(.A(new_n665), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n841), .B1(new_n845), .B2(new_n641), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n840), .B1(new_n846), .B2(new_n616), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n820), .B1(new_n847), .B2(new_n782), .ZN(new_n848));
  OAI21_X1  g647(.A(KEYINPUT112), .B1(new_n848), .B2(new_n442), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n849), .A2(new_n680), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n672), .A2(new_n446), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n829), .A2(new_n665), .A3(new_n832), .ZN(new_n852));
  OAI22_X1  g651(.A1(new_n852), .A2(new_n783), .B1(new_n667), .B2(new_n838), .ZN(new_n853));
  AOI22_X1  g652(.A1(new_n853), .A2(new_n617), .B1(new_n839), .B2(new_n833), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n819), .B1(new_n854), .B2(new_n551), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT112), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n855), .A2(new_n856), .A3(new_n510), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n850), .A2(new_n641), .A3(new_n851), .A4(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(KEYINPUT113), .A3(G113gat), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(KEYINPUT113), .B1(new_n858), .B2(G113gat), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n848), .A2(new_n446), .A3(new_n700), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n718), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n641), .A2(new_n332), .ZN(new_n864));
  OAI22_X1  g663(.A1(new_n860), .A2(new_n861), .B1(new_n863), .B2(new_n864), .ZN(G1340gat));
  NAND4_X1  g664(.A1(new_n850), .A2(new_n666), .A3(new_n851), .A4(new_n857), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT114), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n867), .A3(G120gat), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n867), .B1(new_n866), .B2(G120gat), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n666), .A2(new_n330), .ZN(new_n871));
  OAI22_X1  g670(.A1(new_n869), .A2(new_n870), .B1(new_n863), .B2(new_n871), .ZN(G1341gat));
  OAI21_X1  g671(.A(new_n338), .B1(new_n863), .B2(new_n782), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n850), .A2(new_n851), .A3(new_n857), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n551), .A2(G127gat), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(G1342gat));
  NAND2_X1  g676(.A1(new_n718), .A2(new_n616), .ZN(new_n878));
  XOR2_X1   g677(.A(new_n878), .B(KEYINPUT115), .Z(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n862), .A2(new_n336), .A3(new_n880), .ZN(new_n881));
  XOR2_X1   g680(.A(new_n881), .B(KEYINPUT56), .Z(new_n882));
  OAI21_X1  g681(.A(G134gat), .B1(new_n874), .B2(new_n617), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(G1343gat));
  NAND2_X1  g683(.A1(new_n686), .A2(new_n851), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n853), .A2(new_n617), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT117), .ZN(new_n887));
  AOI22_X1  g686(.A1(new_n886), .A2(new_n887), .B1(new_n839), .B2(new_n833), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n853), .A2(KEYINPUT117), .A3(new_n617), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n551), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI211_X1 g689(.A(KEYINPUT57), .B(new_n442), .C1(new_n890), .C2(new_n820), .ZN(new_n891));
  XNOR2_X1  g690(.A(KEYINPUT116), .B(KEYINPUT57), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n892), .B1(new_n848), .B2(new_n510), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n885), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n316), .B1(new_n894), .B2(new_n641), .ZN(new_n895));
  NAND2_X1  g694(.A1(KEYINPUT118), .A2(KEYINPUT58), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n687), .A2(new_n510), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n855), .A2(new_n380), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n718), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n641), .A2(new_n316), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n896), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g700(.A1(KEYINPUT118), .A2(KEYINPUT58), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT119), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  OR3_X1    g703(.A1(new_n895), .A2(new_n901), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n895), .B2(new_n901), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(G1344gat));
  INV_X1    g706(.A(new_n899), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(new_n314), .A3(new_n666), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT59), .ZN(new_n910));
  AND3_X1   g709(.A1(new_n855), .A2(new_n442), .A3(new_n892), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT57), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n912), .B1(new_n855), .B2(new_n442), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n666), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n915), .A2(new_n885), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n910), .B1(new_n916), .B2(G148gat), .ZN(new_n917));
  AOI211_X1 g716(.A(KEYINPUT59), .B(new_n314), .C1(new_n894), .C2(new_n666), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n909), .B1(new_n917), .B2(new_n918), .ZN(G1345gat));
  AOI21_X1  g718(.A(G155gat), .B1(new_n908), .B2(new_n551), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n782), .A2(new_n320), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n894), .B2(new_n921), .ZN(G1346gat));
  NAND3_X1  g721(.A1(new_n898), .A2(new_n321), .A3(new_n880), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n894), .A2(new_n616), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n923), .B1(new_n925), .B2(new_n321), .ZN(G1347gat));
  NOR2_X1   g725(.A1(new_n718), .A2(new_n380), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n927), .A2(KEYINPUT120), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n927), .A2(KEYINPUT120), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n849), .A2(new_n680), .A3(new_n857), .A4(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(G169gat), .B1(new_n931), .B2(new_n783), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n855), .A2(new_n927), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n933), .A2(new_n505), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n934), .A2(new_n234), .A3(new_n641), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n932), .A2(new_n935), .ZN(G1348gat));
  OAI21_X1  g735(.A(G176gat), .B1(new_n931), .B2(new_n667), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n934), .A2(new_n235), .A3(new_n666), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT121), .ZN(G1349gat));
  OAI21_X1  g739(.A(new_n226), .B1(new_n931), .B2(new_n782), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n934), .A2(new_n229), .A3(new_n551), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g743(.A(G190gat), .B1(new_n931), .B2(new_n617), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT122), .ZN(new_n946));
  OR3_X1    g745(.A1(new_n945), .A2(new_n946), .A3(KEYINPUT61), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n946), .B1(new_n945), .B2(KEYINPUT61), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n945), .A2(KEYINPUT61), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n934), .A2(new_n230), .A3(new_n616), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(G1351gat));
  NAND2_X1  g751(.A1(new_n933), .A2(new_n897), .ZN(new_n953));
  OR3_X1    g752(.A1(new_n953), .A2(G197gat), .A3(new_n783), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n928), .A2(new_n687), .A3(new_n929), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n911), .A2(new_n913), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(new_n641), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n958), .A2(KEYINPUT123), .ZN(new_n959));
  OAI21_X1  g758(.A(G197gat), .B1(new_n958), .B2(KEYINPUT123), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n954), .B1(new_n959), .B2(new_n960), .ZN(G1352gat));
  NOR3_X1   g760(.A1(new_n953), .A2(G204gat), .A3(new_n667), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n962), .B(KEYINPUT62), .ZN(new_n963));
  OAI21_X1  g762(.A(G204gat), .B1(new_n915), .B2(new_n956), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(G1353gat));
  INV_X1    g764(.A(G211gat), .ZN(new_n966));
  OAI21_X1  g765(.A(KEYINPUT57), .B1(new_n848), .B2(new_n510), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n855), .A2(new_n442), .A3(new_n892), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n967), .A2(new_n551), .A3(new_n968), .A4(new_n955), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT124), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n966), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n914), .A2(KEYINPUT124), .A3(new_n551), .A4(new_n955), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n971), .A2(new_n972), .A3(KEYINPUT63), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(KEYINPUT125), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n971), .A2(new_n972), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT63), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT125), .ZN(new_n978));
  NAND4_X1  g777(.A1(new_n971), .A2(new_n972), .A3(new_n978), .A4(KEYINPUT63), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n974), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  NAND4_X1  g779(.A1(new_n933), .A2(new_n966), .A3(new_n551), .A4(new_n897), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(G1354gat));
  NAND3_X1  g781(.A1(new_n957), .A2(G218gat), .A3(new_n616), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n953), .A2(new_n617), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n983), .B1(G218gat), .B2(new_n984), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n985), .B(KEYINPUT126), .ZN(G1355gat));
endmodule


