//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 0 1 1 0 0 0 1 0 0 0 1 0 0 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 1 1 0 0 0 1 1 0 0 1 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n547, new_n548, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n606, new_n608, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1138, new_n1139;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G2106), .ZN(new_n455));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  OAI22_X1  g031(.A1(new_n451), .A2(new_n455), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT65), .Z(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(new_n459), .A2(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G101), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(new_n459), .ZN(new_n463));
  INV_X1    g038(.A(G137), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n462), .A2(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n459), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n465), .A2(new_n468), .ZN(G160));
  AND2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G136), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n472), .A2(new_n459), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  OR2_X1    g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n477), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n474), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G162));
  OAI21_X1  g055(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G114), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(new_n482), .B2(G2105), .ZN(new_n483));
  AND2_X1   g058(.A1(G126), .A2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n484), .B1(new_n470), .B2(new_n471), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT66), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT66), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(new_n484), .C1(new_n470), .C2(new_n471), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n483), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  OAI211_X1 g064(.A(G138), .B(new_n459), .C1(new_n470), .C2(new_n471), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n462), .A2(new_n492), .A3(G138), .A4(new_n459), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G164));
  INV_X1    g071(.A(KEYINPUT67), .ZN(new_n497));
  INV_X1    g072(.A(G543), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(KEYINPUT5), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(KEYINPUT67), .A3(G543), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n499), .A2(new_n501), .B1(KEYINPUT5), .B2(new_n498), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n502), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n502), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n506));
  OR2_X1    g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n505), .A2(new_n511), .ZN(G166));
  NAND3_X1  g087(.A1(new_n502), .A2(G63), .A3(G651), .ZN(new_n513));
  XOR2_X1   g088(.A(new_n513), .B(KEYINPUT68), .Z(new_n514));
  NAND2_X1  g089(.A1(new_n499), .A2(new_n501), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n498), .A2(KEYINPUT5), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n515), .A2(new_n516), .A3(new_n509), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G89), .ZN(new_n519));
  XOR2_X1   g094(.A(KEYINPUT71), .B(KEYINPUT7), .Z(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n520), .B(new_n521), .ZN(new_n522));
  XOR2_X1   g097(.A(KEYINPUT70), .B(G51), .Z(new_n523));
  NAND2_X1  g098(.A1(new_n509), .A2(KEYINPUT69), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT69), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n507), .A2(new_n525), .A3(new_n508), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n524), .A2(G543), .A3(new_n526), .ZN(new_n527));
  OAI211_X1 g102(.A(new_n519), .B(new_n522), .C1(new_n523), .C2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n514), .A2(new_n528), .ZN(G168));
  INV_X1    g104(.A(G52), .ZN(new_n530));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n527), .A2(new_n530), .B1(new_n531), .B2(new_n517), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n502), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n504), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n532), .A2(new_n534), .ZN(G171));
  AOI22_X1  g110(.A1(new_n502), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT72), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n536), .A2(new_n537), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n538), .A2(G651), .A3(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n527), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n541), .A2(G43), .B1(new_n518), .B2(G81), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  NAND4_X1  g120(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(G188));
  INV_X1    g124(.A(KEYINPUT9), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n541), .A2(new_n550), .A3(G53), .ZN(new_n551));
  INV_X1    g126(.A(G53), .ZN(new_n552));
  OAI21_X1  g127(.A(KEYINPUT9), .B1(new_n527), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n517), .A2(KEYINPUT73), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT73), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n502), .A2(new_n556), .A3(new_n509), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n555), .A2(G91), .A3(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n502), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n559), .A2(new_n504), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n554), .A2(new_n558), .A3(new_n560), .ZN(G299));
  INV_X1    g136(.A(G171), .ZN(G301));
  INV_X1    g137(.A(G168), .ZN(G286));
  INV_X1    g138(.A(G166), .ZN(G303));
  NAND3_X1  g139(.A1(new_n555), .A2(G87), .A3(new_n557), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n502), .B2(G74), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n524), .A2(G49), .A3(G543), .A4(new_n526), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(G288));
  NAND2_X1  g143(.A1(new_n502), .A2(G61), .ZN(new_n569));
  NAND2_X1  g144(.A1(G73), .A2(G543), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G651), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n555), .A2(G86), .A3(new_n557), .ZN(new_n573));
  AND2_X1   g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n509), .A2(G48), .A3(G543), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(new_n577));
  OAI21_X1  g152(.A(KEYINPUT74), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT74), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n574), .A2(new_n579), .A3(new_n576), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n580), .ZN(G305));
  INV_X1    g156(.A(G47), .ZN(new_n582));
  INV_X1    g157(.A(G85), .ZN(new_n583));
  OAI22_X1  g158(.A1(new_n527), .A2(new_n582), .B1(new_n583), .B2(new_n517), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n502), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n504), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n502), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n590), .A2(new_n504), .ZN(new_n591));
  INV_X1    g166(.A(G54), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n592), .B2(new_n527), .ZN(new_n593));
  NAND4_X1  g168(.A1(new_n555), .A2(KEYINPUT10), .A3(G92), .A4(new_n557), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n555), .A2(new_n557), .ZN(new_n596));
  INV_X1    g171(.A(G92), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n593), .B1(new_n594), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n589), .B1(new_n599), .B2(G868), .ZN(G284));
  OAI21_X1  g175(.A(new_n589), .B1(new_n599), .B2(G868), .ZN(G321));
  NAND2_X1  g176(.A1(G286), .A2(G868), .ZN(new_n602));
  AND3_X1   g177(.A1(new_n554), .A2(new_n558), .A3(new_n560), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(G868), .B2(new_n603), .ZN(G297));
  OAI21_X1  g179(.A(new_n602), .B1(G868), .B2(new_n603), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n599), .B1(new_n606), .B2(G860), .ZN(G148));
  NOR2_X1   g182(.A1(new_n544), .A2(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n599), .A2(new_n606), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(G868), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT75), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g187(.A1(new_n462), .A2(new_n460), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT13), .ZN(new_n615));
  INV_X1    g190(.A(G2100), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT77), .Z(new_n618));
  NOR2_X1   g193(.A1(new_n615), .A2(new_n616), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT76), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n473), .A2(G135), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n475), .A2(G123), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n459), .A2(G111), .ZN(new_n623));
  OAI21_X1  g198(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n621), .B(new_n622), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(G2096), .Z(new_n626));
  NAND3_X1  g201(.A1(new_n618), .A2(new_n620), .A3(new_n626), .ZN(G156));
  INV_X1    g202(.A(KEYINPUT14), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2427), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2430), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2435), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n628), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(new_n631), .B2(new_n630), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2451), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT16), .ZN(new_n635));
  XNOR2_X1  g210(.A(G1341), .B(G1348), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n633), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  AND3_X1   g216(.A1(new_n640), .A2(G14), .A3(new_n641), .ZN(G401));
  XOR2_X1   g217(.A(KEYINPUT78), .B(KEYINPUT18), .Z(new_n643));
  XOR2_X1   g218(.A(G2084), .B(G2090), .Z(new_n644));
  XNOR2_X1  g219(.A(G2067), .B(G2678), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(KEYINPUT17), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n644), .A2(new_n645), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n643), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2072), .B(G2078), .Z(new_n650));
  INV_X1    g225(.A(new_n643), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n650), .B1(new_n646), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n649), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2096), .B(G2100), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(G227));
  XNOR2_X1  g230(.A(G1956), .B(G2474), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT80), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1961), .B(G1966), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(KEYINPUT79), .B(KEYINPUT19), .Z(new_n661));
  XNOR2_X1  g236(.A(G1971), .B(G1976), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT20), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n658), .A2(new_n659), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n660), .A2(new_n663), .A3(new_n667), .ZN(new_n668));
  OAI211_X1 g243(.A(new_n666), .B(new_n668), .C1(new_n663), .C2(new_n667), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1991), .B(G1996), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1981), .B(G1986), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(G229));
  OAI21_X1  g250(.A(KEYINPUT95), .B1(G29), .B2(G32), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n460), .A2(KEYINPUT93), .A3(G105), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n459), .A2(G105), .A3(G2104), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT93), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI22_X1  g255(.A1(new_n473), .A2(G141), .B1(new_n677), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n475), .A2(G129), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT94), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT26), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(G29), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  MUX2_X1   g265(.A(new_n676), .B(KEYINPUT95), .S(new_n690), .Z(new_n691));
  XOR2_X1   g266(.A(KEYINPUT27), .B(G1996), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G21), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G168), .B2(new_n694), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G1966), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT25), .ZN(new_n698));
  NAND2_X1  g273(.A1(G103), .A2(G2104), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n698), .B1(new_n699), .B2(G2105), .ZN(new_n700));
  NAND4_X1  g275(.A1(new_n459), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n701));
  AOI22_X1  g276(.A1(new_n473), .A2(G139), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  AOI22_X1  g277(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n459), .B2(new_n703), .ZN(new_n704));
  MUX2_X1   g279(.A(G33), .B(new_n704), .S(G29), .Z(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT92), .Z(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G2072), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT31), .B(G11), .Z(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT30), .B(G28), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n708), .B1(new_n689), .B2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT81), .B(G29), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT24), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n712), .A2(G34), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(G34), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n711), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G160), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(new_n689), .ZN(new_n717));
  INV_X1    g292(.A(G2084), .ZN(new_n718));
  OAI221_X1 g293(.A(new_n710), .B1(new_n625), .B2(new_n711), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(new_n718), .B2(new_n717), .ZN(new_n720));
  NAND4_X1  g295(.A1(new_n693), .A2(new_n697), .A3(new_n707), .A4(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n696), .A2(G1966), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT96), .ZN(new_n723));
  INV_X1    g298(.A(new_n711), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n724), .A2(G27), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G164), .B2(new_n724), .ZN(new_n726));
  INV_X1    g301(.A(G2078), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n694), .A2(G5), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G171), .B2(new_n694), .ZN(new_n730));
  INV_X1    g305(.A(G1961), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n728), .B(new_n732), .C1(new_n706), .C2(G2072), .ZN(new_n733));
  NOR3_X1   g308(.A1(new_n721), .A2(new_n723), .A3(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT97), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR4_X1   g311(.A1(new_n721), .A2(KEYINPUT97), .A3(new_n723), .A4(new_n733), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT87), .ZN(new_n738));
  OR3_X1    g313(.A1(new_n738), .A2(G4), .A3(G16), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n738), .B1(G4), .B2(G16), .ZN(new_n740));
  INV_X1    g315(.A(new_n599), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n739), .B(new_n740), .C1(new_n741), .C2(new_n694), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT88), .ZN(new_n743));
  INV_X1    g318(.A(G1348), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n544), .A2(G16), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G16), .B2(G19), .ZN(new_n747));
  INV_X1    g322(.A(G1341), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n724), .A2(G35), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G162), .B2(new_n724), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT29), .B(G2090), .Z(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n711), .A2(G26), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT28), .Z(new_n755));
  NAND2_X1  g330(.A1(new_n473), .A2(G140), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT89), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n475), .A2(G128), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT90), .ZN(new_n759));
  OR2_X1    g334(.A1(G104), .A2(G2105), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n760), .B(G2104), .C1(G116), .C2(new_n459), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT91), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n757), .A2(new_n759), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n755), .B1(new_n763), .B2(G29), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G2067), .ZN(new_n765));
  AND3_X1   g340(.A1(new_n749), .A2(new_n753), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n694), .A2(G20), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT23), .Z(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G299), .B2(G16), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1956), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n766), .B(new_n770), .C1(new_n748), .C2(new_n747), .ZN(new_n771));
  NOR4_X1   g346(.A1(new_n736), .A2(new_n737), .A3(new_n745), .A4(new_n771), .ZN(new_n772));
  MUX2_X1   g347(.A(G6), .B(G305), .S(G16), .Z(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT32), .B(G1981), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT83), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n773), .B(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(G16), .A2(G22), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G166), .B2(G16), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT84), .B(G1971), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n778), .B(new_n779), .Z(new_n780));
  AND2_X1   g355(.A1(new_n780), .A2(KEYINPUT85), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n780), .A2(KEYINPUT85), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n694), .A2(G23), .ZN(new_n783));
  INV_X1    g358(.A(G288), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(new_n694), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT33), .B(G1976), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NOR3_X1   g362(.A1(new_n781), .A2(new_n782), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n776), .A2(new_n788), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT82), .B(KEYINPUT34), .Z(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n776), .A2(new_n790), .A3(new_n788), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n587), .A2(new_n694), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n694), .B2(G24), .ZN(new_n795));
  INV_X1    g370(.A(G1986), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n473), .A2(G131), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n475), .A2(G119), .ZN(new_n799));
  OR2_X1    g374(.A1(G95), .A2(G2105), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n800), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n798), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n803), .A2(new_n724), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G25), .B2(new_n724), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT35), .B(G1991), .Z(new_n806));
  OR2_X1    g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT86), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT36), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n807), .B(new_n808), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n795), .A2(new_n796), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n792), .A2(new_n793), .A3(new_n797), .A4(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(KEYINPUT86), .A2(KEYINPUT36), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n814), .A2(new_n815), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n772), .A2(new_n816), .A3(new_n817), .ZN(G150));
  INV_X1    g393(.A(G150), .ZN(G311));
  NAND2_X1  g394(.A1(new_n599), .A2(G559), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT38), .Z(new_n821));
  NAND2_X1  g396(.A1(new_n502), .A2(G67), .ZN(new_n822));
  NAND2_X1  g397(.A1(G80), .A2(G543), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT98), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n504), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n825), .B2(new_n824), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n541), .A2(G55), .B1(new_n518), .B2(G93), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(new_n543), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n827), .A2(new_n540), .A3(new_n542), .A4(new_n828), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n821), .B(new_n832), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n833), .A2(KEYINPUT39), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n833), .A2(KEYINPUT39), .ZN(new_n835));
  NOR3_X1   g410(.A1(new_n834), .A2(new_n835), .A3(G860), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n829), .A2(G860), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT37), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n836), .A2(new_n838), .ZN(G145));
  NAND2_X1  g414(.A1(new_n473), .A2(G142), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT100), .Z(new_n841));
  INV_X1    g416(.A(G118), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n842), .A2(KEYINPUT101), .A3(G2105), .ZN(new_n843));
  AOI21_X1  g418(.A(KEYINPUT101), .B1(new_n842), .B2(G2105), .ZN(new_n844));
  OAI21_X1  g419(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n475), .A2(G130), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n841), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n802), .B(new_n614), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT102), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n763), .B(G164), .ZN(new_n852));
  AND2_X1   g427(.A1(new_n852), .A2(new_n704), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n852), .A2(new_n704), .ZN(new_n854));
  OR3_X1    g429(.A1(new_n853), .A2(new_n854), .A3(new_n688), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n688), .B1(new_n853), .B2(new_n854), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n851), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  XOR2_X1   g432(.A(G160), .B(KEYINPUT99), .Z(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(G162), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n625), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n855), .A2(new_n856), .A3(new_n850), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AND3_X1   g438(.A1(new_n855), .A2(new_n856), .A3(new_n851), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n860), .B1(new_n864), .B2(new_n857), .ZN(new_n865));
  XOR2_X1   g440(.A(KEYINPUT103), .B(G37), .Z(new_n866));
  NAND3_X1  g441(.A1(new_n863), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g443(.A(new_n832), .B(new_n609), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n741), .A2(KEYINPUT104), .A3(G299), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT104), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n603), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(G299), .A2(KEYINPUT104), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n872), .A2(new_n599), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n869), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT41), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n870), .A2(new_n874), .A3(KEYINPUT41), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n876), .B1(new_n880), .B2(new_n869), .ZN(new_n881));
  OR2_X1    g456(.A1(new_n881), .A2(KEYINPUT42), .ZN(new_n882));
  XOR2_X1   g457(.A(G166), .B(G288), .Z(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n578), .A2(new_n580), .A3(G290), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(G290), .B1(new_n578), .B2(new_n580), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n884), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n887), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n889), .A2(new_n883), .A3(new_n885), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n891), .A2(KEYINPUT105), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n881), .A2(KEYINPUT42), .ZN(new_n893));
  AND3_X1   g468(.A1(new_n882), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n892), .B1(new_n882), .B2(new_n893), .ZN(new_n895));
  OAI21_X1  g470(.A(G868), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n829), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n896), .B1(G868), .B2(new_n897), .ZN(G295));
  OAI21_X1  g473(.A(new_n896), .B1(G868), .B2(new_n897), .ZN(G331));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n830), .A2(G301), .A3(new_n831), .ZN(new_n901));
  AOI21_X1  g476(.A(G301), .B1(new_n830), .B2(new_n831), .ZN(new_n902));
  OAI21_X1  g477(.A(G286), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n832), .A2(G171), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n830), .A2(G301), .A3(new_n831), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n904), .A2(G168), .A3(new_n905), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n878), .A2(new_n879), .A3(new_n903), .A4(new_n906), .ZN(new_n907));
  AND2_X1   g482(.A1(new_n903), .A2(new_n906), .ZN(new_n908));
  OAI211_X1 g483(.A(new_n907), .B(new_n891), .C1(new_n908), .C2(new_n875), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n875), .B1(new_n903), .B2(new_n906), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n910), .B1(new_n880), .B2(new_n908), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n883), .B1(new_n889), .B2(new_n885), .ZN(new_n912));
  NOR3_X1   g487(.A1(new_n886), .A2(new_n884), .A3(new_n887), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT106), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT106), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n888), .A2(new_n890), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n909), .B(new_n866), .C1(new_n911), .C2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n900), .B1(new_n918), .B2(KEYINPUT43), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n914), .A2(new_n916), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n907), .B1(new_n908), .B2(new_n875), .ZN(new_n921));
  AOI21_X1  g496(.A(G37), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT43), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(new_n923), .A3(new_n909), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n919), .A2(KEYINPUT107), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT107), .B1(new_n919), .B2(new_n924), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n923), .B1(new_n922), .B2(new_n909), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n918), .A2(KEYINPUT43), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI22_X1  g504(.A1(new_n925), .A2(new_n926), .B1(KEYINPUT44), .B2(new_n929), .ZN(G397));
  INV_X1    g505(.A(G1384), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n495), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT45), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(G160), .A2(G40), .ZN(new_n935));
  OR3_X1    g510(.A1(new_n934), .A2(KEYINPUT108), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(KEYINPUT108), .B1(new_n934), .B2(new_n935), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n763), .B(G2067), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  XOR2_X1   g515(.A(new_n940), .B(KEYINPUT109), .Z(new_n941));
  XNOR2_X1  g516(.A(new_n688), .B(G1996), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n941), .B1(new_n938), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n938), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n802), .B(new_n806), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n945), .B(KEYINPUT110), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n943), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n587), .B(new_n796), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n947), .B1(new_n938), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(G8), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT111), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n951), .B1(new_n495), .B2(new_n931), .ZN(new_n952));
  AOI211_X1 g527(.A(KEYINPUT111), .B(G1384), .C1(new_n489), .C2(new_n494), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AND2_X1   g529(.A1(G160), .A2(G40), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n950), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n956), .B(KEYINPUT116), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n952), .A2(new_n953), .A3(new_n935), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n577), .A2(G1981), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n572), .A2(new_n573), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n504), .B1(new_n569), .B2(new_n570), .ZN(new_n961));
  INV_X1    g536(.A(G86), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n576), .B1(new_n517), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(G1981), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(KEYINPUT49), .B1(new_n960), .B2(new_n964), .ZN(new_n965));
  NOR3_X1   g540(.A1(new_n958), .A2(new_n965), .A3(new_n950), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n960), .A2(KEYINPUT49), .A3(new_n964), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT115), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT115), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n960), .A2(new_n969), .A3(new_n964), .A4(KEYINPUT49), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  AOI211_X1 g546(.A(G1976), .B(G288), .C1(new_n966), .C2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n960), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n957), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(G1384), .B1(new_n489), .B2(new_n494), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT50), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n977), .B(KEYINPUT113), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n935), .A2(G2090), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT112), .B1(new_n954), .B2(new_n976), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT112), .ZN(new_n981));
  NOR4_X1   g556(.A1(new_n952), .A2(new_n953), .A3(new_n981), .A4(KEYINPUT50), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n978), .B(new_n979), .C1(new_n980), .C2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G1971), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n955), .B1(new_n932), .B2(new_n933), .ZN(new_n985));
  INV_X1    g560(.A(new_n934), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n984), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n950), .B1(new_n983), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(G166), .A2(new_n950), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n989), .B(KEYINPUT55), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n932), .A2(KEYINPUT111), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n975), .A2(new_n951), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n992), .A2(new_n955), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n784), .A2(G1976), .ZN(new_n995));
  INV_X1    g570(.A(G1976), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT52), .B1(G288), .B2(new_n996), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n994), .A2(new_n995), .A3(G8), .A4(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT114), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n956), .A2(KEYINPUT114), .A3(new_n995), .A4(new_n997), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n994), .A2(new_n995), .A3(G8), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n966), .A2(new_n971), .B1(new_n1003), .B2(KEYINPUT52), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n974), .B1(new_n991), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n935), .B1(new_n976), .B2(new_n975), .ZN(new_n1007));
  INV_X1    g582(.A(G2090), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1007), .B(new_n1008), .C1(new_n954), .C2(new_n976), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n987), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n990), .B1(new_n1010), .B2(G8), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1011), .B1(new_n988), .B2(new_n990), .ZN(new_n1012));
  XNOR2_X1  g587(.A(KEYINPUT124), .B(KEYINPUT53), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n985), .A2(new_n986), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1013), .B1(new_n1014), .B2(new_n727), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n955), .B(new_n978), .C1(new_n980), .C2(new_n982), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1015), .B1(new_n1016), .B2(new_n731), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n932), .A2(new_n933), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1018), .A2(new_n935), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1019), .B1(KEYINPUT45), .B2(new_n954), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n727), .A2(KEYINPUT53), .ZN(new_n1021));
  OR2_X1    g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(G301), .B1(new_n1017), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT117), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1002), .A2(new_n1004), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1024), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1012), .B(new_n1023), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  XOR2_X1   g603(.A(KEYINPUT123), .B(KEYINPUT51), .Z(new_n1029));
  NAND2_X1  g604(.A1(G286), .A2(G8), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n1030), .B(KEYINPUT122), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n935), .A2(G2084), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n978), .B(new_n1033), .C1(new_n980), .C2(new_n982), .ZN(new_n1034));
  INV_X1    g609(.A(G1966), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1020), .A2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n950), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1029), .B1(new_n1032), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(G8), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1040), .A2(KEYINPUT51), .A3(new_n1031), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1032), .A2(new_n1039), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1038), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1028), .B1(KEYINPUT62), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT62), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1038), .A2(new_n1041), .A3(new_n1045), .A4(new_n1042), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1006), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  AOI211_X1 g622(.A(new_n950), .B(G286), .C1(new_n1034), .C2(new_n1036), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1012), .B(new_n1048), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT63), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT118), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT118), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1049), .A2(new_n1053), .A3(new_n1050), .ZN(new_n1054));
  OR2_X1    g629(.A1(new_n988), .A2(new_n990), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1005), .A2(new_n1050), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1055), .A2(new_n1056), .A3(new_n991), .A4(new_n1048), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1052), .A2(new_n1054), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1047), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1005), .A2(KEYINPUT117), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(new_n1025), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n1061), .A2(new_n1012), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1018), .ZN(new_n1064));
  XOR2_X1   g639(.A(new_n465), .B(KEYINPUT125), .Z(new_n1065));
  INV_X1    g640(.A(KEYINPUT126), .ZN(new_n1066));
  OAI211_X1 g641(.A(KEYINPUT53), .B(G40), .C1(new_n1066), .C2(G2078), .ZN(new_n1067));
  AOI211_X1 g642(.A(new_n1067), .B(new_n468), .C1(new_n1066), .C2(G2078), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1064), .A2(new_n934), .A3(new_n1065), .A4(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1017), .A2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1070), .A2(G171), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1063), .B1(new_n1071), .B2(new_n1023), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(G171), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1017), .A2(G301), .A3(new_n1022), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1073), .A2(KEYINPUT54), .A3(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1062), .A2(new_n1072), .A3(new_n1075), .A4(new_n1043), .ZN(new_n1076));
  XNOR2_X1  g651(.A(KEYINPUT56), .B(G2072), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1014), .A2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n955), .B1(new_n932), .B2(KEYINPUT50), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n992), .A2(new_n993), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1079), .B1(new_n1080), .B2(KEYINPUT50), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1078), .B1(new_n1081), .B2(G1956), .ZN(new_n1082));
  XNOR2_X1  g657(.A(G299), .B(KEYINPUT57), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT61), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1019), .A2(new_n934), .ZN(new_n1087));
  XNOR2_X1  g662(.A(KEYINPUT58), .B(G1341), .ZN(new_n1088));
  OAI22_X1  g663(.A1(new_n1087), .A2(G1996), .B1(new_n958), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n1090));
  AND4_X1   g665(.A1(KEYINPUT121), .A2(new_n1089), .A3(new_n1090), .A4(new_n544), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT121), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n543), .B1(new_n1092), .B2(KEYINPUT59), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1089), .A2(new_n1093), .B1(KEYINPUT121), .B2(new_n1090), .ZN(new_n1094));
  OAI22_X1  g669(.A1(new_n1085), .A2(new_n1086), .B1(new_n1091), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT61), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT119), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1082), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1083), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n1082), .A2(KEYINPUT119), .A3(new_n1083), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1084), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1095), .B1(new_n1096), .B2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n994), .A2(G2067), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1104), .B1(new_n1016), .B2(new_n744), .ZN(new_n1105));
  OR2_X1    g680(.A1(new_n1105), .A2(KEYINPUT120), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT120), .ZN(new_n1107));
  AOI211_X1 g682(.A(new_n1107), .B(new_n1104), .C1(new_n1016), .C2(new_n744), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT60), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1106), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1105), .A2(KEYINPUT120), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT60), .B1(new_n1112), .B2(new_n1108), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1111), .A2(new_n599), .A3(new_n1113), .ZN(new_n1114));
  OAI211_X1 g689(.A(KEYINPUT60), .B(new_n741), .C1(new_n1112), .C2(new_n1108), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1103), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  NOR3_X1   g691(.A1(new_n1112), .A2(new_n1108), .A3(new_n741), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1084), .ZN(new_n1118));
  OAI22_X1  g693(.A1(new_n1117), .A2(new_n1118), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1076), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n949), .B1(new_n1059), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(G1996), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n938), .A2(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(new_n1123), .B(KEYINPUT46), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n938), .B1(new_n939), .B2(new_n688), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n1126), .B(KEYINPUT47), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n938), .A2(new_n796), .A3(new_n587), .ZN(new_n1128));
  XNOR2_X1  g703(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n1128), .B(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1127), .B1(new_n947), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n943), .A2(new_n806), .A3(new_n803), .ZN(new_n1132));
  OR2_X1    g707(.A1(new_n763), .A2(G2067), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n944), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1121), .A2(new_n1135), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g711(.A1(G401), .A2(new_n457), .A3(G227), .ZN(new_n1138));
  NOR2_X1   g712(.A1(G229), .A2(new_n1138), .ZN(new_n1139));
  OAI211_X1 g713(.A(new_n1139), .B(new_n867), .C1(new_n927), .C2(new_n928), .ZN(G225));
  INV_X1    g714(.A(G225), .ZN(G308));
endmodule


