//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 0 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 1 1 0 0 0 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 1 0 1 0 0 1 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1272,
    new_n1273, new_n1275, new_n1276, new_n1277, new_n1278, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT65), .ZN(new_n214));
  AND2_X1   g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n207), .A2(KEYINPUT64), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT64), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G20), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n214), .A2(new_n215), .A3(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  INV_X1    g0023(.A(G87), .ZN(new_n224));
  INV_X1    g0024(.A(G250), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n209), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n212), .B(new_n220), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G226), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT67), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT68), .ZN(new_n244));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G1), .A2(G13), .ZN(new_n252));
  AND2_X1   g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G13), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n254), .A2(G1), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G20), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n206), .A2(G20), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(G77), .A3(new_n259), .ZN(new_n260));
  NOR3_X1   g0060(.A1(new_n254), .A2(new_n207), .A3(G1), .ZN(new_n261));
  INV_X1    g0061(.A(G77), .ZN(new_n262));
  AOI21_X1  g0062(.A(KEYINPUT72), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n261), .A2(KEYINPUT72), .A3(new_n262), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n251), .A2(new_n252), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT64), .B(G20), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G33), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT15), .B(G87), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT8), .B(G58), .ZN(new_n273));
  NOR2_X1   g0073(.A1(G20), .A2(G33), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  OAI22_X1  g0075(.A1(new_n262), .A2(new_n269), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n268), .B1(new_n272), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT71), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OAI211_X1 g0079(.A(KEYINPUT71), .B(new_n268), .C1(new_n272), .C2(new_n276), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n267), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT3), .B(G33), .ZN(new_n283));
  INV_X1    g0083(.A(G1698), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(G232), .A3(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT70), .B(G107), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n283), .A2(G1698), .ZN(new_n287));
  OAI221_X1 g0087(.A(new_n285), .B1(new_n283), .B2(new_n286), .C1(new_n287), .C2(new_n223), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n252), .B1(G33), .B2(G41), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G179), .ZN(new_n291));
  INV_X1    g0091(.A(G41), .ZN(new_n292));
  INV_X1    g0092(.A(G45), .ZN(new_n293));
  AOI21_X1  g0093(.A(G1), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(G33), .A2(G41), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n295), .A2(G1), .A3(G13), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n294), .A2(new_n296), .A3(G274), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n292), .A2(new_n293), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n206), .A2(new_n299), .B1(new_n215), .B2(new_n295), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n298), .B1(G244), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n290), .A2(new_n291), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n290), .A2(new_n301), .ZN(new_n303));
  INV_X1    g0103(.A(G169), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n282), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n303), .A2(G200), .ZN(new_n307));
  INV_X1    g0107(.A(G190), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n307), .B(new_n281), .C1(new_n308), .C2(new_n303), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n283), .A2(G222), .A3(new_n284), .ZN(new_n311));
  INV_X1    g0111(.A(G223), .ZN(new_n312));
  OAI221_X1 g0112(.A(new_n311), .B1(new_n262), .B2(new_n283), .C1(new_n287), .C2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(new_n289), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n298), .B1(G226), .B2(new_n300), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n291), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n261), .A2(new_n201), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n259), .A2(G50), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n318), .B1(new_n257), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT69), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI211_X1 g0122(.A(KEYINPUT69), .B(new_n318), .C1(new_n257), .C2(new_n319), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n325));
  INV_X1    g0125(.A(G150), .ZN(new_n326));
  OAI221_X1 g0126(.A(new_n325), .B1(new_n326), .B2(new_n275), .C1(new_n270), .C2(new_n273), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n268), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n317), .B(new_n329), .C1(G169), .C2(new_n316), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n329), .B(KEYINPUT9), .ZN(new_n331));
  INV_X1    g0131(.A(G200), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n332), .B1(new_n314), .B2(new_n315), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n333), .B1(G190), .B2(new_n316), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT10), .ZN(new_n335));
  AND3_X1   g0135(.A1(new_n331), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n335), .B1(new_n331), .B2(new_n334), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n310), .B(new_n330), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n261), .A2(new_n222), .ZN(new_n339));
  XNOR2_X1  g0139(.A(new_n339), .B(KEYINPUT12), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n258), .A2(G68), .A3(new_n259), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n274), .A2(G50), .B1(G20), .B2(new_n222), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(new_n270), .B2(new_n262), .ZN(new_n344));
  AND3_X1   g0144(.A1(new_n344), .A2(KEYINPUT11), .A3(new_n268), .ZN(new_n345));
  AOI21_X1  g0145(.A(KEYINPUT11), .B1(new_n344), .B2(new_n268), .ZN(new_n346));
  NOR3_X1   g0146(.A1(new_n342), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT14), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n283), .A2(G232), .A3(G1698), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n283), .A2(G226), .A3(new_n284), .ZN(new_n351));
  NAND2_X1  g0151(.A1(G33), .A2(G97), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n289), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n298), .B1(G238), .B2(new_n300), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT13), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n356), .B1(new_n354), .B2(new_n355), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n349), .B(G169), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n359), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n361), .A2(G179), .A3(new_n357), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n361), .A2(new_n357), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n349), .B1(new_n364), .B2(G169), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n348), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(G200), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n361), .A2(G190), .A3(new_n357), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n367), .A2(new_n347), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n273), .B1(new_n206), .B2(G20), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n258), .A2(new_n371), .B1(new_n261), .B2(new_n273), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  XNOR2_X1  g0173(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT7), .ZN(new_n375));
  AND2_X1   g0175(.A1(KEYINPUT3), .A2(G33), .ZN(new_n376));
  NOR2_X1   g0176(.A1(KEYINPUT3), .A2(G33), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n375), .B1(new_n378), .B2(new_n269), .ZN(new_n379));
  NOR4_X1   g0179(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT7), .A4(G20), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n379), .A2(new_n380), .A3(new_n222), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n202), .A2(new_n222), .ZN(new_n382));
  NOR2_X1   g0182(.A1(G58), .A2(G68), .ZN(new_n383));
  OAI21_X1  g0183(.A(G20), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n274), .A2(G159), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n374), .B1(new_n381), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT7), .B1(new_n283), .B2(G20), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n378), .A2(new_n269), .A3(new_n375), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(new_n389), .A3(G68), .ZN(new_n390));
  AND3_X1   g0190(.A1(new_n384), .A2(KEYINPUT16), .A3(new_n385), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n253), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n373), .B1(new_n387), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n312), .A2(new_n284), .ZN(new_n394));
  INV_X1    g0194(.A(G226), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(G1698), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n394), .B(new_n396), .C1(new_n376), .C2(new_n377), .ZN(new_n397));
  NAND2_X1  g0197(.A1(G33), .A2(G87), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n296), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n296), .A2(G232), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n297), .A2(new_n401), .ZN(new_n402));
  NOR3_X1   g0202(.A1(new_n399), .A2(new_n402), .A3(new_n291), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n397), .A2(new_n398), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n289), .ZN(new_n405));
  INV_X1    g0205(.A(G274), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n406), .B1(new_n215), .B2(new_n295), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n300), .A2(G232), .B1(new_n407), .B2(new_n294), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n403), .B1(new_n409), .B2(G169), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT18), .B1(new_n393), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n390), .A2(new_n391), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n268), .ZN(new_n413));
  INV_X1    g0213(.A(new_n374), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT7), .B1(new_n219), .B2(new_n283), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n378), .A2(new_n375), .A3(new_n207), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n415), .A2(G68), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n386), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n414), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n372), .B1(new_n413), .B2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT18), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n409), .A2(G169), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n409), .B2(new_n291), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n420), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n411), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n405), .A2(new_n308), .A3(new_n408), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n332), .B1(new_n399), .B2(new_n402), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n429), .B(new_n372), .C1(new_n413), .C2(new_n419), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT17), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n387), .A2(new_n392), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n433), .A2(KEYINPUT17), .A3(new_n372), .A4(new_n429), .ZN(new_n434));
  AND3_X1   g0234(.A1(new_n432), .A2(KEYINPUT74), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(KEYINPUT74), .B1(new_n432), .B2(new_n434), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n426), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n338), .A2(new_n370), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n286), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n415), .A2(new_n416), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT6), .ZN(new_n441));
  NOR3_X1   g0241(.A1(new_n441), .A2(G97), .A3(G107), .ZN(new_n442));
  INV_X1    g0242(.A(G97), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(KEYINPUT6), .ZN(new_n444));
  INV_X1    g0244(.A(G107), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n445), .A2(KEYINPUT76), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n445), .A2(KEYINPUT76), .ZN(new_n447));
  OAI22_X1  g0247(.A1(new_n442), .A2(new_n444), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  XNOR2_X1  g0248(.A(KEYINPUT76), .B(G107), .ZN(new_n449));
  INV_X1    g0249(.A(new_n444), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n443), .A2(new_n445), .A3(KEYINPUT6), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n448), .A2(new_n452), .A3(new_n219), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n274), .A2(G77), .ZN(new_n454));
  XNOR2_X1  g0254(.A(new_n454), .B(KEYINPUT75), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n440), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n268), .ZN(new_n457));
  INV_X1    g0257(.A(G33), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n253), .B(new_n256), .C1(G1), .C2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n459), .A2(new_n443), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n256), .A2(G97), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n457), .A2(new_n462), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n206), .B(G45), .C1(new_n292), .C2(KEYINPUT5), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT78), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT5), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G41), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT78), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n467), .A2(new_n468), .A3(new_n206), .A4(G45), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n466), .A2(G41), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n465), .A2(new_n469), .A3(new_n407), .A4(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT79), .ZN(new_n473));
  OAI211_X1 g0273(.A(G257), .B(new_n296), .C1(new_n464), .C2(new_n470), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n473), .B1(new_n472), .B2(new_n474), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT80), .ZN(new_n479));
  OAI211_X1 g0279(.A(G244), .B(new_n284), .C1(new_n376), .C2(new_n377), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT4), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT77), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n283), .A2(G244), .A3(new_n284), .A4(new_n482), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G33), .A2(G283), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n283), .A2(G250), .A3(G1698), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n484), .A2(new_n485), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n289), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n478), .A2(new_n479), .A3(G190), .A4(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n472), .A2(new_n474), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(KEYINPUT79), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n492), .A2(new_n489), .A3(new_n475), .ZN(new_n493));
  AOI21_X1  g0293(.A(KEYINPUT80), .B1(new_n493), .B2(G200), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n493), .A2(new_n308), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n463), .B(new_n490), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n493), .A2(new_n304), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n457), .A2(new_n462), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n492), .A2(new_n489), .A3(new_n291), .A4(new_n475), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n271), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(new_n256), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n459), .A2(new_n224), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n269), .A2(new_n283), .A3(G68), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n216), .A2(new_n218), .A3(G33), .A4(G97), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT19), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n216), .B(new_n218), .C1(new_n506), .C2(new_n352), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n445), .A2(KEYINPUT70), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT70), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G107), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n509), .A2(new_n511), .A3(new_n224), .A4(new_n443), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT81), .ZN(new_n513));
  AND3_X1   g0313(.A1(new_n508), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n513), .B1(new_n508), .B2(new_n512), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n504), .B(new_n507), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  AOI211_X1 g0316(.A(new_n502), .B(new_n503), .C1(new_n516), .C2(new_n268), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n225), .B1(new_n293), .B2(G1), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n206), .A2(new_n406), .A3(G45), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n296), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(G238), .B(new_n284), .C1(new_n376), .C2(new_n377), .ZN(new_n522));
  OAI211_X1 g0322(.A(G244), .B(G1698), .C1(new_n376), .C2(new_n377), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G116), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n521), .B1(new_n525), .B2(new_n289), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n526), .A2(new_n332), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n527), .B1(G190), .B2(new_n526), .ZN(new_n528));
  INV_X1    g0328(.A(new_n502), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n459), .A2(new_n271), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n507), .A2(new_n504), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n508), .A2(new_n512), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT81), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n508), .A2(new_n512), .A3(new_n513), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n532), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n529), .B(new_n531), .C1(new_n536), .C2(new_n253), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n526), .A2(G169), .ZN(new_n538));
  AOI211_X1 g0338(.A(G179), .B(new_n521), .C1(new_n525), .C2(new_n289), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n517), .A2(new_n528), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n496), .A2(new_n500), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n269), .A2(new_n283), .A3(G87), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT22), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT22), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n269), .A2(new_n283), .A3(new_n545), .A4(G87), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n524), .A2(G20), .ZN(new_n548));
  NOR2_X1   g0348(.A1(KEYINPUT23), .A2(G107), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n548), .B1(new_n219), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT82), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n509), .A2(new_n511), .A3(G20), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT23), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n551), .B1(new_n550), .B2(new_n553), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n547), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT24), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(KEYINPUT24), .B(new_n547), .C1(new_n554), .C2(new_n555), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n558), .A2(new_n268), .A3(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(G257), .B(G1698), .C1(new_n376), .C2(new_n377), .ZN(new_n561));
  OAI211_X1 g0361(.A(G250), .B(new_n284), .C1(new_n376), .C2(new_n377), .ZN(new_n562));
  XNOR2_X1  g0362(.A(KEYINPUT84), .B(G294), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n561), .B(new_n562), .C1(new_n458), .C2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n464), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n289), .B1(new_n565), .B2(new_n471), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n564), .A2(new_n289), .B1(new_n566), .B2(G264), .ZN(new_n567));
  AND3_X1   g0367(.A1(new_n567), .A2(G190), .A3(new_n472), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n332), .B1(new_n567), .B2(new_n472), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n261), .A2(new_n445), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT83), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n571), .A2(new_n572), .A3(KEYINPUT25), .ZN(new_n573));
  XOR2_X1   g0373(.A(KEYINPUT83), .B(KEYINPUT25), .Z(new_n574));
  OAI221_X1 g0374(.A(new_n573), .B1(new_n571), .B2(new_n574), .C1(new_n459), .C2(new_n445), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n560), .A2(new_n570), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n567), .A2(new_n472), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n304), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n567), .A2(new_n291), .A3(new_n472), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(new_n560), .B2(new_n576), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT21), .ZN(new_n583));
  INV_X1    g0383(.A(G116), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n261), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n459), .B2(new_n584), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n269), .B(new_n486), .C1(G33), .C2(new_n443), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n251), .A2(new_n252), .B1(G20), .B2(new_n584), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT20), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n587), .A2(KEYINPUT20), .A3(new_n588), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n586), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(G264), .B(G1698), .C1(new_n376), .C2(new_n377), .ZN(new_n594));
  OAI211_X1 g0394(.A(G257), .B(new_n284), .C1(new_n376), .C2(new_n377), .ZN(new_n595));
  OR2_X1    g0395(.A1(KEYINPUT3), .A2(G33), .ZN(new_n596));
  NAND2_X1  g0396(.A1(KEYINPUT3), .A2(G33), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n596), .A2(G303), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n594), .A2(new_n595), .A3(new_n598), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n599), .A2(new_n289), .ZN(new_n600));
  OAI211_X1 g0400(.A(G270), .B(new_n296), .C1(new_n464), .C2(new_n470), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n472), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(G169), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n583), .B1(new_n593), .B2(new_n603), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n472), .A2(new_n601), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n599), .A2(new_n289), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(G190), .A3(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n600), .A2(new_n602), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n593), .B(new_n607), .C1(new_n608), .C2(new_n332), .ZN(new_n609));
  NOR3_X1   g0409(.A1(new_n600), .A2(new_n602), .A3(new_n291), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n458), .A2(G1), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n257), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(G116), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n587), .A2(KEYINPUT20), .A3(new_n588), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT20), .B1(new_n587), .B2(new_n588), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n613), .B(new_n585), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n304), .B1(new_n605), .B2(new_n606), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n618), .A2(new_n616), .A3(KEYINPUT21), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n604), .A2(new_n609), .A3(new_n617), .A4(new_n619), .ZN(new_n620));
  NOR3_X1   g0420(.A1(new_n577), .A2(new_n582), .A3(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n438), .A2(new_n542), .A3(new_n621), .ZN(G372));
  AOI211_X1 g0422(.A(new_n502), .B(new_n530), .C1(new_n516), .C2(new_n268), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n526), .A2(new_n291), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n624), .B1(G169), .B2(new_n526), .ZN(new_n625));
  INV_X1    g0425(.A(new_n503), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n529), .B(new_n626), .C1(new_n536), .C2(new_n253), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n526), .A2(G190), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n628), .B1(new_n332), .B2(new_n526), .ZN(new_n629));
  OAI22_X1  g0429(.A1(new_n623), .A2(new_n625), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT26), .ZN(new_n631));
  NOR3_X1   g0431(.A1(new_n630), .A2(new_n500), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n498), .A2(new_n499), .ZN(new_n633));
  AOI21_X1  g0433(.A(G169), .B1(new_n478), .B2(new_n489), .ZN(new_n634));
  OAI21_X1  g0434(.A(KEYINPUT85), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT85), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n497), .A2(new_n636), .A3(new_n498), .A4(new_n499), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n635), .A2(new_n541), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n632), .B1(new_n631), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n537), .A2(new_n540), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n253), .B1(new_n556), .B2(new_n557), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n575), .B1(new_n641), .B2(new_n559), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n570), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n604), .A2(new_n617), .A3(new_n619), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n643), .B1(new_n582), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n493), .A2(G200), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n492), .A2(new_n489), .A3(new_n475), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n646), .A2(new_n479), .B1(new_n647), .B2(G190), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n490), .A2(new_n463), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n541), .B(new_n500), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n640), .B1(new_n645), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n438), .B1(new_n639), .B2(new_n651), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n282), .A2(new_n302), .A3(new_n305), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n369), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n366), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT74), .ZN(new_n656));
  INV_X1    g0456(.A(new_n434), .ZN(new_n657));
  AOI21_X1  g0457(.A(KEYINPUT17), .B1(new_n393), .B2(new_n429), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n432), .A2(KEYINPUT74), .A3(new_n434), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n425), .B1(new_n655), .B2(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n662), .A2(KEYINPUT86), .ZN(new_n663));
  OAI22_X1  g0463(.A1(new_n662), .A2(KEYINPUT86), .B1(new_n337), .B2(new_n336), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n652), .B(new_n330), .C1(new_n663), .C2(new_n664), .ZN(G369));
  INV_X1    g0465(.A(KEYINPUT88), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n269), .A2(new_n255), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(KEYINPUT87), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT87), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n269), .A2(new_n669), .A3(new_n255), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT27), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n668), .A2(new_n673), .A3(new_n670), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n672), .A2(G213), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(G343), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n666), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NOR3_X1   g0478(.A1(new_n675), .A2(new_n666), .A3(new_n676), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(new_n593), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n644), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n620), .B2(new_n681), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G330), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n549), .ZN(new_n686));
  OAI22_X1  g0486(.A1(new_n269), .A2(new_n686), .B1(G20), .B2(new_n524), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT23), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n688), .B1(new_n286), .B2(G20), .ZN(new_n689));
  OAI21_X1  g0489(.A(KEYINPUT82), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n550), .A2(new_n553), .A3(new_n551), .ZN(new_n691));
  AOI22_X1  g0491(.A1(new_n690), .A2(new_n691), .B1(new_n544), .B2(new_n546), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n268), .B1(new_n692), .B2(KEYINPUT24), .ZN(new_n693));
  INV_X1    g0493(.A(new_n559), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n576), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n581), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n643), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n680), .A2(new_n642), .ZN(new_n699));
  OAI22_X1  g0499(.A1(new_n698), .A2(new_n699), .B1(new_n697), .B2(new_n680), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n685), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n680), .A2(new_n644), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n703), .B1(new_n582), .B2(new_n680), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n701), .A2(new_n704), .ZN(G399));
  INV_X1    g0505(.A(new_n210), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(G41), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(new_n206), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n512), .A2(G116), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n708), .A2(new_n709), .B1(new_n214), .B2(new_n707), .ZN(new_n710));
  XOR2_X1   g0510(.A(new_n710), .B(KEYINPUT28), .Z(new_n711));
  OAI21_X1  g0511(.A(new_n680), .B1(new_n651), .B2(new_n639), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT29), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n635), .A2(KEYINPUT26), .A3(new_n541), .A4(new_n637), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n631), .B1(new_n630), .B2(new_n500), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  XOR2_X1   g0518(.A(new_n640), .B(KEYINPUT90), .Z(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n645), .B2(new_n650), .ZN(new_n720));
  OAI211_X1 g0520(.A(KEYINPUT29), .B(new_n680), .C1(new_n718), .C2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n714), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(G330), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT30), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n608), .A2(G179), .A3(new_n526), .A4(new_n567), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n724), .B1(new_n725), .B2(new_n493), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n567), .A2(new_n526), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n647), .A2(new_n610), .A3(KEYINPUT30), .A4(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT89), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n525), .A2(new_n289), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(new_n520), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n729), .A2(new_n731), .B1(new_n567), .B2(new_n472), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n526), .A2(KEYINPUT89), .ZN(new_n733));
  AOI21_X1  g0533(.A(G179), .B1(new_n605), .B2(new_n606), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n732), .A2(new_n733), .A3(new_n493), .A4(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n726), .A2(new_n728), .A3(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n679), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n677), .ZN(new_n738));
  AND3_X1   g0538(.A1(new_n736), .A2(KEYINPUT31), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(KEYINPUT31), .B1(new_n736), .B2(new_n738), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n621), .A2(new_n542), .A3(new_n680), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n723), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n722), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n711), .B1(new_n746), .B2(G1), .ZN(new_n747));
  XOR2_X1   g0547(.A(new_n747), .B(KEYINPUT91), .Z(G364));
  NOR3_X1   g0548(.A1(new_n219), .A2(new_n254), .A3(new_n293), .ZN(new_n749));
  OR2_X1    g0549(.A1(new_n749), .A2(KEYINPUT92), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(KEYINPUT92), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n708), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n706), .A2(new_n378), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G355), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n757), .B1(G116), .B2(new_n210), .ZN(new_n758));
  OR2_X1    g0558(.A1(new_n246), .A2(new_n293), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n706), .A2(new_n283), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n761), .B1(new_n214), .B2(new_n293), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n758), .B1(new_n759), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G13), .A2(G33), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(G20), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n252), .B1(G20), .B2(new_n304), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n755), .B1(new_n763), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n219), .A2(new_n308), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n772), .A2(KEYINPUT93), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n332), .A2(G179), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n772), .A2(KEYINPUT93), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n773), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(G179), .A2(G200), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n773), .A2(new_n775), .A3(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI22_X1  g0580(.A1(G283), .A2(new_n777), .B1(new_n780), .B2(G329), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT96), .Z(new_n782));
  NAND3_X1  g0582(.A1(new_n774), .A2(G20), .A3(G190), .ZN(new_n783));
  INV_X1    g0583(.A(G303), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n378), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n771), .A2(new_n291), .A3(new_n332), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  XOR2_X1   g0587(.A(KEYINPUT33), .B(G317), .Z(new_n788));
  AOI21_X1  g0588(.A(new_n269), .B1(G190), .B2(new_n778), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n787), .A2(new_n788), .B1(new_n563), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n269), .A2(new_n291), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G190), .A2(G200), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n785), .B(new_n790), .C1(G311), .C2(new_n793), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n791), .A2(G190), .A3(new_n332), .ZN(new_n795));
  INV_X1    g0595(.A(G322), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n791), .A2(G190), .A3(G200), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n797), .B1(G326), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n782), .A2(new_n794), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n777), .A2(G107), .ZN(new_n802));
  OAI211_X1 g0602(.A(new_n802), .B(new_n283), .C1(new_n224), .C2(new_n783), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT95), .ZN(new_n804));
  XOR2_X1   g0604(.A(KEYINPUT94), .B(G159), .Z(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n780), .A2(new_n806), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n807), .A2(KEYINPUT32), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(KEYINPUT32), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n201), .A2(new_n798), .B1(new_n795), .B2(new_n202), .ZN(new_n810));
  INV_X1    g0610(.A(new_n793), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n811), .A2(new_n262), .B1(new_n789), .B2(new_n443), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n810), .B(new_n812), .C1(G68), .C2(new_n786), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n808), .A2(new_n809), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n801), .B1(new_n804), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n770), .B1(new_n815), .B2(new_n767), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT97), .Z(new_n817));
  INV_X1    g0617(.A(new_n766), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n683), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n685), .A2(new_n755), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(G330), .B2(new_n683), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(G396));
  NOR2_X1   g0623(.A1(new_n738), .A2(new_n306), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n282), .B1(new_n678), .B2(new_n679), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n653), .B1(new_n825), .B2(new_n309), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n712), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n826), .A2(new_n824), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n680), .B(new_n828), .C1(new_n651), .C2(new_n639), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n755), .B1(new_n830), .B2(new_n744), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n744), .B2(new_n830), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n767), .A2(new_n764), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n754), .B1(new_n262), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n767), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n777), .A2(G87), .ZN(new_n836));
  INV_X1    g0636(.A(G311), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n836), .B1(new_n837), .B2(new_n779), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n378), .B1(new_n445), .B2(new_n783), .C1(new_n789), .C2(new_n443), .ZN(new_n839));
  INV_X1    g0639(.A(G283), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n584), .A2(new_n811), .B1(new_n787), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(G294), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n842), .A2(new_n795), .B1(new_n798), .B2(new_n784), .ZN(new_n843));
  NOR4_X1   g0643(.A1(new_n838), .A2(new_n839), .A3(new_n841), .A4(new_n843), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n793), .A2(new_n806), .B1(new_n786), .B2(G150), .ZN(new_n845));
  INV_X1    g0645(.A(G137), .ZN(new_n846));
  INV_X1    g0646(.A(G143), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n845), .B1(new_n846), .B2(new_n798), .C1(new_n847), .C2(new_n795), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT34), .ZN(new_n849));
  OR2_X1    g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n777), .A2(G68), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n283), .B1(new_n783), .B2(new_n201), .ZN(new_n852));
  INV_X1    g0652(.A(new_n789), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n852), .B1(new_n853), .B2(G58), .ZN(new_n854));
  INV_X1    g0654(.A(G132), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n851), .B(new_n854), .C1(new_n855), .C2(new_n779), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(new_n849), .B2(new_n848), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n844), .B1(new_n850), .B2(new_n857), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n834), .B1(new_n828), .B2(new_n765), .C1(new_n835), .C2(new_n858), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n832), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(G384));
  NOR3_X1   g0661(.A1(new_n269), .A2(new_n584), .A3(new_n252), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n448), .A2(new_n452), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(KEYINPUT98), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT35), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n862), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(new_n866), .B2(new_n865), .ZN(new_n868));
  XNOR2_X1  g0668(.A(KEYINPUT99), .B(KEYINPUT36), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n868), .B(new_n869), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n214), .B(G77), .C1(new_n202), .C2(new_n222), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n201), .A2(G68), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n206), .B(G13), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n741), .A2(new_n742), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n680), .A2(new_n347), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n370), .A2(new_n876), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n366), .B(new_n369), .C1(new_n347), .C2(new_n680), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n875), .A2(new_n879), .A3(new_n828), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT38), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n414), .B1(new_n390), .B2(new_n418), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n373), .B1(new_n884), .B2(new_n392), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n430), .B1(new_n885), .B2(new_n675), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n885), .A2(new_n410), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT37), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n420), .A2(new_n423), .ZN(new_n889));
  INV_X1    g0689(.A(new_n675), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n420), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT37), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n889), .A2(new_n891), .A3(new_n892), .A4(new_n430), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n882), .B1(new_n888), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n425), .B1(new_n659), .B2(new_n660), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n372), .B1(new_n413), .B2(new_n883), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n890), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n894), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT101), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n897), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n437), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n902), .A2(KEYINPUT101), .A3(new_n894), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n889), .A2(new_n891), .A3(new_n430), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT37), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n893), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n432), .A2(new_n434), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n420), .B(new_n890), .C1(new_n425), .C2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g0709(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n900), .A2(new_n903), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n881), .A2(new_n912), .A3(KEYINPUT40), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT40), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n888), .A2(new_n893), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT38), .B1(new_n902), .B2(new_n915), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n890), .A2(new_n896), .B1(new_n393), .B2(new_n429), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n896), .A2(new_n423), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n892), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n893), .ZN(new_n920));
  OAI21_X1  g0720(.A(KEYINPUT38), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(new_n437), .B2(new_n901), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n916), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n914), .B1(new_n923), .B2(new_n880), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n913), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT104), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n438), .A2(new_n875), .ZN(new_n927));
  OAI21_X1  g0727(.A(G330), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(new_n927), .B2(new_n926), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n364), .A2(G169), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(KEYINPUT14), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n931), .A2(new_n362), .A3(new_n360), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n932), .A2(new_n348), .A3(new_n680), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(KEYINPUT39), .B1(new_n916), .B2(new_n922), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT102), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT39), .B1(new_n909), .B2(new_n910), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n900), .A2(new_n903), .A3(new_n937), .ZN(new_n938));
  AND3_X1   g0738(.A1(new_n935), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n936), .B1(new_n935), .B2(new_n938), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n934), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n824), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n829), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n879), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n944), .A2(new_n923), .B1(new_n426), .B2(new_n890), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n941), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n330), .B1(new_n664), .B2(new_n663), .ZN(new_n948));
  INV_X1    g0748(.A(new_n640), .ZN(new_n949));
  AND3_X1   g0749(.A1(new_n604), .A2(new_n617), .A3(new_n619), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n697), .A2(new_n950), .B1(new_n642), .B2(new_n570), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n949), .B1(new_n542), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n638), .A2(new_n631), .ZN(new_n953));
  INV_X1    g0753(.A(new_n632), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n738), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n721), .B(new_n438), .C1(new_n956), .C2(KEYINPUT29), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(KEYINPUT103), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT103), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n714), .A2(new_n959), .A3(new_n438), .A4(new_n721), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n948), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n947), .B(new_n961), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n929), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(G1), .B1(new_n219), .B2(new_n254), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n929), .B2(new_n962), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n874), .B1(new_n963), .B2(new_n965), .ZN(G367));
  NOR2_X1   g0766(.A1(new_n752), .A2(new_n206), .ZN(new_n967));
  INV_X1    g0767(.A(new_n702), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n700), .A2(new_n968), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n969), .A2(KEYINPUT106), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n969), .A2(KEYINPUT106), .ZN(new_n971));
  NOR3_X1   g0771(.A1(new_n970), .A2(new_n971), .A3(new_n703), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n684), .B(KEYINPUT107), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n972), .B1(KEYINPUT107), .B2(new_n685), .ZN(new_n975));
  AND3_X1   g0775(.A1(new_n974), .A2(new_n746), .A3(new_n975), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n496), .B(new_n500), .C1(new_n680), .C2(new_n463), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n680), .A2(new_n500), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n704), .A2(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT45), .Z(new_n981));
  NOR2_X1   g0781(.A1(new_n704), .A2(new_n979), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT44), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n984), .A2(new_n685), .A3(new_n700), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n976), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n981), .A2(new_n701), .A3(new_n983), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT108), .Z(new_n988));
  AOI21_X1  g0788(.A(new_n745), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n707), .B(KEYINPUT41), .Z(new_n990));
  OAI21_X1  g0790(.A(new_n967), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n500), .B1(new_n977), .B2(new_n697), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT105), .ZN(new_n993));
  AND2_X1   g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n992), .A2(new_n993), .ZN(new_n995));
  NOR3_X1   g0795(.A1(new_n994), .A2(new_n995), .A3(new_n738), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n979), .A2(new_n703), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT42), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT43), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n738), .A2(new_n627), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(new_n630), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n996), .A2(new_n998), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n999), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1002), .B(new_n1003), .Z(new_n1004));
  AOI21_X1  g0804(.A(new_n701), .B1(new_n977), .B2(new_n978), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n991), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n789), .A2(new_n222), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n783), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n378), .B(new_n1008), .C1(G58), .C2(new_n1009), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1010), .B1(new_n201), .B2(new_n811), .C1(new_n787), .C2(new_n805), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n777), .A2(G77), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n846), .B2(new_n779), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n847), .A2(new_n798), .B1(new_n795), .B2(new_n326), .ZN(new_n1014));
  NOR3_X1   g0814(.A1(new_n1011), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT109), .Z(new_n1016));
  AOI21_X1  g0816(.A(KEYINPUT46), .B1(new_n1009), .B2(G116), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1017), .A2(new_n283), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1009), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1018), .B(new_n1019), .C1(new_n784), .C2(new_n795), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(G311), .B2(new_n799), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n840), .A2(new_n811), .B1(new_n787), .B2(new_n563), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(new_n439), .B2(new_n853), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n780), .A2(G317), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n777), .A2(G97), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1021), .A2(new_n1023), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1016), .A2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT47), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n767), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1001), .A2(new_n766), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n241), .A2(new_n760), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n769), .B1(new_n706), .B2(new_n501), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n754), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1029), .A2(new_n1030), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1007), .A2(new_n1034), .ZN(G387));
  AOI21_X1  g0835(.A(new_n761), .B1(new_n237), .B2(G45), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n709), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1036), .B1(new_n1037), .B2(new_n756), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n273), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n201), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT50), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n293), .B1(new_n222), .B2(new_n262), .ZN(new_n1042));
  NOR3_X1   g0842(.A1(new_n1041), .A2(new_n1037), .A3(new_n1042), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n1038), .A2(new_n1043), .B1(G107), .B2(new_n210), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n754), .B1(new_n1044), .B2(new_n768), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n700), .B2(new_n818), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n283), .B1(new_n783), .B2(new_n262), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n787), .A2(new_n273), .B1(new_n789), .B2(new_n271), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n1047), .B(new_n1048), .C1(G68), .C2(new_n793), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n795), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G50), .A2(new_n1050), .B1(new_n799), .B2(G159), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n780), .A2(G150), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1049), .A2(new_n1025), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n283), .B1(new_n780), .B2(G326), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n853), .A2(G283), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(G303), .A2(new_n793), .B1(new_n786), .B2(G311), .ZN(new_n1056));
  INV_X1    g0856(.A(G317), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1056), .B1(new_n1057), .B2(new_n795), .C1(new_n796), .C2(new_n798), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT110), .Z(new_n1059));
  OAI221_X1 g0859(.A(new_n1055), .B1(new_n563), .B2(new_n783), .C1(new_n1059), .C2(KEYINPUT48), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(KEYINPUT48), .B2(new_n1059), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT111), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT49), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1054), .B1(new_n584), .B2(new_n776), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1064));
  AND2_X1   g0864(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1053), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1046), .B1(new_n1066), .B2(new_n767), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n974), .A2(new_n975), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n967), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n707), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n976), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n746), .B2(new_n1068), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1070), .A2(new_n1073), .ZN(G393));
  XOR2_X1   g0874(.A(new_n985), .B(KEYINPUT112), .Z(new_n1075));
  NAND3_X1  g0875(.A1(new_n1075), .A2(new_n988), .A3(new_n1069), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n768), .B1(new_n443), .B2(new_n210), .C1(new_n761), .C2(new_n249), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n755), .A2(new_n1077), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n779), .A2(new_n847), .B1(new_n222), .B2(new_n783), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT114), .ZN(new_n1080));
  INV_X1    g0880(.A(G159), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n326), .A2(new_n798), .B1(new_n795), .B2(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT51), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n378), .B1(new_n793), .B2(new_n1039), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n789), .A2(new_n262), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(G50), .B2(new_n786), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1083), .A2(new_n836), .A3(new_n1084), .A4(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n780), .A2(G322), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n378), .B1(new_n783), .B2(new_n840), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n793), .B2(G294), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(G303), .A2(new_n786), .B1(new_n853), .B2(G116), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n802), .A2(new_n1088), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n837), .A2(new_n795), .B1(new_n798), .B2(new_n1057), .ZN(new_n1093));
  XOR2_X1   g0893(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n1094));
  XNOR2_X1  g0894(.A(new_n1093), .B(new_n1094), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n1080), .A2(new_n1087), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1078), .B1(new_n1096), .B2(new_n767), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT116), .Z(new_n1098));
  NOR2_X1   g0898(.A1(new_n979), .A2(new_n818), .ZN(new_n1099));
  OR2_X1    g0899(.A1(new_n1099), .A2(KEYINPUT113), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(KEYINPUT113), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1098), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n976), .B1(new_n1075), .B2(new_n988), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n986), .A2(new_n988), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n707), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1076), .B(new_n1102), .C1(new_n1103), .C2(new_n1105), .ZN(G390));
  NAND2_X1  g0906(.A1(new_n736), .A2(new_n738), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT31), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n736), .A2(KEYINPUT31), .A3(new_n738), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AND4_X1   g0911(.A1(new_n604), .A2(new_n609), .A3(new_n617), .A4(new_n619), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1112), .A2(new_n643), .A3(new_n697), .ZN(new_n1113));
  NOR3_X1   g0913(.A1(new_n1113), .A2(new_n650), .A3(new_n738), .ZN(new_n1114));
  OAI211_X1 g0914(.A(G330), .B(new_n828), .C1(new_n1111), .C2(new_n1114), .ZN(new_n1115));
  AND2_X1   g0915(.A1(new_n877), .A2(new_n878), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n934), .B1(new_n943), .B2(new_n879), .ZN(new_n1118));
  NOR3_X1   g0918(.A1(new_n939), .A2(new_n940), .A3(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n640), .B(KEYINPUT90), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(new_n542), .B2(new_n951), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n738), .B1(new_n1121), .B2(new_n717), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n826), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n824), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n933), .B(new_n912), .C1(new_n1124), .C2(new_n1116), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1117), .B1(new_n1119), .B2(new_n1126), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n900), .A2(new_n903), .A3(new_n937), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT39), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n897), .B1(new_n661), .B2(new_n426), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n915), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n882), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1129), .B1(new_n1132), .B2(new_n898), .ZN(new_n1133));
  OAI21_X1  g0933(.A(KEYINPUT102), .B1(new_n1128), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n944), .A2(new_n933), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n935), .A2(new_n938), .A3(new_n936), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT117), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n743), .A2(KEYINPUT117), .A3(new_n828), .A4(new_n879), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1137), .A2(new_n1125), .A3(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1127), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1139), .A2(new_n1124), .A3(new_n1140), .A4(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n879), .B1(new_n743), .B2(new_n828), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n943), .B1(new_n1117), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n743), .A2(new_n438), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n1148), .A2(new_n961), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1071), .B1(new_n1143), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1127), .A2(new_n1150), .A3(new_n1142), .ZN(new_n1153));
  AND2_X1   g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1134), .A2(new_n764), .A3(new_n1136), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n789), .A2(new_n1081), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(KEYINPUT54), .B(G143), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n811), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT53), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n783), .B2(new_n326), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1009), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n1156), .B(new_n1158), .C1(new_n1160), .C2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(G125), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n1162), .B1(new_n201), .B2(new_n776), .C1(new_n1163), .C2(new_n779), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n378), .B1(new_n786), .B2(G137), .ZN(new_n1165));
  INV_X1    g0965(.A(G128), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n1165), .B1(new_n1166), .B2(new_n798), .C1(new_n855), .C2(new_n795), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(G97), .A2(new_n793), .B1(new_n786), .B2(new_n439), .ZN(new_n1168));
  XOR2_X1   g0968(.A(new_n1168), .B(KEYINPUT118), .Z(new_n1169));
  OAI211_X1 g0969(.A(new_n1169), .B(new_n851), .C1(new_n842), .C2(new_n779), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n283), .B(new_n1085), .C1(G87), .C2(new_n1009), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1171), .B1(new_n584), .B2(new_n795), .C1(new_n840), .C2(new_n798), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n1164), .A2(new_n1167), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n767), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n754), .B1(new_n273), .B2(new_n833), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1155), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n1143), .B2(new_n967), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1154), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(G378));
  INV_X1    g0979(.A(KEYINPUT122), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n890), .A2(new_n329), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n336), .A2(new_n337), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n330), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1182), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NOR3_X1   g0986(.A1(new_n1183), .A2(new_n1184), .A3(new_n1182), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1188), .B(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT121), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n913), .A2(new_n924), .A3(G330), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n941), .A2(new_n946), .A3(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1194), .B1(new_n941), .B2(new_n946), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1193), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1194), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n933), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1198), .B1(new_n1199), .B2(new_n945), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1193), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n941), .A2(new_n946), .A3(new_n1194), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n961), .A2(new_n1149), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1197), .A2(new_n1203), .B1(new_n1153), .B2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1180), .B1(new_n1206), .B2(KEYINPUT57), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1071), .B1(new_n1206), .B2(KEYINPUT57), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT57), .ZN(new_n1209));
  AND3_X1   g1009(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1201), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  AND3_X1   g1012(.A1(new_n1137), .A2(new_n1125), .A3(new_n1141), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1117), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n1137), .B2(new_n1125), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1213), .A2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1204), .B1(new_n1216), .B2(new_n1150), .ZN(new_n1217));
  OAI211_X1 g1017(.A(KEYINPUT122), .B(new_n1209), .C1(new_n1212), .C2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1207), .A2(new_n1208), .A3(new_n1218), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1212), .A2(new_n967), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1191), .A2(new_n764), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n378), .A2(new_n292), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n1222), .B(new_n1008), .C1(G77), .C2(new_n1009), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1223), .B1(new_n443), .B2(new_n787), .C1(new_n271), .C2(new_n811), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n777), .A2(G58), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n840), .B2(new_n779), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n445), .A2(new_n795), .B1(new_n798), .B2(new_n584), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(new_n1224), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  XOR2_X1   g1028(.A(new_n1228), .B(KEYINPUT58), .Z(new_n1229));
  OAI211_X1 g1029(.A(new_n1222), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n846), .A2(new_n811), .B1(new_n787), .B2(new_n855), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n789), .A2(new_n326), .B1(new_n783), .B2(new_n1157), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n1163), .A2(new_n798), .B1(new_n795), .B2(new_n1166), .ZN(new_n1233));
  NOR3_X1   g1033(.A1(new_n1231), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1235), .A2(KEYINPUT59), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n458), .B(new_n292), .C1(new_n776), .C2(new_n805), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(G124), .B2(new_n780), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT59), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1238), .B1(new_n1239), .B2(new_n1234), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1229), .B(new_n1230), .C1(new_n1236), .C2(new_n1240), .ZN(new_n1241));
  XOR2_X1   g1041(.A(new_n1241), .B(KEYINPUT119), .Z(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n767), .ZN(new_n1243));
  XOR2_X1   g1043(.A(new_n1243), .B(KEYINPUT120), .Z(new_n1244));
  INV_X1    g1044(.A(new_n833), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n755), .B1(G50), .B2(new_n1245), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1244), .A2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1220), .B1(new_n1221), .B2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1219), .A2(new_n1248), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1249), .B(KEYINPUT123), .ZN(G375));
  NAND2_X1  g1050(.A1(new_n1116), .A2(new_n764), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n378), .B1(new_n783), .B2(new_n443), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n286), .A2(new_n811), .B1(new_n787), .B2(new_n584), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n1252), .B(new_n1253), .C1(new_n501), .C2(new_n853), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(G283), .A2(new_n1050), .B1(new_n799), .B2(G294), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n780), .A2(G303), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1254), .A2(new_n1012), .A3(new_n1255), .A4(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n283), .B1(new_n783), .B2(new_n1081), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n787), .A2(new_n1157), .B1(new_n789), .B2(new_n201), .ZN(new_n1259));
  AOI211_X1 g1059(.A(new_n1258), .B(new_n1259), .C1(G150), .C2(new_n793), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(G132), .A2(new_n799), .B1(new_n1050), .B2(G137), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n780), .A2(G128), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1260), .A2(new_n1225), .A3(new_n1261), .A4(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n835), .B1(new_n1257), .B2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n755), .B1(G68), .B2(new_n1245), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1265), .B(KEYINPUT124), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n1148), .A2(new_n1069), .B1(new_n1251), .B2(new_n1267), .ZN(new_n1268));
  OR2_X1    g1068(.A1(new_n1150), .A2(new_n990), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1205), .A2(new_n1148), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1268), .B1(new_n1269), .B2(new_n1270), .ZN(G381));
  NAND4_X1  g1071(.A1(new_n1070), .A2(new_n1073), .A3(new_n822), .A4(new_n860), .ZN(new_n1272));
  OR4_X1    g1072(.A1(G387), .A2(new_n1272), .A3(G390), .A4(G381), .ZN(new_n1273));
  OR3_X1    g1073(.A1(G375), .A2(new_n1273), .A3(G378), .ZN(G407));
  NOR2_X1   g1074(.A1(G375), .A2(G378), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n676), .A2(G213), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1278), .A2(G407), .A3(G213), .ZN(G409));
  INV_X1    g1079(.A(new_n1034), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1280), .B1(new_n991), .B2(new_n1006), .ZN(new_n1281));
  OR2_X1    g1081(.A1(new_n1281), .A2(G390), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(G390), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT126), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1285), .B1(new_n1281), .B2(G390), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(G393), .B(G396), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1284), .A2(new_n1288), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1282), .A2(new_n1283), .A3(KEYINPUT126), .A4(new_n1287), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1219), .A2(G378), .A3(new_n1248), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1247), .A2(new_n1221), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1293), .B1(new_n967), .B2(new_n1212), .ZN(new_n1294));
  NOR3_X1   g1094(.A1(new_n1212), .A2(new_n1217), .A3(new_n990), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1178), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1292), .A2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1276), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1270), .B1(new_n1151), .B2(KEYINPUT60), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1204), .A2(KEYINPUT60), .A3(new_n1147), .A4(new_n1145), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n707), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1268), .B1(new_n1299), .B2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n860), .ZN(new_n1303));
  OAI211_X1 g1103(.A(G384), .B(new_n1268), .C1(new_n1299), .C2(new_n1301), .ZN(new_n1304));
  OR2_X1    g1104(.A1(new_n1276), .A2(KEYINPUT125), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1303), .A2(new_n1304), .A3(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1306), .A2(G2897), .A3(new_n1277), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1277), .A2(G2897), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1303), .A2(new_n1304), .A3(new_n1308), .A4(new_n1305), .ZN(new_n1309));
  AND2_X1   g1109(.A1(new_n1307), .A2(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(KEYINPUT61), .B1(new_n1298), .B2(new_n1310), .ZN(new_n1311));
  AND2_X1   g1111(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1297), .A2(new_n1276), .A3(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT63), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1277), .B1(new_n1292), .B2(new_n1296), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1316), .A2(KEYINPUT63), .A3(new_n1312), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1291), .A2(new_n1311), .A3(new_n1315), .A4(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1291), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT61), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1307), .A2(new_n1309), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1320), .B1(new_n1316), .B2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT62), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1313), .A2(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1316), .A2(KEYINPUT62), .A3(new_n1312), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1322), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1319), .B1(new_n1326), .B2(KEYINPUT127), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1325), .ZN(new_n1328));
  AOI21_X1  g1128(.A(KEYINPUT62), .B1(new_n1316), .B2(new_n1312), .ZN(new_n1329));
  OAI211_X1 g1129(.A(KEYINPUT127), .B(new_n1311), .C1(new_n1328), .C2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1330), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1318), .B1(new_n1327), .B2(new_n1331), .ZN(G405));
  INV_X1    g1132(.A(new_n1312), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1290), .ZN(new_n1334));
  AOI22_X1  g1134(.A1(new_n1282), .A2(new_n1283), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1333), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1289), .A2(new_n1312), .A3(new_n1290), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1178), .B1(new_n1219), .B2(new_n1248), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1275), .A2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1338), .A2(new_n1340), .ZN(new_n1341));
  OAI211_X1 g1141(.A(new_n1336), .B(new_n1337), .C1(new_n1275), .C2(new_n1339), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1341), .A2(new_n1342), .ZN(G402));
endmodule


