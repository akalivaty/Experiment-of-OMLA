//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 1 0 0 0 1 0 1 0 1 1 1 1 0 0 0 0 1 1 1 1 0 1 0 0 1 0 1 1 0 0 1 1 1 1 0 0 1 0 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n796, new_n797, new_n798, new_n799,
    new_n801, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n979, new_n980, new_n981, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1010, new_n1011, new_n1012;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT90), .B(G197gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(KEYINPUT11), .B(G169gat), .Z(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT12), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G43gat), .B(G50gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT15), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT91), .B(G50gat), .ZN(new_n212));
  INV_X1    g011(.A(G43gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI21_X1  g013(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(KEYINPUT14), .B(G29gat), .ZN(new_n217));
  INV_X1    g016(.A(G36gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G29gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n220), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n211), .B1(new_n216), .B2(new_n222), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n210), .B1(new_n219), .B2(new_n221), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT17), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G15gat), .B(G22gat), .ZN(new_n226));
  INV_X1    g025(.A(G1gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT16), .ZN(new_n228));
  AND2_X1   g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n226), .A2(G1gat), .ZN(new_n230));
  NOR3_X1   g029(.A1(new_n229), .A2(new_n230), .A3(G8gat), .ZN(new_n231));
  INV_X1    g030(.A(G8gat), .ZN(new_n232));
  XOR2_X1   g031(.A(G15gat), .B(G22gat), .Z(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(new_n227), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n226), .A2(new_n228), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n232), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n231), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT17), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n211), .ZN(new_n239));
  AOI22_X1  g038(.A1(new_n219), .A2(new_n221), .B1(new_n214), .B2(new_n215), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n238), .B(new_n239), .C1(new_n240), .C2(new_n211), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n237), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT92), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT93), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n239), .B1(new_n240), .B2(new_n211), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n245), .B1(new_n246), .B2(new_n237), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n223), .A2(new_n224), .ZN(new_n248));
  OAI21_X1  g047(.A(G8gat), .B1(new_n229), .B2(new_n230), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n234), .A2(new_n232), .A3(new_n235), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n248), .A2(KEYINPUT93), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n247), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(G229gat), .A2(G233gat), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n225), .A2(KEYINPUT92), .A3(new_n237), .A4(new_n241), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n244), .A2(new_n253), .A3(new_n254), .A4(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT18), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n246), .A2(new_n237), .ZN(new_n260));
  NOR3_X1   g059(.A1(new_n246), .A2(new_n237), .A3(new_n245), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT93), .B1(new_n248), .B2(new_n251), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT94), .B(KEYINPUT13), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(new_n254), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n266), .B1(new_n256), .B2(new_n257), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n208), .B1(new_n259), .B2(new_n267), .ZN(new_n268));
  AND2_X1   g067(.A1(new_n253), .A2(new_n255), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n269), .A2(KEYINPUT18), .A3(new_n254), .A4(new_n244), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n270), .A2(new_n258), .A3(new_n266), .A4(new_n207), .ZN(new_n271));
  AND2_X1   g070(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(G155gat), .ZN(new_n273));
  INV_X1    g072(.A(G162gat), .ZN(new_n274));
  OAI21_X1  g073(.A(KEYINPUT2), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(G141gat), .A2(G148gat), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(G141gat), .A2(G148gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n275), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  AND2_X1   g078(.A1(G155gat), .A2(G162gat), .ZN(new_n280));
  NOR2_X1   g079(.A1(G155gat), .A2(G162gat), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT79), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n277), .A2(new_n284), .A3(new_n278), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n279), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n278), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n287), .A2(new_n276), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n288), .B(new_n275), .C1(new_n282), .C2(new_n284), .ZN(new_n289));
  AND3_X1   g088(.A1(new_n286), .A2(KEYINPUT80), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT80), .B1(new_n286), .B2(new_n289), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT3), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT82), .B(KEYINPUT3), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n293), .B1(new_n286), .B2(new_n289), .ZN(new_n294));
  AND2_X1   g093(.A1(KEYINPUT71), .A2(G120gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(KEYINPUT71), .A2(G120gat), .ZN(new_n296));
  OAI21_X1  g095(.A(G113gat), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G113gat), .ZN(new_n298));
  INV_X1    g097(.A(G120gat), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT1), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(G127gat), .B(G134gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n297), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G134gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G127gat), .ZN(new_n304));
  INV_X1    g103(.A(G127gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G134gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n298), .A2(new_n299), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT1), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n309), .B1(G113gat), .B2(G120gat), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n307), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  AND3_X1   g110(.A1(new_n302), .A2(KEYINPUT81), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(KEYINPUT81), .B1(new_n302), .B2(new_n311), .ZN(new_n313));
  NOR3_X1   g112(.A1(new_n294), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n292), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n286), .A2(new_n289), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n307), .A2(new_n310), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n300), .B1(new_n298), .B2(new_n299), .ZN(new_n318));
  AOI22_X1  g117(.A1(new_n317), .A2(new_n297), .B1(new_n318), .B2(new_n307), .ZN(new_n319));
  AND3_X1   g118(.A1(new_n316), .A2(KEYINPUT4), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT4), .B1(new_n316), .B2(new_n319), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AND2_X1   g121(.A1(new_n315), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT5), .ZN(new_n324));
  NAND2_X1  g123(.A1(G225gat), .A2(G233gat), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n323), .A2(KEYINPUT85), .A3(new_n324), .A4(new_n325), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n315), .A2(new_n324), .A3(new_n322), .A4(new_n325), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT85), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n315), .A2(new_n325), .A3(new_n322), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT80), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n286), .A2(KEYINPUT80), .A3(new_n289), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n312), .A2(new_n313), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n316), .A2(new_n319), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n325), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n324), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n326), .A2(new_n329), .B1(new_n330), .B2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G57gat), .B(G85gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n342), .B(KEYINPUT84), .ZN(new_n343));
  XOR2_X1   g142(.A(KEYINPUT83), .B(KEYINPUT0), .Z(new_n344));
  XNOR2_X1  g143(.A(new_n343), .B(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G1gat), .B(G29gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n345), .B(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT6), .B1(new_n341), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n340), .A2(new_n330), .ZN(new_n349));
  AND2_X1   g148(.A1(new_n327), .A2(new_n328), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n327), .A2(new_n328), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n349), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n347), .B(KEYINPUT88), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n326), .A2(new_n329), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n347), .B1(new_n356), .B2(new_n349), .ZN(new_n357));
  AOI22_X1  g156(.A1(new_n348), .A2(new_n355), .B1(KEYINPUT6), .B2(new_n357), .ZN(new_n358));
  XOR2_X1   g157(.A(G8gat), .B(G36gat), .Z(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(KEYINPUT77), .ZN(new_n360));
  XNOR2_X1  g159(.A(G64gat), .B(G92gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT75), .B(G211gat), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT22), .B1(new_n363), .B2(G218gat), .ZN(new_n364));
  XOR2_X1   g163(.A(G197gat), .B(G204gat), .Z(new_n365));
  OR2_X1    g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  XOR2_X1   g165(.A(G211gat), .B(G218gat), .Z(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n368), .A2(KEYINPUT76), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n366), .B(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT27), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT27), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n373), .A2(KEYINPUT68), .A3(G183gat), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT67), .ZN(new_n375));
  INV_X1    g174(.A(G190gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n372), .A2(new_n374), .A3(new_n377), .A4(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT28), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT69), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n379), .A2(KEYINPUT69), .A3(new_n380), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n373), .A2(G183gat), .ZN(new_n385));
  INV_X1    g184(.A(G183gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT27), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n385), .A2(new_n387), .A3(KEYINPUT28), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n377), .A2(new_n378), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n383), .A2(new_n384), .A3(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(G169gat), .ZN(new_n393));
  INV_X1    g192(.A(G176gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT26), .ZN(new_n396));
  NAND2_X1  g195(.A1(G169gat), .A2(G176gat), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(G183gat), .A2(G190gat), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n393), .A2(new_n394), .A3(KEYINPUT26), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n392), .A2(new_n402), .ZN(new_n403));
  AND2_X1   g202(.A1(G226gat), .A2(G233gat), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT24), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n405), .A2(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n406), .B1(KEYINPUT66), .B2(new_n405), .ZN(new_n407));
  NAND3_X1  g206(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n407), .B(new_n408), .C1(G183gat), .C2(new_n389), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n393), .A2(new_n394), .A3(KEYINPUT23), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT23), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n411), .B1(G169gat), .B2(G176gat), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n410), .A2(new_n412), .A3(new_n397), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT25), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n409), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT65), .ZN(new_n417));
  OR2_X1    g216(.A1(new_n408), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n419), .A2(new_n399), .B1(new_n408), .B2(new_n417), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n413), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n416), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n403), .A2(new_n404), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT70), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n390), .B1(new_n381), .B2(new_n382), .ZN(new_n426));
  AOI211_X1 g225(.A(new_n425), .B(new_n401), .C1(new_n426), .C2(new_n384), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT70), .B1(new_n392), .B2(new_n402), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n423), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n404), .A2(KEYINPUT29), .ZN(new_n430));
  AOI211_X1 g229(.A(new_n370), .B(new_n424), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n364), .A2(new_n365), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(new_n369), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n404), .B(new_n423), .C1(new_n427), .C2(new_n428), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n421), .A2(new_n422), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n435), .B1(new_n409), .B2(new_n415), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n401), .B1(new_n426), .B2(new_n384), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n430), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n433), .B1(new_n434), .B2(new_n438), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n431), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT37), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n362), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n424), .B1(new_n429), .B2(new_n430), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n441), .B1(new_n443), .B2(new_n370), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n434), .A2(new_n438), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n433), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT38), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  AOI22_X1  g246(.A1(new_n442), .A2(new_n447), .B1(new_n440), .B2(new_n362), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n440), .A2(new_n441), .ZN(new_n449));
  INV_X1    g248(.A(new_n362), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n445), .A2(new_n370), .ZN(new_n451));
  INV_X1    g250(.A(new_n424), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n379), .A2(KEYINPUT69), .A3(new_n380), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT69), .B1(new_n379), .B2(new_n380), .ZN(new_n454));
  NOR3_X1   g253(.A1(new_n453), .A2(new_n454), .A3(new_n390), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n425), .B1(new_n455), .B2(new_n401), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n437), .A2(KEYINPUT70), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n436), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n430), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n452), .B(new_n433), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n451), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n450), .B1(new_n461), .B2(KEYINPUT37), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT38), .B1(new_n449), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n358), .A2(new_n448), .A3(new_n463), .ZN(new_n464));
  AND2_X1   g263(.A1(G228gat), .A2(G233gat), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n433), .B1(KEYINPUT29), .B2(new_n294), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT29), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT3), .B1(new_n370), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n334), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n465), .B(new_n466), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n466), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n366), .A2(new_n368), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n432), .A2(new_n367), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(new_n467), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n293), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n316), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n470), .B1(new_n465), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(KEYINPUT87), .A2(G22gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(G78gat), .B(G106gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n480), .B(G50gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(KEYINPUT86), .B(KEYINPUT31), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n481), .B(new_n482), .ZN(new_n483));
  MUX2_X1   g282(.A(new_n479), .B(G22gat), .S(new_n483), .Z(new_n484));
  XNOR2_X1  g283(.A(new_n478), .B(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n450), .B1(new_n431), .B2(new_n439), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT78), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n461), .A2(KEYINPUT78), .A3(new_n450), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n451), .A2(new_n460), .A3(new_n362), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT30), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT30), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n451), .A2(new_n460), .A3(new_n492), .A4(new_n362), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n488), .A2(new_n489), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n315), .A2(new_n322), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT89), .B1(new_n495), .B2(new_n339), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n495), .A2(KEYINPUT89), .A3(new_n339), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n336), .A2(new_n325), .A3(new_n337), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n497), .A2(KEYINPUT39), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT39), .ZN(new_n501));
  INV_X1    g300(.A(new_n498), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n501), .B1(new_n502), .B2(new_n496), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n500), .A2(new_n503), .A3(new_n353), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT40), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n500), .A2(new_n503), .A3(KEYINPUT40), .A4(new_n353), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n506), .A2(new_n355), .A3(new_n507), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n464), .B(new_n485), .C1(new_n494), .C2(new_n508), .ZN(new_n509));
  XOR2_X1   g308(.A(new_n478), .B(new_n484), .Z(new_n510));
  INV_X1    g309(.A(new_n347), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n352), .A2(KEYINPUT6), .A3(new_n511), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n349), .B(new_n347), .C1(new_n350), .C2(new_n351), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT6), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n512), .B1(new_n515), .B2(new_n357), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n488), .A2(new_n489), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n491), .A2(new_n493), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n510), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n429), .A2(new_n319), .ZN(new_n522));
  NAND2_X1  g321(.A1(G227gat), .A2(G233gat), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n319), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n525), .B(new_n423), .C1(new_n427), .C2(new_n428), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n522), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT32), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT33), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(KEYINPUT72), .B(G71gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(G99gat), .ZN(new_n532));
  XOR2_X1   g331(.A(G15gat), .B(G43gat), .Z(new_n533));
  XOR2_X1   g332(.A(new_n532), .B(new_n533), .Z(new_n534));
  NAND3_X1  g333(.A1(new_n528), .A2(new_n530), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n534), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n527), .B(KEYINPUT32), .C1(new_n529), .C2(new_n536), .ZN(new_n537));
  AND2_X1   g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT34), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n458), .A2(new_n525), .ZN(new_n540));
  INV_X1    g339(.A(new_n526), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n539), .B(new_n523), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT74), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n524), .B1(new_n522), .B2(new_n526), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT74), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(new_n545), .A3(new_n539), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n523), .B1(new_n540), .B2(new_n541), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT34), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n543), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n538), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n537), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n543), .A2(new_n546), .A3(new_n548), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(KEYINPUT36), .B1(new_n550), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n551), .A2(KEYINPUT73), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT73), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n535), .A2(new_n556), .A3(new_n537), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n555), .A2(new_n557), .A3(new_n552), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT36), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n559), .B1(new_n538), .B2(new_n549), .ZN(new_n560));
  AND2_X1   g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n509), .B(new_n521), .C1(new_n554), .C2(new_n561), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n494), .A2(new_n516), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n485), .B1(new_n551), .B2(new_n552), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n563), .A2(new_n558), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT35), .ZN(new_n567));
  AND3_X1   g366(.A1(new_n550), .A2(new_n485), .A3(new_n553), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n341), .A2(new_n353), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n512), .B1(new_n569), .B2(new_n515), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT35), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n570), .A2(new_n494), .A3(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n567), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n272), .B1(new_n562), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT21), .ZN(new_n577));
  NAND2_X1  g376(.A1(G71gat), .A2(G78gat), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT9), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(G57gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(G64gat), .ZN(new_n582));
  INV_X1    g381(.A(G64gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(G57gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(G71gat), .ZN(new_n586));
  INV_X1    g385(.A(G78gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AND3_X1   g387(.A1(new_n588), .A2(KEYINPUT96), .A3(new_n578), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT96), .B1(new_n588), .B2(new_n578), .ZN(new_n590));
  OAI211_X1 g389(.A(new_n580), .B(new_n585), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n585), .A2(new_n580), .ZN(new_n592));
  NAND3_X1  g391(.A1(KEYINPUT95), .A2(G71gat), .A3(G78gat), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT95), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n592), .A2(new_n588), .A3(new_n593), .A4(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n237), .B1(new_n577), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT97), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(new_n273), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n600), .B(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n597), .A2(new_n577), .ZN(new_n605));
  NAND2_X1  g404(.A1(G231gat), .A2(G233gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  OR2_X1    g406(.A1(new_n607), .A2(new_n305), .ZN(new_n608));
  XOR2_X1   g407(.A(G183gat), .B(G211gat), .Z(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n607), .A2(new_n305), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n608), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n610), .B1(new_n608), .B2(new_n611), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n604), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n600), .B(new_n602), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n607), .B(new_n305), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(new_n609), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n616), .A2(new_n618), .A3(new_n612), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(G190gat), .B(G218gat), .Z(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(G99gat), .A2(G106gat), .ZN(new_n623));
  INV_X1    g422(.A(G85gat), .ZN(new_n624));
  INV_X1    g423(.A(G92gat), .ZN(new_n625));
  AOI22_X1  g424(.A1(KEYINPUT8), .A2(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND4_X1  g425(.A1(KEYINPUT98), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n627));
  NAND3_X1  g426(.A1(KEYINPUT98), .A2(G85gat), .A3(G92gat), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT7), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n626), .A2(new_n627), .A3(new_n630), .ZN(new_n631));
  OR2_X1    g430(.A1(G99gat), .A2(G106gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n623), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n626), .A2(new_n633), .A3(new_n627), .A4(new_n630), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AND2_X1   g436(.A1(G232gat), .A2(G233gat), .ZN(new_n638));
  AOI22_X1  g437(.A1(new_n248), .A2(new_n637), .B1(KEYINPUT41), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n635), .A2(new_n636), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n225), .A2(new_n241), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n622), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n638), .A2(KEYINPUT41), .ZN(new_n644));
  XNOR2_X1  g443(.A(G134gat), .B(G162gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n639), .A2(new_n641), .A3(new_n622), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n643), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n646), .ZN(new_n649));
  INV_X1    g448(.A(new_n647), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n649), .B1(new_n650), .B2(new_n642), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(G230gat), .A2(G233gat), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n631), .A2(KEYINPUT99), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT99), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n626), .A2(new_n656), .A3(new_n627), .A4(new_n630), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n633), .A2(KEYINPUT100), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT100), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n632), .A2(new_n659), .A3(new_n623), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n655), .A2(new_n657), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT101), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AND3_X1   g463(.A1(new_n591), .A2(new_n596), .A3(new_n636), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n655), .A2(KEYINPUT101), .A3(new_n661), .A4(new_n657), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT10), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n597), .A2(new_n640), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n637), .A2(KEYINPUT10), .A3(new_n591), .A4(new_n596), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n654), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n653), .B1(new_n667), .B2(new_n669), .ZN(new_n673));
  XNOR2_X1  g472(.A(G120gat), .B(G148gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(G176gat), .B(G204gat), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n674), .B(new_n675), .Z(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  OR3_X1    g476(.A1(new_n672), .A2(new_n673), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n677), .B1(new_n672), .B2(new_n673), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n620), .A2(new_n652), .A3(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n576), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n684), .A2(new_n516), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(new_n227), .ZN(G1324gat));
  INV_X1    g485(.A(KEYINPUT42), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n684), .A2(new_n494), .ZN(new_n688));
  XOR2_X1   g487(.A(KEYINPUT16), .B(G8gat), .Z(new_n689));
  AOI21_X1  g488(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(G8gat), .B1(new_n684), .B2(new_n494), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT102), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n687), .A2(KEYINPUT102), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n693), .B1(new_n689), .B2(new_n694), .ZN(new_n695));
  AOI22_X1  g494(.A1(new_n690), .A2(new_n691), .B1(new_n688), .B2(new_n695), .ZN(G1325gat));
  AOI21_X1  g495(.A(new_n554), .B1(new_n558), .B2(new_n560), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(G15gat), .B1(new_n684), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n550), .A2(new_n553), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n268), .A2(new_n271), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n485), .B1(new_n508), .B2(new_n494), .ZN(new_n703));
  AND3_X1   g502(.A1(new_n358), .A2(new_n448), .A3(new_n463), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n521), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n705), .A2(new_n697), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n545), .B1(new_n544), .B2(new_n539), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n544), .A2(new_n539), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AOI22_X1  g508(.A1(new_n551), .A2(KEYINPUT73), .B1(new_n709), .B2(new_n546), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n564), .B1(new_n710), .B2(new_n557), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n571), .B1(new_n711), .B2(new_n563), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n700), .A2(new_n572), .A3(new_n510), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OAI211_X1 g513(.A(new_n701), .B(new_n702), .C1(new_n706), .C2(new_n714), .ZN(new_n715));
  OR2_X1    g514(.A1(new_n682), .A2(G15gat), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n699), .B1(new_n715), .B2(new_n716), .ZN(G1326gat));
  NOR2_X1   g516(.A1(new_n684), .A2(new_n485), .ZN(new_n718));
  XOR2_X1   g517(.A(KEYINPUT43), .B(G22gat), .Z(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1327gat));
  AOI21_X1  g519(.A(new_n652), .B1(new_n562), .B2(new_n575), .ZN(new_n721));
  INV_X1    g520(.A(new_n620), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n681), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n723), .A2(new_n272), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n725), .A2(G29gat), .A3(new_n516), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n726), .B(KEYINPUT45), .Z(new_n727));
  OAI21_X1  g526(.A(KEYINPUT103), .B1(new_n712), .B2(new_n713), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT103), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n567), .A2(new_n574), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n706), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n652), .A2(KEYINPUT44), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n734));
  OAI22_X1  g533(.A1(new_n731), .A2(new_n733), .B1(new_n721), .B2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n724), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n736), .A2(new_n516), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n727), .B1(new_n220), .B2(new_n738), .ZN(G1328gat));
  INV_X1    g538(.A(new_n652), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n722), .A2(new_n740), .A3(new_n681), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT46), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n218), .B1(new_n742), .B2(KEYINPUT104), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n741), .A2(new_n494), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n576), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n742), .A2(KEYINPUT104), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n745), .B(new_n746), .Z(new_n747));
  NOR3_X1   g546(.A1(new_n736), .A2(new_n494), .A3(new_n737), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n747), .B1(new_n748), .B2(new_n218), .ZN(G1329gat));
  INV_X1    g548(.A(KEYINPUT109), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n741), .A2(G43gat), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(KEYINPUT107), .B1(new_n715), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT107), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n576), .A2(new_n754), .A3(new_n701), .A4(new_n751), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT47), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n728), .A2(new_n730), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n733), .B1(new_n758), .B2(new_n562), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n562), .A2(new_n575), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n734), .B1(new_n760), .B2(new_n740), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n697), .B(new_n724), .C1(new_n759), .C2(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n213), .B1(new_n762), .B2(KEYINPUT108), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT108), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n735), .A2(new_n764), .A3(new_n697), .A4(new_n724), .ZN(new_n765));
  AOI211_X1 g564(.A(new_n750), .B(new_n757), .C1(new_n763), .C2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n762), .A2(KEYINPUT108), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n767), .A2(G43gat), .A3(new_n765), .ZN(new_n768));
  INV_X1    g567(.A(new_n757), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT109), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT106), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n762), .A2(new_n771), .A3(G43gat), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n771), .B1(new_n762), .B2(G43gat), .ZN(new_n773));
  INV_X1    g572(.A(new_n756), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  XOR2_X1   g574(.A(KEYINPUT105), .B(KEYINPUT47), .Z(new_n776));
  OAI22_X1  g575(.A1(new_n766), .A2(new_n770), .B1(new_n775), .B2(new_n776), .ZN(G1330gat));
  NAND2_X1  g576(.A1(new_n510), .A2(new_n212), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT110), .ZN(new_n779));
  OAI22_X1  g578(.A1(new_n725), .A2(new_n778), .B1(new_n779), .B2(KEYINPUT48), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n735), .A2(new_n510), .A3(new_n724), .ZN(new_n781));
  INV_X1    g580(.A(new_n212), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n779), .A2(KEYINPUT48), .ZN(new_n784));
  XOR2_X1   g583(.A(new_n783), .B(new_n784), .Z(G1331gat));
  NAND2_X1  g584(.A1(new_n758), .A2(new_n562), .ZN(new_n786));
  NOR4_X1   g585(.A1(new_n722), .A2(new_n702), .A3(new_n740), .A4(new_n681), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(new_n516), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(new_n581), .ZN(G1332gat));
  NOR2_X1   g589(.A1(new_n788), .A2(new_n494), .ZN(new_n791));
  NOR2_X1   g590(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n792));
  AND2_X1   g591(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n794), .B1(new_n791), .B2(new_n792), .ZN(G1333gat));
  OAI21_X1  g594(.A(G71gat), .B1(new_n788), .B2(new_n698), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n701), .A2(new_n586), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n796), .B1(new_n788), .B2(new_n797), .ZN(new_n798));
  XOR2_X1   g597(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n799));
  XNOR2_X1  g598(.A(new_n798), .B(new_n799), .ZN(G1334gat));
  NOR2_X1   g599(.A1(new_n788), .A2(new_n485), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(new_n587), .ZN(G1335gat));
  NAND2_X1  g601(.A1(new_n722), .A2(new_n272), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n803), .A2(new_n681), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n735), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(G85gat), .B1(new_n805), .B2(new_n516), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n803), .A2(new_n652), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n786), .A2(KEYINPUT51), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(KEYINPUT51), .B1(new_n786), .B2(new_n807), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n517), .A2(new_n624), .A3(new_n680), .ZN(new_n811));
  XOR2_X1   g610(.A(new_n811), .B(KEYINPUT112), .Z(new_n812));
  OAI21_X1  g611(.A(new_n806), .B1(new_n810), .B2(new_n812), .ZN(G1336gat));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n494), .A2(G92gat), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n680), .B(new_n815), .C1(new_n808), .C2(new_n809), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n814), .B1(new_n816), .B2(KEYINPUT113), .ZN(new_n817));
  OAI21_X1  g616(.A(G92gat), .B1(new_n805), .B2(new_n494), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n816), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n817), .B(new_n819), .ZN(G1337gat));
  INV_X1    g619(.A(G99gat), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n805), .A2(new_n821), .A3(new_n698), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n701), .B(new_n680), .C1(new_n808), .C2(new_n809), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n822), .B1(new_n821), .B2(new_n823), .ZN(G1338gat));
  NAND3_X1  g623(.A1(new_n735), .A2(new_n510), .A3(new_n804), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(G106gat), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n485), .A2(G106gat), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n680), .B(new_n827), .C1(new_n808), .C2(new_n809), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT114), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n826), .B(KEYINPUT115), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n829), .B1(KEYINPUT115), .B2(KEYINPUT53), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n832), .B1(new_n825), .B2(G106gat), .ZN(new_n833));
  AOI22_X1  g632(.A1(new_n830), .A2(new_n831), .B1(new_n828), .B2(new_n833), .ZN(G1339gat));
  INV_X1    g633(.A(KEYINPUT116), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n671), .A2(new_n654), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n670), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT54), .ZN(new_n838));
  OAI21_X1  g637(.A(KEYINPUT55), .B1(new_n838), .B2(new_n672), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n670), .A2(new_n671), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n840), .A2(new_n841), .A3(new_n653), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n677), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n678), .B1(new_n839), .B2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n672), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n841), .B1(new_n670), .B2(new_n836), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n676), .B1(new_n672), .B2(new_n841), .ZN(new_n848));
  AOI21_X1  g647(.A(KEYINPUT55), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n835), .B1(new_n844), .B2(new_n849), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n672), .A2(new_n673), .A3(new_n677), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT55), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n852), .B1(new_n845), .B2(new_n846), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n851), .B1(new_n853), .B2(new_n848), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n838), .A2(new_n672), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n852), .B1(new_n843), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n854), .A2(new_n856), .A3(KEYINPUT116), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n850), .A2(new_n857), .A3(new_n702), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n254), .B1(new_n269), .B2(new_n244), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n263), .A2(new_n265), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n206), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n680), .A2(new_n861), .A3(new_n271), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n740), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n740), .A2(new_n861), .A3(new_n271), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n865), .A2(new_n850), .A3(new_n857), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n722), .B1(new_n863), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n682), .A2(new_n702), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n871), .A2(new_n517), .A3(new_n494), .A4(new_n568), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n872), .A2(new_n298), .A3(new_n272), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n516), .B1(new_n868), .B2(new_n870), .ZN(new_n874));
  INV_X1    g673(.A(new_n711), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n875), .A2(new_n520), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n702), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n873), .B1(new_n298), .B2(new_n879), .ZN(G1340gat));
  OAI21_X1  g679(.A(G120gat), .B1(new_n872), .B2(new_n681), .ZN(new_n881));
  OR3_X1    g680(.A1(new_n681), .A2(new_n296), .A3(new_n295), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n881), .B1(new_n877), .B2(new_n882), .ZN(G1341gat));
  OAI21_X1  g682(.A(G127gat), .B1(new_n872), .B2(new_n722), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n620), .A2(new_n305), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n884), .B1(new_n877), .B2(new_n885), .ZN(G1342gat));
  NOR3_X1   g685(.A1(new_n877), .A2(G134gat), .A3(new_n652), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n888), .A2(KEYINPUT56), .ZN(new_n889));
  OAI21_X1  g688(.A(G134gat), .B1(new_n872), .B2(new_n652), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(KEYINPUT56), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(G1343gat));
  NOR3_X1   g691(.A1(new_n697), .A2(new_n516), .A3(new_n520), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT57), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n485), .A2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n854), .A2(new_n856), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n862), .B1(new_n272), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n652), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n620), .B1(new_n899), .B2(new_n866), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT117), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n869), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n702), .A2(new_n856), .A3(new_n854), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n740), .B1(new_n903), .B2(new_n862), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n722), .B1(new_n867), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT117), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n896), .B1(new_n902), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(KEYINPUT57), .B1(new_n871), .B2(new_n510), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n893), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(G141gat), .B1(new_n909), .B2(new_n272), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n697), .A2(new_n520), .A3(new_n485), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n874), .A2(new_n911), .ZN(new_n912));
  OR3_X1    g711(.A1(new_n912), .A2(G141gat), .A3(new_n272), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g714(.A(KEYINPUT121), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n896), .B1(new_n868), .B2(new_n870), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n897), .A2(new_n864), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n918), .B1(new_n898), .B2(new_n652), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n870), .B1(new_n919), .B2(new_n620), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT119), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI211_X1 g721(.A(new_n870), .B(KEYINPUT119), .C1(new_n919), .C2(new_n620), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n922), .A2(new_n510), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n917), .B1(new_n924), .B2(new_n894), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n893), .A2(new_n680), .ZN(new_n926));
  OAI21_X1  g725(.A(KEYINPUT120), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(new_n926), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT120), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n485), .B1(new_n920), .B2(new_n921), .ZN(new_n930));
  AOI21_X1  g729(.A(KEYINPUT57), .B1(new_n930), .B2(new_n923), .ZN(new_n931));
  OAI211_X1 g730(.A(new_n928), .B(new_n929), .C1(new_n931), .C2(new_n917), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n927), .A2(G148gat), .A3(new_n932), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n680), .B(new_n893), .C1(new_n907), .C2(new_n908), .ZN(new_n934));
  INV_X1    g733(.A(G148gat), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n935), .A2(KEYINPUT59), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(KEYINPUT118), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT118), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n934), .A2(new_n939), .A3(new_n936), .ZN(new_n940));
  AOI22_X1  g739(.A1(new_n933), .A2(KEYINPUT59), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n912), .A2(G148gat), .A3(new_n681), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n916), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(new_n942), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n938), .A2(new_n940), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT59), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n924), .A2(new_n894), .ZN(new_n947));
  INV_X1    g746(.A(new_n917), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n926), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n935), .B1(new_n949), .B2(new_n929), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n946), .B1(new_n950), .B2(new_n927), .ZN(new_n951));
  OAI211_X1 g750(.A(KEYINPUT121), .B(new_n944), .C1(new_n945), .C2(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n943), .A2(new_n952), .ZN(G1345gat));
  NOR3_X1   g752(.A1(new_n912), .A2(G155gat), .A3(new_n722), .ZN(new_n954));
  INV_X1    g753(.A(new_n909), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(new_n620), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n954), .B1(new_n956), .B2(G155gat), .ZN(new_n957));
  XOR2_X1   g756(.A(new_n957), .B(KEYINPUT122), .Z(G1346gat));
  INV_X1    g757(.A(new_n912), .ZN(new_n959));
  AOI21_X1  g758(.A(G162gat), .B1(new_n959), .B2(new_n740), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n652), .A2(new_n274), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n960), .B1(new_n955), .B2(new_n961), .ZN(G1347gat));
  AND4_X1   g761(.A1(new_n516), .A2(new_n871), .A3(new_n520), .A4(new_n568), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n393), .B1(new_n963), .B2(new_n702), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT123), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n517), .B1(new_n868), .B2(new_n870), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n875), .A2(new_n494), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(new_n968), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n969), .A2(new_n393), .A3(new_n702), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n965), .A2(new_n970), .ZN(G1348gat));
  NAND3_X1  g770(.A1(new_n969), .A2(new_n394), .A3(new_n680), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n963), .A2(new_n680), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n972), .B1(new_n973), .B2(new_n394), .ZN(G1349gat));
  AOI21_X1  g773(.A(new_n386), .B1(new_n963), .B2(new_n620), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n620), .A2(new_n385), .A3(new_n387), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n975), .B1(new_n969), .B2(new_n976), .ZN(new_n977));
  XOR2_X1   g776(.A(new_n977), .B(KEYINPUT60), .Z(G1350gat));
  AOI21_X1  g777(.A(new_n376), .B1(new_n963), .B2(new_n740), .ZN(new_n979));
  XNOR2_X1  g778(.A(new_n979), .B(KEYINPUT61), .ZN(new_n980));
  NOR3_X1   g779(.A1(new_n968), .A2(new_n389), .A3(new_n652), .ZN(new_n981));
  OR2_X1    g780(.A1(new_n980), .A2(new_n981), .ZN(G1351gat));
  NAND3_X1  g781(.A1(new_n698), .A2(new_n516), .A3(new_n520), .ZN(new_n983));
  XNOR2_X1  g782(.A(new_n983), .B(KEYINPUT125), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n984), .A2(new_n925), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n985), .A2(new_n702), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n986), .A2(G197gat), .ZN(new_n987));
  NOR3_X1   g786(.A1(new_n697), .A2(new_n494), .A3(new_n485), .ZN(new_n988));
  AND2_X1   g787(.A1(new_n966), .A2(new_n988), .ZN(new_n989));
  INV_X1    g788(.A(G197gat), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n989), .A2(new_n990), .A3(new_n702), .ZN(new_n991));
  XNOR2_X1  g790(.A(new_n991), .B(KEYINPUT124), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n987), .A2(new_n992), .ZN(new_n993));
  INV_X1    g792(.A(KEYINPUT126), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n987), .A2(KEYINPUT126), .A3(new_n992), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(G1352gat));
  INV_X1    g796(.A(new_n989), .ZN(new_n998));
  NOR3_X1   g797(.A1(new_n998), .A2(G204gat), .A3(new_n681), .ZN(new_n999));
  XNOR2_X1  g798(.A(new_n999), .B(KEYINPUT62), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n680), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1001), .A2(G204gat), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1000), .A2(new_n1002), .ZN(G1353gat));
  NOR3_X1   g802(.A1(new_n925), .A2(new_n722), .A3(new_n983), .ZN(new_n1004));
  INV_X1    g803(.A(G211gat), .ZN(new_n1005));
  NOR2_X1   g804(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g805(.A(new_n1006), .B(KEYINPUT63), .ZN(new_n1007));
  OR2_X1    g806(.A1(new_n722), .A2(new_n363), .ZN(new_n1008));
  OAI21_X1  g807(.A(new_n1007), .B1(new_n998), .B2(new_n1008), .ZN(G1354gat));
  AOI21_X1  g808(.A(G218gat), .B1(new_n989), .B2(new_n740), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n740), .A2(G218gat), .ZN(new_n1011));
  XOR2_X1   g810(.A(new_n1011), .B(KEYINPUT127), .Z(new_n1012));
  AOI21_X1  g811(.A(new_n1010), .B1(new_n985), .B2(new_n1012), .ZN(G1355gat));
endmodule


