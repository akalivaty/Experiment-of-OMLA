//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 0 1 1 0 0 1 1 0 1 1 0 1 0 1 0 1 1 1 1 0 1 1 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 1 0 0 1 0 1 1 0 1 1 1 1 0 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995;
  INV_X1    g000(.A(G125), .ZN(new_n187));
  OR3_X1    g001(.A1(new_n187), .A2(KEYINPUT16), .A3(G140), .ZN(new_n188));
  XOR2_X1   g002(.A(G125), .B(G140), .Z(new_n189));
  INV_X1    g003(.A(KEYINPUT16), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n188), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  OAI211_X1 g007(.A(G146), .B(new_n188), .C1(new_n189), .C2(new_n190), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT68), .B(G128), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(KEYINPUT23), .A3(G119), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  AOI21_X1  g012(.A(KEYINPUT23), .B1(new_n198), .B2(G119), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n198), .A2(G119), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n197), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G110), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n200), .B1(new_n196), .B2(G119), .ZN(new_n204));
  XOR2_X1   g018(.A(KEYINPUT24), .B(G110), .Z(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n195), .A2(new_n203), .A3(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(G125), .B(G140), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(new_n192), .ZN(new_n209));
  XOR2_X1   g023(.A(KEYINPUT78), .B(G110), .Z(new_n210));
  NOR2_X1   g024(.A1(new_n202), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n204), .A2(new_n205), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n194), .B(new_n209), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n207), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT80), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT80), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n207), .A2(new_n213), .A3(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G953), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(G221), .A3(G234), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n219), .B(KEYINPUT79), .ZN(new_n220));
  XOR2_X1   g034(.A(KEYINPUT22), .B(G137), .Z(new_n221));
  XNOR2_X1  g035(.A(new_n220), .B(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n215), .A2(new_n217), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n215), .B1(new_n217), .B2(new_n222), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G217), .ZN(new_n227));
  INV_X1    g041(.A(G902), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n227), .B1(G234), .B2(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(G902), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT81), .B1(new_n226), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT81), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n233), .B(new_n230), .C1(new_n224), .C2(new_n225), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n217), .A2(new_n222), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(KEYINPUT80), .A3(new_n214), .ZN(new_n236));
  AOI21_X1  g050(.A(G902), .B1(new_n236), .B2(new_n223), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT25), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n229), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  AOI211_X1 g053(.A(KEYINPUT25), .B(G902), .C1(new_n236), .C2(new_n223), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n232), .B(new_n234), .C1(new_n239), .C2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT29), .ZN(new_n242));
  NAND2_X1  g056(.A1(KEYINPUT11), .A2(G134), .ZN(new_n243));
  OAI21_X1  g057(.A(KEYINPUT66), .B1(new_n243), .B2(G137), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT66), .ZN(new_n245));
  INV_X1    g059(.A(G137), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n245), .A2(new_n246), .A3(KEYINPUT11), .A4(G134), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G134), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT65), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT65), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G134), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n250), .A2(new_n252), .A3(G137), .ZN(new_n253));
  AOI21_X1  g067(.A(G137), .B1(new_n250), .B2(new_n252), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n248), .B(new_n253), .C1(new_n254), .C2(KEYINPUT11), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G131), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT11), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT65), .B(G134), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n257), .B1(new_n258), .B2(G137), .ZN(new_n259));
  INV_X1    g073(.A(G131), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n259), .A2(new_n260), .A3(new_n248), .A4(new_n253), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n192), .A2(G143), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT64), .ZN(new_n264));
  INV_X1    g078(.A(G143), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n264), .B1(new_n265), .B2(G146), .ZN(new_n266));
  NOR3_X1   g080(.A1(new_n192), .A2(KEYINPUT64), .A3(G143), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n263), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  AND2_X1   g082(.A1(KEYINPUT0), .A2(G128), .ZN(new_n269));
  NOR2_X1   g083(.A1(KEYINPUT0), .A2(G128), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(G143), .B(G146), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n268), .A2(new_n271), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n262), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n246), .A2(G134), .ZN(new_n275));
  OAI21_X1  g089(.A(G131), .B1(new_n254), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n261), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT1), .B1(new_n265), .B2(G146), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT67), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT67), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n263), .A2(new_n280), .A3(KEYINPUT1), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n198), .A2(KEYINPUT68), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT68), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G128), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n279), .A2(new_n281), .A3(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n198), .A2(KEYINPUT1), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n286), .A2(new_n268), .B1(new_n272), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(KEYINPUT71), .B1(new_n277), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n286), .A2(new_n268), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n265), .A2(G146), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n287), .A2(new_n263), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT71), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n293), .A2(new_n294), .A3(new_n261), .A4(new_n276), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n274), .A2(new_n289), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT72), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT2), .ZN(new_n298));
  INV_X1    g112(.A(G113), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(new_n299), .A3(KEYINPUT69), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT69), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n301), .B1(KEYINPUT2), .B2(G113), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(KEYINPUT2), .A2(G113), .ZN(new_n304));
  XNOR2_X1  g118(.A(G116), .B(G119), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n305), .B1(new_n303), .B2(new_n304), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT70), .ZN(new_n308));
  NOR3_X1   g122(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n303), .A2(new_n304), .ZN(new_n310));
  INV_X1    g124(.A(new_n305), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI22_X1  g126(.A1(new_n300), .A2(new_n302), .B1(KEYINPUT2), .B2(G113), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n305), .ZN(new_n314));
  AOI21_X1  g128(.A(KEYINPUT70), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n297), .B1(new_n309), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n308), .B1(new_n306), .B2(new_n307), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n312), .A2(KEYINPUT70), .A3(new_n314), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n318), .A3(KEYINPUT72), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  OR2_X1    g134(.A1(new_n296), .A2(new_n320), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n274), .A2(new_n289), .A3(KEYINPUT30), .A4(new_n295), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n309), .A2(new_n315), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT30), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n277), .A2(new_n288), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n272), .A2(new_n269), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n291), .A2(KEYINPUT64), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n264), .A2(new_n265), .A3(G146), .ZN(new_n328));
  AOI22_X1  g142(.A1(new_n327), .A2(new_n328), .B1(G143), .B2(new_n192), .ZN(new_n329));
  INV_X1    g143(.A(new_n271), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n326), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n331), .B1(new_n256), .B2(new_n261), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n324), .B1(new_n325), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n322), .A2(new_n323), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n321), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G237), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT73), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT73), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G237), .ZN(new_n339));
  AOI21_X1  g153(.A(G953), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G210), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n341), .B(KEYINPUT27), .ZN(new_n342));
  XNOR2_X1  g156(.A(KEYINPUT26), .B(G101), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n342), .B(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n335), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n323), .B1(new_n325), .B2(new_n332), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT74), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT74), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n323), .B(new_n349), .C1(new_n325), .C2(new_n332), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n296), .A2(new_n320), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT28), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n293), .A2(new_n261), .A3(new_n276), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n316), .A2(new_n274), .A3(new_n319), .A4(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT75), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT28), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n356), .B1(new_n355), .B2(new_n357), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n353), .A2(new_n360), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n242), .B(new_n346), .C1(new_n361), .C2(new_n345), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n355), .A2(new_n357), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT75), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n296), .A2(new_n320), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n357), .B1(new_n321), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n345), .A2(new_n242), .ZN(new_n370));
  AOI21_X1  g184(.A(G902), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n362), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(G472), .A2(G902), .ZN(new_n373));
  XOR2_X1   g187(.A(new_n373), .B(KEYINPUT76), .Z(new_n374));
  AND2_X1   g188(.A1(new_n348), .A2(new_n350), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n357), .B1(new_n375), .B2(new_n321), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n345), .B1(new_n376), .B2(new_n366), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT31), .ZN(new_n378));
  INV_X1    g192(.A(new_n334), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n344), .B1(new_n296), .B2(new_n320), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n321), .A2(new_n334), .A3(KEYINPUT31), .A4(new_n344), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n374), .B1(new_n377), .B2(new_n383), .ZN(new_n384));
  AOI22_X1  g198(.A1(new_n372), .A2(G472), .B1(new_n384), .B2(KEYINPUT32), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT77), .ZN(new_n386));
  AOI22_X1  g200(.A1(new_n361), .A2(new_n345), .B1(new_n381), .B2(new_n382), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n386), .B1(new_n387), .B2(new_n374), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT32), .ZN(new_n389));
  INV_X1    g203(.A(new_n374), .ZN(new_n390));
  INV_X1    g204(.A(new_n383), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n344), .B1(new_n353), .B2(new_n360), .ZN(new_n392));
  OAI211_X1 g206(.A(KEYINPUT77), .B(new_n390), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n388), .A2(new_n389), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n241), .B1(new_n385), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT82), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n396), .A2(KEYINPUT3), .ZN(new_n397));
  INV_X1    g211(.A(G104), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(G107), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n396), .A2(KEYINPUT3), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n397), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n398), .A2(G107), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT3), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(KEYINPUT82), .ZN(new_n404));
  INV_X1    g218(.A(G107), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G104), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n402), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(G101), .B1(new_n401), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n405), .A2(G104), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n409), .B1(new_n397), .B2(new_n399), .ZN(new_n410));
  INV_X1    g224(.A(G101), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n403), .A2(KEYINPUT82), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n404), .B1(new_n412), .B2(new_n406), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n410), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n408), .A2(KEYINPUT4), .A3(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(KEYINPUT83), .B(KEYINPUT4), .ZN(new_n416));
  OAI211_X1 g230(.A(G101), .B(new_n416), .C1(new_n401), .C2(new_n407), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n317), .A2(new_n415), .A3(new_n318), .A4(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n305), .A2(KEYINPUT5), .ZN(new_n419));
  INV_X1    g233(.A(G116), .ZN(new_n420));
  NOR3_X1   g234(.A1(new_n420), .A2(KEYINPUT5), .A3(G119), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n421), .A2(new_n299), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(G101), .B1(new_n399), .B2(new_n409), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n414), .A2(new_n314), .A3(new_n423), .A4(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n418), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(G110), .B(G122), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n418), .A2(new_n425), .A3(new_n427), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n429), .A2(KEYINPUT6), .A3(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT6), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n426), .A2(new_n432), .A3(new_n428), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT86), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n434), .B1(new_n273), .B2(new_n187), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n288), .A2(new_n187), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n331), .A2(KEYINPUT86), .A3(G125), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n218), .A2(G224), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n438), .B(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n431), .A2(new_n433), .A3(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n436), .B1(new_n187), .B2(new_n273), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n439), .A2(KEYINPUT7), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AND2_X1   g259(.A1(new_n430), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n438), .ZN(new_n447));
  INV_X1    g261(.A(new_n444), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT87), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n425), .A2(new_n449), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n313), .A2(new_n305), .B1(new_n419), .B2(new_n422), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n451), .A2(KEYINPUT87), .A3(new_n414), .A4(new_n424), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n414), .A2(new_n424), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n314), .A2(new_n423), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n450), .A2(new_n452), .A3(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n427), .B(KEYINPUT8), .ZN(new_n457));
  AOI22_X1  g271(.A1(new_n447), .A2(new_n448), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(G902), .B1(new_n446), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n442), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(G210), .B1(G237), .B2(G902), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n442), .A2(new_n459), .A3(new_n461), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(KEYINPUT88), .A3(new_n464), .ZN(new_n465));
  OR2_X1    g279(.A1(new_n464), .A2(KEYINPUT88), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(G214), .B1(G237), .B2(G902), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(KEYINPUT9), .B(G234), .ZN(new_n471));
  OAI21_X1  g285(.A(G221), .B1(new_n471), .B2(G902), .ZN(new_n472));
  XNOR2_X1  g286(.A(G110), .B(G140), .ZN(new_n473));
  INV_X1    g287(.A(G227), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(G953), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n473), .B(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n198), .B1(new_n263), .B2(KEYINPUT1), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n292), .B1(new_n477), .B2(new_n272), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n414), .A2(new_n424), .A3(new_n478), .ZN(new_n479));
  XOR2_X1   g293(.A(KEYINPUT85), .B(KEYINPUT10), .Z(new_n480));
  NAND3_X1  g294(.A1(new_n414), .A2(KEYINPUT10), .A3(new_n424), .ZN(new_n481));
  OAI22_X1  g295(.A1(new_n479), .A2(new_n480), .B1(new_n288), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n415), .A2(new_n273), .A3(new_n417), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(KEYINPUT84), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT84), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n415), .A2(new_n485), .A3(new_n273), .A4(new_n417), .ZN(new_n486));
  AOI211_X1 g300(.A(new_n262), .B(new_n482), .C1(new_n484), .C2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n262), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n484), .A2(new_n486), .ZN(new_n489));
  INV_X1    g303(.A(new_n482), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n476), .B1(new_n487), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n482), .B1(new_n484), .B2(new_n486), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n476), .B1(new_n493), .B2(new_n488), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n288), .A2(new_n453), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n414), .A2(new_n478), .A3(new_n424), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n497), .A2(KEYINPUT12), .A3(new_n262), .ZN(new_n498));
  AOI21_X1  g312(.A(KEYINPUT12), .B1(new_n497), .B2(new_n262), .ZN(new_n499));
  OR2_X1    g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  AOI211_X1 g315(.A(G469), .B(G902), .C1(new_n492), .C2(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n498), .A2(new_n499), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n476), .B1(new_n487), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n489), .A2(new_n490), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n262), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n494), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n504), .A2(new_n507), .A3(G469), .ZN(new_n508));
  NAND2_X1  g322(.A1(G469), .A2(G902), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n472), .B1(new_n502), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(G234), .A2(G237), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(G952), .A3(new_n218), .ZN(new_n514));
  XOR2_X1   g328(.A(KEYINPUT21), .B(G898), .Z(new_n515));
  NAND3_X1  g329(.A1(new_n513), .A2(G902), .A3(G953), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  XOR2_X1   g331(.A(new_n517), .B(KEYINPUT97), .Z(new_n518));
  AOI21_X1  g332(.A(KEYINPUT13), .B1(new_n265), .B2(G128), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n519), .B(KEYINPUT93), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n198), .A2(G143), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n196), .A2(G143), .B1(KEYINPUT13), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n249), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n196), .A2(G143), .ZN(new_n524));
  INV_X1    g338(.A(new_n521), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n258), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(G122), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(G116), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n420), .A2(G122), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(G107), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n528), .A2(new_n529), .A3(new_n405), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n526), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n523), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n528), .A2(KEYINPUT14), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n530), .A2(new_n536), .A3(G107), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n528), .B(new_n529), .C1(KEYINPUT14), .C2(new_n405), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n524), .A2(new_n525), .ZN(new_n540));
  INV_X1    g354(.A(new_n258), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n539), .B1(new_n542), .B2(new_n526), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n471), .A2(new_n227), .A3(G953), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n535), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT93), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n519), .B(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n521), .A2(KEYINPUT13), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n549), .B1(new_n285), .B2(new_n265), .ZN(new_n550));
  OAI21_X1  g364(.A(G134), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n551), .A2(new_n526), .A3(new_n533), .ZN(new_n552));
  INV_X1    g366(.A(new_n526), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n258), .B1(new_n524), .B2(new_n525), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n538), .B(new_n537), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n544), .B1(new_n552), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n228), .B1(new_n546), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(G478), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n558), .A2(KEYINPUT15), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n557), .A2(KEYINPUT94), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT94), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n545), .B1(new_n535), .B2(new_n543), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n552), .A2(new_n555), .A3(new_n544), .ZN(new_n563));
  AOI21_X1  g377(.A(G902), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n559), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n561), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n560), .A2(new_n566), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n228), .B(new_n565), .C1(new_n546), .C2(new_n556), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT95), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n564), .A2(KEYINPUT95), .A3(new_n565), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AND3_X1   g386(.A1(new_n567), .A2(new_n572), .A3(KEYINPUT96), .ZN(new_n573));
  AOI21_X1  g387(.A(KEYINPUT96), .B1(new_n567), .B2(new_n572), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n518), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(G113), .B(G122), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(new_n398), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n340), .A2(G143), .A3(G214), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(G143), .B1(new_n340), .B2(G214), .ZN(new_n580));
  OAI21_X1  g394(.A(G131), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n340), .A2(G214), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n265), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n583), .A2(new_n260), .A3(new_n578), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n194), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n208), .B(KEYINPUT19), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n586), .B1(new_n192), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n577), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT90), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n583), .A2(new_n590), .A3(new_n578), .ZN(new_n591));
  NAND2_X1  g405(.A1(KEYINPUT18), .A2(G131), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n583), .A2(new_n590), .A3(new_n578), .A4(new_n592), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n189), .A2(G146), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n209), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(KEYINPUT89), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT89), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n596), .A2(new_n209), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n594), .A2(new_n595), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n589), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(G475), .A2(G902), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT17), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n581), .A2(new_n605), .A3(new_n584), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n260), .B1(new_n583), .B2(new_n578), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n195), .B1(new_n607), .B2(KEYINPUT17), .ZN(new_n608));
  AOI22_X1  g422(.A1(new_n591), .A2(new_n593), .B1(new_n598), .B2(new_n600), .ZN(new_n609));
  AOI22_X1  g423(.A1(new_n606), .A2(new_n608), .B1(new_n609), .B2(new_n595), .ZN(new_n610));
  INV_X1    g424(.A(new_n577), .ZN(new_n611));
  OAI211_X1 g425(.A(new_n603), .B(new_n604), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(KEYINPUT20), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT91), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n612), .A2(KEYINPUT91), .A3(KEYINPUT20), .ZN(new_n616));
  INV_X1    g430(.A(new_n606), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n193), .B(new_n194), .C1(new_n581), .C2(new_n605), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n602), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AOI22_X1  g433(.A1(new_n619), .A2(new_n577), .B1(new_n602), .B2(new_n589), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT20), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n620), .A2(new_n621), .A3(new_n604), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n615), .A2(new_n616), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n611), .A2(KEYINPUT92), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n228), .B1(new_n619), .B2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n624), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n610), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(G475), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n575), .A2(new_n629), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n470), .A2(new_n512), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n395), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G101), .ZN(G3));
  NOR2_X1   g447(.A1(new_n511), .A2(new_n241), .ZN(new_n634));
  OAI21_X1  g448(.A(G472), .B1(new_n387), .B2(G902), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n634), .A2(new_n388), .A3(new_n393), .A4(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n558), .A2(new_n228), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n639), .B1(new_n557), .B2(G478), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n546), .A2(new_n556), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT33), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n640), .B1(new_n642), .B2(G478), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n629), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n469), .B1(new_n463), .B2(new_n464), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n518), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n644), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n637), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(new_n398), .ZN(new_n650));
  XNOR2_X1  g464(.A(KEYINPUT98), .B(KEYINPUT34), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G6));
  INV_X1    g466(.A(KEYINPUT101), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT100), .ZN(new_n654));
  OAI211_X1 g468(.A(new_n654), .B(G475), .C1(new_n625), .C2(new_n627), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(G902), .B1(new_n610), .B2(new_n626), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n619), .A2(new_n624), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n654), .B1(new_n659), .B2(G475), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT99), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n620), .A2(new_n662), .A3(new_n621), .A4(new_n604), .ZN(new_n663));
  OAI21_X1  g477(.A(KEYINPUT99), .B1(new_n612), .B2(KEYINPUT20), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n615), .A2(new_n616), .A3(new_n663), .A4(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n567), .A2(new_n572), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT96), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n567), .A2(new_n572), .A3(KEYINPUT96), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n661), .A2(new_n665), .A3(new_n668), .A4(new_n669), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n653), .B1(new_n670), .B2(new_n647), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n628), .A2(KEYINPUT100), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n655), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n673), .A2(new_n573), .A3(new_n574), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n674), .A2(KEYINPUT101), .A3(new_n518), .A4(new_n665), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n671), .A2(new_n675), .A3(new_n645), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n637), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT102), .ZN(new_n678));
  XNOR2_X1  g492(.A(KEYINPUT35), .B(G107), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G9));
  NOR2_X1   g494(.A1(new_n222), .A2(KEYINPUT36), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n214), .B(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  OAI22_X1  g497(.A1(new_n239), .A2(new_n240), .B1(new_n231), .B2(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n470), .A2(new_n630), .A3(new_n512), .A4(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n388), .A2(new_n635), .A3(new_n393), .ZN(new_n686));
  OR2_X1    g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT37), .B(G110), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G12));
  NAND2_X1  g503(.A1(new_n385), .A2(new_n394), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n492), .A2(new_n501), .ZN(new_n691));
  INV_X1    g505(.A(G469), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n691), .A2(new_n692), .A3(new_n228), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n693), .A2(new_n509), .A3(new_n508), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n694), .A2(new_n684), .A3(new_n645), .A4(new_n472), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n573), .A2(new_n574), .ZN(new_n696));
  OR2_X1    g510(.A1(new_n516), .A2(G900), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n514), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n696), .A2(new_n665), .A3(new_n661), .A4(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n690), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G128), .ZN(G30));
  XNOR2_X1  g516(.A(new_n698), .B(KEYINPUT39), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n512), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g518(.A(new_n704), .B(KEYINPUT40), .Z(new_n705));
  XOR2_X1   g519(.A(new_n467), .B(KEYINPUT38), .Z(new_n706));
  INV_X1    g520(.A(new_n684), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n345), .B1(new_n321), .B2(new_n334), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n321), .A2(new_n367), .ZN(new_n710));
  OAI211_X1 g524(.A(new_n709), .B(KEYINPUT103), .C1(new_n344), .C2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT103), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n710), .A2(new_n344), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n712), .B1(new_n713), .B2(new_n708), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n711), .A2(new_n714), .A3(new_n228), .ZN(new_n715));
  AOI22_X1  g529(.A1(G472), .A2(new_n715), .B1(new_n384), .B2(KEYINPUT32), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n394), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n696), .A2(new_n629), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n718), .A2(new_n468), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n706), .A2(new_n707), .A3(new_n717), .A4(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT104), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n705), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n720), .A2(new_n721), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(new_n265), .ZN(G45));
  NAND3_X1  g539(.A1(new_n629), .A2(new_n643), .A3(new_n698), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n695), .A2(new_n726), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n690), .A2(new_n727), .ZN(new_n728));
  XOR2_X1   g542(.A(KEYINPUT105), .B(G146), .Z(new_n729));
  XNOR2_X1  g543(.A(new_n728), .B(new_n729), .ZN(G48));
  AOI21_X1  g544(.A(new_n692), .B1(new_n691), .B2(new_n228), .ZN(new_n731));
  INV_X1    g545(.A(new_n472), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n731), .A2(new_n502), .A3(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n395), .A2(new_n648), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(KEYINPUT41), .B(G113), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G15));
  NAND3_X1  g550(.A1(new_n676), .A2(new_n395), .A3(new_n733), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G116), .ZN(G18));
  NAND2_X1  g552(.A1(new_n733), .A2(new_n645), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n690), .A2(new_n630), .A3(new_n684), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G119), .ZN(G21));
  NAND4_X1  g556(.A1(new_n718), .A2(new_n518), .A3(new_n645), .A4(new_n733), .ZN(new_n743));
  INV_X1    g557(.A(new_n241), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n383), .B1(new_n369), .B2(new_n344), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n390), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n744), .A2(new_n635), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(KEYINPUT106), .B1(new_n743), .B2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n696), .A2(new_n629), .A3(new_n518), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n739), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n747), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT106), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n748), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G122), .ZN(G24));
  AND3_X1   g569(.A1(new_n635), .A2(new_n684), .A3(new_n746), .ZN(new_n756));
  INV_X1    g570(.A(new_n726), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n740), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G125), .ZN(G27));
  OAI21_X1  g573(.A(new_n389), .B1(new_n387), .B2(new_n374), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n241), .B1(new_n385), .B2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT107), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n511), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n694), .A2(KEYINPUT107), .A3(new_n472), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n469), .B1(new_n465), .B2(new_n466), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n761), .A2(new_n766), .A3(KEYINPUT42), .A4(new_n757), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n766), .A2(new_n690), .A3(new_n744), .A4(new_n757), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT108), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT42), .ZN(new_n770));
  AND3_X1   g584(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n769), .B1(new_n768), .B2(new_n770), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n767), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  XOR2_X1   g587(.A(KEYINPUT109), .B(G131), .Z(new_n774));
  XNOR2_X1  g588(.A(new_n773), .B(new_n774), .ZN(G33));
  INV_X1    g589(.A(new_n699), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n395), .A2(new_n776), .A3(new_n766), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G134), .ZN(G36));
  AND2_X1   g592(.A1(new_n504), .A2(new_n507), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n779), .A2(KEYINPUT45), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(KEYINPUT45), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(G469), .A3(new_n781), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n782), .A2(new_n509), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(KEYINPUT46), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n784), .B(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT111), .ZN(new_n787));
  OR3_X1    g601(.A1(new_n783), .A2(new_n787), .A3(KEYINPUT46), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n787), .B1(new_n783), .B2(KEYINPUT46), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n786), .A2(new_n693), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT112), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n790), .A2(new_n791), .A3(new_n472), .A4(new_n703), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n784), .B(KEYINPUT110), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n788), .A2(new_n693), .A3(new_n789), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n472), .B(new_n703), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(KEYINPUT112), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n623), .A2(new_n628), .A3(new_n643), .ZN(new_n798));
  XOR2_X1   g612(.A(new_n798), .B(KEYINPUT43), .Z(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(new_n686), .A3(new_n684), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT44), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n765), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n802), .A2(KEYINPUT113), .A3(new_n765), .ZN(new_n806));
  AOI22_X1  g620(.A1(new_n805), .A2(new_n806), .B1(new_n801), .B2(new_n800), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n797), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(KEYINPUT114), .B(G137), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n808), .B(new_n809), .ZN(G39));
  NAND3_X1  g624(.A1(new_n790), .A2(KEYINPUT47), .A3(new_n472), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n472), .B1(new_n793), .B2(new_n794), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT47), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n467), .A2(new_n468), .ZN(new_n816));
  NOR4_X1   g630(.A1(new_n690), .A2(new_n744), .A3(new_n726), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G140), .ZN(G42));
  NOR2_X1   g633(.A1(new_n731), .A2(new_n502), .ZN(new_n820));
  XOR2_X1   g634(.A(new_n820), .B(KEYINPUT49), .Z(new_n821));
  OR4_X1    g635(.A1(new_n241), .A2(new_n798), .A3(new_n469), .A4(new_n732), .ZN(new_n822));
  OR4_X1    g636(.A1(new_n717), .A2(new_n706), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n514), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n799), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n820), .A2(new_n472), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n816), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n825), .A2(new_n761), .A3(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(KEYINPUT48), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n218), .A2(G952), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n825), .A2(new_n751), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n830), .B1(new_n831), .B2(new_n740), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n827), .A2(new_n744), .A3(new_n824), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n833), .A2(new_n717), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT123), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n829), .B(new_n832), .C1(new_n644), .C2(new_n835), .ZN(new_n836));
  OR3_X1    g650(.A1(new_n835), .A2(new_n629), .A3(new_n643), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n706), .A2(new_n468), .A3(new_n826), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n831), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT50), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n825), .A2(new_n756), .A3(new_n827), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n837), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT51), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n820), .A2(new_n732), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n811), .A2(new_n814), .A3(new_n846), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n831), .A2(new_n765), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n836), .B1(new_n845), .B2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT122), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n847), .A2(new_n851), .A3(new_n848), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n851), .B1(new_n847), .B2(new_n848), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n852), .A2(new_n853), .A3(new_n843), .ZN(new_n854));
  XNOR2_X1  g668(.A(KEYINPUT121), .B(KEYINPUT51), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n850), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n395), .A2(new_n631), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n623), .A2(new_n628), .A3(new_n666), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n644), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n860), .A2(new_n470), .A3(new_n518), .ZN(new_n861));
  OAI22_X1  g675(.A1(new_n861), .A2(new_n636), .B1(new_n685), .B2(new_n686), .ZN(new_n862));
  OAI21_X1  g676(.A(KEYINPUT115), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  OR2_X1    g677(.A1(new_n636), .A2(new_n861), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT115), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n864), .A2(new_n687), .A3(new_n865), .A4(new_n632), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  AND4_X1   g681(.A1(new_n734), .A2(new_n754), .A3(new_n737), .A4(new_n741), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n766), .A2(new_n757), .A3(new_n756), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n777), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(new_n698), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n666), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n661), .A2(new_n665), .A3(new_n872), .ZN(new_n873));
  NOR4_X1   g687(.A1(new_n816), .A2(new_n511), .A3(new_n707), .A4(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT116), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n874), .A2(new_n690), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n874), .A2(new_n690), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT116), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n870), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n773), .A2(new_n867), .A3(new_n868), .A4(new_n879), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n718), .A2(new_n645), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n511), .A2(new_n871), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n717), .A2(new_n881), .A3(new_n882), .A4(new_n707), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n690), .B1(new_n700), .B2(new_n727), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n883), .A2(new_n884), .A3(new_n758), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT52), .B1(new_n885), .B2(KEYINPUT117), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n885), .A2(KEYINPUT117), .A3(KEYINPUT52), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OAI211_X1 g703(.A(KEYINPUT118), .B(new_n857), .C1(new_n880), .C2(new_n889), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n867), .A2(new_n868), .A3(new_n879), .ZN(new_n891));
  XOR2_X1   g705(.A(KEYINPUT119), .B(KEYINPUT53), .Z(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n885), .B(KEYINPUT52), .Z(new_n894));
  NAND4_X1  g708(.A1(new_n891), .A2(new_n773), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n890), .A2(new_n895), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n885), .A2(KEYINPUT117), .A3(KEYINPUT52), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n897), .A2(new_n886), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n754), .A2(new_n737), .A3(new_n734), .A4(new_n741), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n863), .B2(new_n866), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n898), .A2(new_n900), .A3(new_n773), .A4(new_n879), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT118), .B1(new_n901), .B2(new_n857), .ZN(new_n902));
  OAI21_X1  g716(.A(KEYINPUT54), .B1(new_n896), .B2(new_n902), .ZN(new_n903));
  OR2_X1    g717(.A1(new_n901), .A2(new_n857), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT54), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n891), .A2(new_n773), .A3(new_n894), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n892), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n904), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n903), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT120), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT120), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n903), .A2(new_n911), .A3(new_n908), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n856), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(G952), .A2(G953), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n823), .B1(new_n913), .B2(new_n914), .ZN(G75));
  NOR2_X1   g729(.A1(new_n218), .A2(G952), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n228), .B1(new_n904), .B2(new_n907), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT56), .B1(new_n918), .B2(G210), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n431), .A2(new_n433), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT124), .Z(new_n921));
  XNOR2_X1  g735(.A(new_n441), .B(KEYINPUT55), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n921), .B(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n917), .B1(new_n919), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n924), .B1(new_n919), .B2(new_n923), .ZN(G51));
  XOR2_X1   g739(.A(new_n691), .B(KEYINPUT125), .Z(new_n926));
  INV_X1    g740(.A(new_n908), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n905), .B1(new_n904), .B2(new_n907), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n509), .B(KEYINPUT57), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n926), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n904), .A2(new_n907), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(G902), .ZN(new_n933));
  OR2_X1    g747(.A1(new_n933), .A2(new_n782), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n916), .B1(new_n931), .B2(new_n934), .ZN(G54));
  AND3_X1   g749(.A1(new_n918), .A2(KEYINPUT58), .A3(G475), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n936), .A2(new_n620), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n917), .B1(new_n936), .B2(new_n620), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n937), .A2(new_n938), .ZN(G60));
  XNOR2_X1  g753(.A(new_n638), .B(KEYINPUT59), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n642), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n917), .B1(new_n929), .B2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n940), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n910), .A2(new_n912), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n942), .B1(new_n944), .B2(new_n642), .ZN(G63));
  INV_X1    g759(.A(KEYINPUT61), .ZN(new_n946));
  NAND2_X1  g760(.A1(G217), .A2(G902), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT60), .Z(new_n948));
  NAND2_X1  g762(.A1(new_n932), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n226), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n917), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n949), .A2(new_n683), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n946), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n932), .A2(new_n682), .A3(new_n948), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n950), .A2(KEYINPUT61), .A3(new_n917), .A4(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n953), .A2(new_n955), .ZN(G66));
  AOI21_X1  g770(.A(new_n218), .B1(new_n515), .B2(G224), .ZN(new_n957));
  INV_X1    g771(.A(new_n900), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n957), .B1(new_n958), .B2(new_n218), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n921), .B1(G898), .B2(new_n218), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT126), .Z(new_n961));
  XNOR2_X1  g775(.A(new_n959), .B(new_n961), .ZN(G69));
  NAND2_X1  g776(.A1(new_n322), .A2(new_n333), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(new_n587), .Z(new_n964));
  INV_X1    g778(.A(G900), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n964), .B1(new_n965), .B2(new_n218), .ZN(new_n966));
  AOI22_X1  g780(.A1(new_n797), .A2(new_n807), .B1(new_n815), .B2(new_n817), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n797), .A2(new_n761), .A3(new_n881), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n884), .A2(new_n758), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n773), .A2(new_n777), .A3(new_n969), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n967), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n966), .B1(new_n971), .B2(new_n218), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n218), .B1(G227), .B2(G900), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n969), .B1(new_n722), .B2(new_n723), .ZN(new_n974));
  OR2_X1    g788(.A1(new_n974), .A2(KEYINPUT62), .ZN(new_n975));
  AOI211_X1 g789(.A(new_n816), .B(new_n704), .C1(new_n644), .C2(new_n859), .ZN(new_n976));
  AOI22_X1  g790(.A1(new_n974), .A2(KEYINPUT62), .B1(new_n395), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n967), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n964), .B1(new_n978), .B2(new_n218), .ZN(new_n979));
  OR3_X1    g793(.A1(new_n972), .A2(new_n973), .A3(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n973), .B1(new_n972), .B2(new_n979), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(G72));
  NAND3_X1  g796(.A1(new_n321), .A2(new_n345), .A3(new_n334), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n967), .A2(new_n900), .A3(new_n968), .A4(new_n970), .ZN(new_n984));
  NAND2_X1  g798(.A1(G472), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT63), .Z(new_n986));
  AOI21_X1  g800(.A(new_n983), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n967), .A2(new_n900), .A3(new_n975), .A4(new_n977), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n709), .B1(new_n988), .B2(new_n986), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n987), .A2(new_n989), .A3(new_n916), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT127), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n346), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n346), .A2(new_n991), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n993), .B1(new_n379), .B2(new_n380), .ZN(new_n994));
  OAI221_X1 g808(.A(new_n986), .B1(new_n992), .B2(new_n994), .C1(new_n896), .C2(new_n902), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n990), .A2(new_n995), .ZN(G57));
endmodule


