//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 1 1 1 1 0 0 0 0 1 1 1 1 1 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957;
  INV_X1    g000(.A(G475), .ZN(new_n187));
  INV_X1    g001(.A(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  AND3_X1   g003(.A1(new_n188), .A2(new_n189), .A3(G214), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT88), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n188), .A2(new_n189), .A3(G214), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT88), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n191), .A2(new_n192), .A3(new_n195), .ZN(new_n196));
  OR2_X1    g010(.A1(new_n196), .A2(KEYINPUT89), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n190), .A2(G143), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(KEYINPUT89), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n197), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G131), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT17), .ZN(new_n202));
  INV_X1    g016(.A(G131), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n197), .A2(new_n203), .A3(new_n198), .A4(new_n199), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n201), .A2(new_n202), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G140), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G125), .ZN(new_n207));
  INV_X1    g021(.A(G125), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G140), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n207), .A2(new_n209), .A3(KEYINPUT79), .A4(KEYINPUT16), .ZN(new_n210));
  AND3_X1   g024(.A1(new_n207), .A2(new_n209), .A3(KEYINPUT16), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT79), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n212), .B1(new_n207), .B2(KEYINPUT16), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n210), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G146), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G146), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n217), .B(new_n210), .C1(new_n211), .C2(new_n213), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n200), .A2(KEYINPUT17), .A3(G131), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n205), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT18), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n200), .B1(new_n223), .B2(new_n203), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n203), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n197), .A2(new_n225), .A3(new_n198), .A4(new_n199), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n207), .A2(new_n209), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n228), .A2(G146), .ZN(new_n229));
  OR2_X1    g043(.A1(new_n229), .A2(KEYINPUT90), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(G146), .ZN(new_n231));
  XOR2_X1   g045(.A(new_n230), .B(new_n231), .Z(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n227), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n222), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(G113), .B(G122), .ZN(new_n236));
  INV_X1    g050(.A(G104), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n236), .B(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n222), .A2(new_n234), .A3(new_n238), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G902), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n187), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n232), .B1(new_n224), .B2(new_n226), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n228), .B(KEYINPUT19), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n215), .B1(new_n246), .B2(G146), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n247), .B1(new_n201), .B2(new_n204), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n239), .B1(new_n245), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n241), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT91), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT20), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(G475), .B1(new_n241), .B2(new_n249), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(new_n243), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n251), .A2(new_n252), .A3(new_n243), .A4(new_n254), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n244), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G116), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(KEYINPUT14), .A3(G122), .ZN(new_n261));
  XNOR2_X1  g075(.A(G116), .B(G122), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  OAI211_X1 g077(.A(G107), .B(new_n261), .C1(new_n263), .C2(KEYINPUT14), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n264), .B(KEYINPUT94), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n192), .A2(G128), .ZN(new_n266));
  INV_X1    g080(.A(G128), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n267), .A2(G143), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G134), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n269), .B(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G107), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n262), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n273), .B(KEYINPUT93), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n265), .A2(new_n271), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n268), .A2(KEYINPUT13), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n276), .B(KEYINPUT92), .ZN(new_n277));
  INV_X1    g091(.A(new_n266), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n278), .B1(new_n268), .B2(KEYINPUT13), .ZN(new_n279));
  OAI21_X1  g093(.A(G134), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n269), .A2(new_n270), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n262), .B(new_n272), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  XOR2_X1   g097(.A(KEYINPUT9), .B(G234), .Z(new_n284));
  NAND3_X1  g098(.A1(new_n284), .A2(G217), .A3(new_n189), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  AND3_X1   g100(.A1(new_n275), .A2(new_n283), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n286), .B1(new_n275), .B2(new_n283), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n243), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT95), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G478), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n292), .A2(KEYINPUT15), .ZN(new_n293));
  OAI211_X1 g107(.A(KEYINPUT95), .B(new_n243), .C1(new_n287), .C2(new_n288), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n291), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT96), .ZN(new_n296));
  OR3_X1    g110(.A1(new_n289), .A2(new_n296), .A3(new_n293), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n296), .B1(new_n289), .B2(new_n293), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n295), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n189), .A2(G952), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n300), .B1(G234), .B2(G237), .ZN(new_n301));
  XOR2_X1   g115(.A(KEYINPUT21), .B(G898), .Z(new_n302));
  XNOR2_X1  g116(.A(new_n302), .B(KEYINPUT97), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  AOI211_X1 g118(.A(new_n243), .B(new_n189), .C1(G234), .C2(G237), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n301), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NOR3_X1   g120(.A1(new_n259), .A2(new_n299), .A3(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(KEYINPUT3), .B1(new_n237), .B2(G107), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT3), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(new_n272), .A3(G104), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n237), .A2(G107), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n308), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  OR2_X1    g126(.A1(new_n312), .A2(G101), .ZN(new_n313));
  INV_X1    g127(.A(new_n311), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n237), .A2(G107), .ZN(new_n315));
  OAI21_X1  g129(.A(G101), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  AND2_X1   g130(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n192), .B(G146), .C1(new_n267), .C2(KEYINPUT1), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n267), .A2(new_n217), .A3(G143), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OR2_X1    g134(.A1(new_n320), .A2(KEYINPUT85), .ZN(new_n321));
  XNOR2_X1  g135(.A(G143), .B(G146), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT1), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(new_n323), .A3(G128), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n320), .A2(KEYINPUT85), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n321), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n317), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n320), .A2(KEYINPUT67), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT67), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n318), .A2(new_n329), .A3(new_n319), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(new_n324), .A3(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n327), .B1(new_n331), .B2(new_n317), .ZN(new_n332));
  OAI21_X1  g146(.A(KEYINPUT66), .B1(new_n270), .B2(G137), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT11), .ZN(new_n334));
  INV_X1    g148(.A(G137), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n335), .A2(G134), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT11), .ZN(new_n338));
  OAI211_X1 g152(.A(KEYINPUT66), .B(new_n338), .C1(new_n270), .C2(G137), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n334), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G131), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n334), .A2(new_n203), .A3(new_n337), .A4(new_n339), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n332), .A2(KEYINPUT12), .A3(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT86), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT68), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n341), .A2(KEYINPUT68), .A3(new_n342), .ZN(new_n349));
  AND2_X1   g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n332), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT12), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n332), .A2(KEYINPUT86), .A3(KEYINPUT12), .A4(new_n343), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n346), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n327), .A2(new_n356), .ZN(new_n357));
  AND2_X1   g171(.A1(KEYINPUT0), .A2(G128), .ZN(new_n358));
  NOR2_X1   g172(.A1(KEYINPUT0), .A2(G128), .ZN(new_n359));
  NOR3_X1   g173(.A1(new_n322), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(KEYINPUT65), .B1(new_n322), .B2(new_n358), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NOR4_X1   g176(.A1(new_n322), .A2(KEYINPUT65), .A3(new_n358), .A4(new_n359), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT4), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n312), .A2(new_n365), .A3(G101), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n312), .A2(G101), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n313), .A2(new_n367), .A3(KEYINPUT4), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n364), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n317), .A2(KEYINPUT10), .A3(new_n331), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n357), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n371), .A2(new_n350), .ZN(new_n372));
  XNOR2_X1  g186(.A(G110), .B(G140), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n189), .A2(G227), .ZN(new_n374));
  XOR2_X1   g188(.A(new_n373), .B(new_n374), .Z(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n372), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n355), .A2(new_n377), .ZN(new_n378));
  OR2_X1    g192(.A1(new_n371), .A2(new_n350), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n371), .A2(new_n350), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n378), .B1(new_n381), .B2(new_n375), .ZN(new_n382));
  INV_X1    g196(.A(G469), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n383), .A3(new_n243), .ZN(new_n384));
  NAND2_X1  g198(.A1(G469), .A2(G902), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT87), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n379), .A2(new_n386), .A3(new_n375), .ZN(new_n387));
  OAI21_X1  g201(.A(KEYINPUT87), .B1(new_n372), .B2(new_n376), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n380), .A3(new_n388), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n355), .A2(new_n379), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n389), .B(G469), .C1(new_n390), .C2(new_n375), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n384), .A2(new_n385), .A3(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(G214), .B1(G237), .B2(G902), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n364), .A2(G125), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n331), .A2(new_n208), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G224), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(G953), .ZN(new_n399));
  OR2_X1    g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n397), .A2(new_n399), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n400), .B(new_n401), .C1(KEYINPUT7), .C2(new_n399), .ZN(new_n402));
  XOR2_X1   g216(.A(G116), .B(G119), .Z(new_n403));
  XNOR2_X1  g217(.A(KEYINPUT2), .B(G113), .ZN(new_n404));
  XOR2_X1   g218(.A(new_n403), .B(new_n404), .Z(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(new_n366), .A3(new_n368), .ZN(new_n407));
  XOR2_X1   g221(.A(G110), .B(G122), .Z(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT5), .ZN(new_n410));
  INV_X1    g224(.A(G119), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(new_n411), .A3(G116), .ZN(new_n412));
  OAI211_X1 g226(.A(G113), .B(new_n412), .C1(new_n403), .C2(new_n410), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n413), .B1(new_n403), .B2(new_n404), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n313), .A2(new_n316), .ZN(new_n415));
  OR2_X1    g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n407), .A2(new_n409), .A3(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n414), .B(new_n415), .ZN(new_n418));
  XOR2_X1   g232(.A(new_n408), .B(KEYINPUT8), .Z(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OR3_X1    g234(.A1(new_n397), .A2(KEYINPUT7), .A3(new_n399), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n402), .A2(new_n417), .A3(new_n420), .A4(new_n421), .ZN(new_n422));
  AND2_X1   g236(.A1(new_n400), .A2(new_n401), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n407), .A2(new_n416), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT6), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(new_n425), .A3(new_n408), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n424), .A2(new_n408), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(KEYINPUT6), .A3(new_n417), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n423), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n422), .A2(new_n243), .A3(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(G210), .B1(G237), .B2(G902), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n422), .A2(new_n243), .A3(new_n429), .A4(new_n431), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n394), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n284), .ZN(new_n436));
  OAI21_X1  g250(.A(G221), .B1(new_n436), .B2(G902), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n437), .B(KEYINPUT84), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n392), .A2(new_n435), .A3(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n307), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT83), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n215), .A2(new_n218), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT77), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n445), .B(KEYINPUT23), .C1(new_n267), .C2(G119), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n411), .A2(KEYINPUT77), .A3(G128), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(KEYINPUT78), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n267), .A2(G119), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT78), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n445), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT23), .ZN(new_n452));
  AOI22_X1  g266(.A1(new_n448), .A2(new_n449), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(G110), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT76), .ZN(new_n455));
  NOR3_X1   g269(.A1(new_n455), .A2(new_n267), .A3(G119), .ZN(new_n456));
  AOI21_X1  g270(.A(KEYINPUT76), .B1(new_n411), .B2(G128), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n449), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(KEYINPUT24), .B(G110), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n444), .B(new_n454), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT81), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n458), .A2(new_n459), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n462), .B1(new_n453), .B2(G110), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT80), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n229), .B1(new_n214), .B2(G146), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n464), .B1(new_n463), .B2(new_n465), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n460), .B(new_n461), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n469), .B(KEYINPUT22), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(new_n335), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n463), .A2(new_n465), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT80), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n463), .A2(new_n465), .A3(new_n464), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n461), .B1(new_n476), .B2(new_n460), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n460), .B1(new_n466), .B2(new_n467), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT81), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n480), .A2(new_n468), .A3(new_n471), .ZN(new_n481));
  AOI21_X1  g295(.A(G902), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n483));
  NAND2_X1  g297(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NOR3_X1   g299(.A1(new_n482), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n472), .A2(new_n477), .ZN(new_n487));
  AOI211_X1 g301(.A(new_n461), .B(new_n471), .C1(new_n476), .C2(new_n460), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n243), .B(new_n483), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(G234), .ZN(new_n490));
  OAI21_X1  g304(.A(G217), .B1(new_n490), .B2(G902), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(KEYINPUT75), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n443), .B1(new_n486), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n478), .A2(new_n481), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n243), .ZN(new_n496));
  INV_X1    g310(.A(new_n483), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n497), .A3(new_n484), .ZN(new_n498));
  INV_X1    g312(.A(new_n492), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n499), .B1(new_n482), .B2(new_n483), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n498), .A2(new_n500), .A3(KEYINPUT83), .ZN(new_n501));
  AOI21_X1  g315(.A(G902), .B1(new_n490), .B2(G217), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n495), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n494), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT32), .ZN(new_n505));
  NOR2_X1   g319(.A1(G472), .A2(G902), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(G101), .ZN(new_n509));
  INV_X1    g323(.A(G210), .ZN(new_n510));
  NOR3_X1   g324(.A1(new_n510), .A2(G237), .A3(G953), .ZN(new_n511));
  XOR2_X1   g325(.A(new_n509), .B(new_n511), .Z(new_n512));
  NAND3_X1  g326(.A1(new_n348), .A2(new_n349), .A3(new_n364), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n270), .A2(G137), .ZN(new_n514));
  OAI21_X1  g328(.A(G131), .B1(new_n336), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n331), .A2(new_n342), .A3(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n513), .A2(new_n405), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT69), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT69), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n513), .A2(new_n519), .A3(new_n405), .A4(new_n516), .ZN(new_n520));
  OR2_X1    g334(.A1(new_n360), .A2(new_n361), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT65), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n360), .A2(new_n522), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n343), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n516), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n406), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n518), .A2(new_n520), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT28), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT28), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n517), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n512), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  AND2_X1   g345(.A1(new_n518), .A2(new_n520), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n513), .A2(KEYINPUT30), .A3(new_n516), .ZN(new_n533));
  XOR2_X1   g347(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n534));
  OAI21_X1  g348(.A(new_n534), .B1(new_n524), .B2(new_n525), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n533), .A2(new_n535), .A3(new_n406), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n532), .A2(KEYINPUT70), .A3(new_n512), .A4(new_n536), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n536), .A2(new_n518), .A3(new_n520), .A4(new_n512), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT70), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n531), .B1(new_n541), .B2(KEYINPUT31), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n536), .A2(new_n518), .A3(new_n520), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT31), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n543), .A2(KEYINPUT71), .A3(new_n544), .A4(new_n512), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT71), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n546), .B1(new_n538), .B2(KEYINPUT31), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n507), .B1(new_n542), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT72), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n505), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n538), .A2(new_n539), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n538), .A2(new_n539), .ZN(new_n553));
  OAI21_X1  g367(.A(KEYINPUT31), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n531), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(new_n548), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n506), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n557), .A2(KEYINPUT72), .A3(KEYINPUT32), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n551), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n530), .ZN(new_n560));
  INV_X1    g374(.A(new_n512), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT29), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n518), .A2(new_n520), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT73), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n513), .A2(new_n516), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n406), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n518), .A2(KEYINPUT73), .A3(new_n520), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n567), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AOI211_X1 g385(.A(new_n560), .B(new_n564), .C1(new_n571), .C2(KEYINPUT28), .ZN(new_n572));
  OAI21_X1  g386(.A(KEYINPUT74), .B1(new_n572), .B2(G902), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(KEYINPUT28), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n574), .A2(new_n530), .A3(new_n563), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT74), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(new_n576), .A3(new_n243), .ZN(new_n577));
  INV_X1    g391(.A(new_n543), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n561), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n528), .A2(new_n530), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n579), .B(new_n562), .C1(new_n580), .C2(new_n561), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n573), .A2(new_n577), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(G472), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n504), .B1(new_n559), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n442), .A2(new_n584), .ZN(new_n585));
  XOR2_X1   g399(.A(KEYINPUT98), .B(G101), .Z(new_n586));
  XNOR2_X1  g400(.A(new_n585), .B(new_n586), .ZN(G3));
  INV_X1    g401(.A(new_n504), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n392), .A2(new_n439), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(G472), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n591), .B1(new_n556), .B2(new_n243), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n592), .A2(new_n549), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n291), .A2(new_n292), .A3(new_n294), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT99), .B1(new_n287), .B2(new_n288), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(KEYINPUT33), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT33), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(G902), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n597), .B1(new_n603), .B2(G478), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n258), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n306), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n435), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(KEYINPUT100), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT100), .ZN(new_n610));
  NOR4_X1   g424(.A1(new_n607), .A2(new_n258), .A3(new_n604), .A4(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n595), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT34), .B(G104), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G6));
  XNOR2_X1  g429(.A(new_n255), .B(KEYINPUT20), .ZN(new_n616));
  INV_X1    g430(.A(new_n244), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AND3_X1   g432(.A1(new_n618), .A2(new_n299), .A3(new_n608), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n595), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT35), .B(G107), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G9));
  NOR2_X1   g436(.A1(new_n471), .A2(KEYINPUT36), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n479), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n502), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(KEYINPUT101), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n494), .A2(new_n501), .A3(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT102), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n442), .A2(new_n593), .A3(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT37), .B(G110), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT103), .B(KEYINPUT104), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G12));
  NAND2_X1  g448(.A1(new_n559), .A2(new_n583), .ZN(new_n635));
  INV_X1    g449(.A(G900), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n301), .B1(new_n305), .B2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n616), .A2(new_n299), .A3(new_n617), .A4(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n440), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n635), .A2(new_n629), .A3(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT105), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n635), .A2(KEYINPUT105), .A3(new_n629), .A4(new_n640), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G128), .ZN(G30));
  AOI22_X1  g460(.A1(new_n571), .A2(new_n561), .B1(new_n537), .B2(new_n540), .ZN(new_n647));
  OAI21_X1  g461(.A(G472), .B1(new_n647), .B2(G902), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n559), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n637), .B(KEYINPUT39), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n589), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n650), .B1(KEYINPUT40), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n653), .A2(KEYINPUT40), .ZN(new_n655));
  INV_X1    g469(.A(new_n299), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n258), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n433), .A2(new_n434), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT38), .ZN(new_n661));
  INV_X1    g475(.A(new_n627), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n654), .A2(new_n393), .A3(new_n659), .A4(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G143), .ZN(G45));
  NAND2_X1  g479(.A1(new_n605), .A2(new_n638), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n635), .A2(new_n441), .A3(new_n629), .A4(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G146), .ZN(G48));
  NAND2_X1  g483(.A1(new_n382), .A2(new_n243), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(G469), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n671), .A2(new_n384), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n439), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n612), .A2(new_n584), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT41), .B(G113), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G15));
  NAND3_X1  g491(.A1(new_n584), .A2(new_n619), .A3(new_n674), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G116), .ZN(G18));
  INV_X1    g493(.A(new_n435), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n673), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n635), .A2(new_n307), .A3(new_n629), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G119), .ZN(G21));
  AOI21_X1  g497(.A(new_n560), .B1(new_n571), .B2(KEYINPUT28), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n554), .B1(new_n684), .B2(new_n512), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT106), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  OAI211_X1 g501(.A(new_n554), .B(KEYINPUT106), .C1(new_n684), .C2(new_n512), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n687), .A2(new_n548), .A3(new_n688), .ZN(new_n689));
  AOI211_X1 g503(.A(new_n504), .B(new_n592), .C1(new_n689), .C2(new_n506), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n690), .A2(new_n608), .A3(new_n657), .A4(new_n674), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G122), .ZN(G24));
  AOI21_X1  g506(.A(new_n592), .B1(new_n689), .B2(new_n506), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n667), .A2(new_n693), .A3(new_n681), .A4(new_n627), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G125), .ZN(G27));
  NAND3_X1  g509(.A1(new_n433), .A2(new_n393), .A3(new_n434), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n385), .B(KEYINPUT107), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n384), .A2(new_n391), .A3(new_n698), .ZN(new_n699));
  AND3_X1   g513(.A1(new_n697), .A2(new_n439), .A3(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n635), .A2(new_n588), .A3(new_n667), .A4(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(KEYINPUT108), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT42), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n584), .A2(new_n704), .A3(new_n667), .A4(new_n700), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n557), .A2(new_n505), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n549), .A2(KEYINPUT32), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n583), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  AND2_X1   g523(.A1(new_n709), .A2(new_n588), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n667), .A2(new_n700), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n710), .A2(KEYINPUT42), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n706), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G131), .ZN(G33));
  INV_X1    g528(.A(new_n639), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n584), .A2(new_n715), .A3(new_n700), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G134), .ZN(G36));
  INV_X1    g531(.A(new_n604), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n258), .A2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT43), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(KEYINPUT109), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n719), .B(KEYINPUT43), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT109), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT110), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n727), .B1(new_n593), .B2(new_n662), .ZN(new_n728));
  OAI211_X1 g542(.A(KEYINPUT110), .B(new_n627), .C1(new_n592), .C2(new_n549), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n726), .A2(KEYINPUT44), .A3(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AOI22_X1  g547(.A1(new_n722), .A2(new_n725), .B1(new_n728), .B2(new_n729), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(KEYINPUT111), .A3(KEYINPUT44), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n389), .B1(new_n390), .B2(new_n375), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT45), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n737), .A2(new_n738), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n739), .A2(G469), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n698), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT46), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n741), .A2(KEYINPUT46), .A3(new_n698), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n744), .A2(new_n384), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n439), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n747), .A2(new_n651), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n734), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT44), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n736), .A2(new_n697), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G137), .ZN(G39));
  INV_X1    g568(.A(KEYINPUT47), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(KEYINPUT112), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n747), .A2(new_n756), .ZN(new_n757));
  AOI22_X1  g571(.A1(new_n746), .A2(new_n439), .B1(KEYINPUT112), .B2(new_n755), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n757), .B1(new_n758), .B2(new_n756), .ZN(new_n759));
  NOR4_X1   g573(.A1(new_n635), .A2(new_n666), .A3(new_n588), .A4(new_n696), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT113), .ZN(new_n761));
  OR2_X1    g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n759), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(new_n206), .ZN(G42));
  INV_X1    g579(.A(new_n672), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(KEYINPUT49), .ZN(new_n767));
  XOR2_X1   g581(.A(new_n767), .B(KEYINPUT114), .Z(new_n768));
  AOI21_X1  g582(.A(new_n649), .B1(KEYINPUT49), .B2(new_n766), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n768), .A2(new_n393), .A3(new_n439), .A4(new_n769), .ZN(new_n770));
  NOR4_X1   g584(.A1(new_n770), .A2(new_n504), .A3(new_n661), .A4(new_n719), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(KEYINPUT115), .ZN(new_n772));
  INV_X1    g586(.A(new_n301), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n723), .A2(new_n773), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n774), .A2(new_n690), .A3(new_n697), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n672), .A2(new_n438), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n759), .A2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT120), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n775), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(KEYINPUT120), .B1(new_n759), .B2(new_n776), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n661), .A2(new_n393), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n774), .A2(new_n674), .A3(new_n690), .A4(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n673), .A2(new_n773), .A3(new_n696), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n721), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT119), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n693), .A2(new_n627), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n650), .A2(new_n588), .A3(new_n786), .ZN(new_n791));
  OR3_X1    g605(.A1(new_n791), .A2(new_n259), .A3(new_n718), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n785), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  OAI21_X1  g607(.A(KEYINPUT51), .B1(new_n781), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT51), .B1(new_n777), .B2(new_n775), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n795), .A2(new_n785), .A3(new_n790), .A4(new_n792), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n300), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n668), .A2(new_n694), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n637), .A2(KEYINPUT116), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n699), .A2(new_n439), .A3(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n637), .A2(KEYINPUT116), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n800), .A2(new_n662), .A3(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(KEYINPUT117), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n658), .A2(new_n680), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n804), .A2(new_n649), .A3(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n645), .A2(new_n798), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT52), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n635), .A2(new_n629), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n589), .A2(new_n656), .A3(new_n638), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n809), .A2(new_n618), .A3(new_n697), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n711), .A2(new_n789), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n811), .A2(new_n716), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT52), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n645), .A2(new_n798), .A3(new_n806), .A4(new_n814), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n808), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n259), .A2(new_n718), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n817), .B1(new_n656), .B2(new_n259), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n595), .A2(new_n608), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n819), .A2(new_n585), .A3(new_n630), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n675), .A2(new_n691), .A3(new_n678), .A4(new_n682), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(new_n713), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n816), .A2(KEYINPUT53), .A3(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n808), .A2(new_n813), .A3(new_n815), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n826), .B1(new_n827), .B2(new_n823), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(KEYINPUT54), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n774), .A2(new_n681), .A3(new_n690), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n668), .A2(new_n694), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n832), .B1(new_n643), .B2(new_n644), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n814), .B1(new_n833), .B2(new_n806), .ZN(new_n834));
  INV_X1    g648(.A(new_n815), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT118), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n821), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n838), .A2(new_n820), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n706), .A2(new_n712), .ZN(new_n840));
  OAI21_X1  g654(.A(KEYINPUT53), .B1(new_n821), .B2(new_n837), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n836), .A2(new_n813), .A3(new_n839), .A4(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n843), .A2(new_n828), .A3(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n797), .A2(new_n830), .A3(new_n831), .A4(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n791), .A2(new_n817), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n788), .A2(new_n710), .ZN(new_n848));
  XOR2_X1   g662(.A(new_n848), .B(KEYINPUT48), .Z(new_n849));
  NOR3_X1   g663(.A1(new_n846), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(G952), .A2(G953), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n772), .B1(new_n850), .B2(new_n851), .ZN(G75));
  NAND2_X1  g666(.A1(new_n428), .A2(new_n426), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(new_n423), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(KEYINPUT55), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT56), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n855), .B1(KEYINPUT121), .B2(new_n856), .ZN(new_n857));
  AOI211_X1 g671(.A(new_n510), .B(new_n243), .C1(new_n843), .C2(new_n828), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n857), .B1(new_n858), .B2(KEYINPUT56), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n189), .A2(G952), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n843), .A2(new_n828), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n862), .A2(G210), .A3(G902), .ZN(new_n863));
  INV_X1    g677(.A(new_n857), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n863), .A2(new_n856), .A3(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n859), .A2(new_n861), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT122), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT122), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n859), .A2(new_n865), .A3(new_n868), .A4(new_n861), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n867), .A2(new_n869), .ZN(G51));
  NAND2_X1  g684(.A1(new_n862), .A2(KEYINPUT54), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(new_n845), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n698), .A2(KEYINPUT57), .ZN(new_n873));
  OR2_X1    g687(.A1(new_n698), .A2(KEYINPUT57), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n382), .ZN(new_n876));
  INV_X1    g690(.A(new_n862), .ZN(new_n877));
  OR3_X1    g691(.A1(new_n877), .A2(new_n243), .A3(new_n741), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n860), .B1(new_n876), .B2(new_n878), .ZN(G54));
  NOR2_X1   g693(.A1(new_n877), .A2(new_n243), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT58), .ZN(new_n881));
  OAI21_X1  g695(.A(KEYINPUT123), .B1(new_n881), .B2(new_n187), .ZN(new_n882));
  OR3_X1    g696(.A1(new_n881), .A2(new_n187), .A3(KEYINPUT123), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n880), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(new_n250), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n880), .A2(new_n250), .A3(new_n882), .A4(new_n883), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n886), .A2(new_n861), .A3(new_n887), .ZN(G60));
  NAND2_X1  g702(.A1(G478), .A2(G902), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n889), .B(KEYINPUT59), .Z(new_n890));
  AOI21_X1  g704(.A(new_n890), .B1(new_n830), .B2(new_n845), .ZN(new_n891));
  INV_X1    g705(.A(new_n600), .ZN(new_n892));
  INV_X1    g706(.A(new_n602), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n861), .B1(new_n891), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n894), .A2(new_n890), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n872), .A2(KEYINPUT124), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT124), .B1(new_n872), .B2(new_n897), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n896), .A2(new_n898), .A3(new_n899), .ZN(G63));
  NAND2_X1  g714(.A1(G217), .A2(G902), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT60), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n862), .A2(new_n624), .A3(new_n903), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n904), .A2(new_n861), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n478), .B(new_n481), .C1(new_n877), .C2(new_n902), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT61), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n905), .A2(KEYINPUT61), .A3(new_n906), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(G66));
  OAI21_X1  g725(.A(G953), .B1(new_n304), .B2(new_n398), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n912), .B1(new_n822), .B2(G953), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n853), .B1(G898), .B2(new_n189), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n913), .B(new_n914), .ZN(G69));
  INV_X1    g729(.A(new_n764), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n753), .A2(new_n716), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n748), .A2(new_n710), .A3(new_n805), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n713), .A2(new_n833), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(KEYINPUT126), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n696), .B1(new_n733), .B2(new_n735), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n764), .B1(new_n921), .B2(new_n752), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT126), .ZN(new_n923));
  INV_X1    g737(.A(new_n919), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n922), .A2(new_n923), .A3(new_n716), .A4(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n920), .A2(new_n189), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n533), .A2(new_n535), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(new_n246), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n926), .B(new_n928), .C1(new_n636), .C2(new_n189), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n928), .B(KEYINPUT125), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n833), .A2(new_n664), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT62), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n931), .B(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n653), .A2(new_n696), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n584), .A2(new_n818), .A3(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n933), .A2(new_n922), .A3(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n930), .B1(new_n937), .B2(G953), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n929), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n940), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n929), .A2(new_n942), .A3(new_n938), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n941), .A2(new_n943), .ZN(G72));
  NAND3_X1  g758(.A1(new_n920), .A2(new_n822), .A3(new_n925), .ZN(new_n945));
  NAND2_X1  g759(.A1(G472), .A2(G902), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT63), .Z(new_n947));
  NAND2_X1  g761(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n948), .A2(new_n561), .A3(new_n543), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n829), .A2(new_n947), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n541), .A2(new_n579), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n860), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n933), .A2(new_n922), .A3(new_n822), .A4(new_n935), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n561), .B1(new_n953), .B2(new_n947), .ZN(new_n954));
  AOI21_X1  g768(.A(KEYINPUT127), .B1(new_n954), .B2(new_n578), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n954), .A2(KEYINPUT127), .A3(new_n578), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n949), .B(new_n952), .C1(new_n955), .C2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(G57));
endmodule


