

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579;

  XOR2_X1 U321 ( .A(G92GAT), .B(G85GAT), .Z(n289) );
  XOR2_X1 U322 ( .A(n434), .B(n433), .Z(n548) );
  NOR2_X1 U323 ( .A1(n520), .A2(n448), .ZN(n555) );
  XOR2_X1 U324 ( .A(n459), .B(KEYINPUT28), .Z(n515) );
  XNOR2_X1 U325 ( .A(n449), .B(G176GAT), .ZN(n450) );
  XNOR2_X1 U326 ( .A(n451), .B(n450), .ZN(G1349GAT) );
  XOR2_X1 U327 ( .A(KEYINPUT86), .B(G176GAT), .Z(n291) );
  XNOR2_X1 U328 ( .A(G120GAT), .B(KEYINPUT20), .ZN(n290) );
  XNOR2_X1 U329 ( .A(n291), .B(n290), .ZN(n309) );
  XOR2_X1 U330 ( .A(G190GAT), .B(G99GAT), .Z(n293) );
  XNOR2_X1 U331 ( .A(G43GAT), .B(G134GAT), .ZN(n292) );
  XNOR2_X1 U332 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U333 ( .A(G127GAT), .B(G71GAT), .Z(n295) );
  XNOR2_X1 U334 ( .A(G169GAT), .B(G15GAT), .ZN(n294) );
  XNOR2_X1 U335 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U336 ( .A(n297), .B(n296), .Z(n307) );
  XNOR2_X1 U337 ( .A(KEYINPUT19), .B(KEYINPUT84), .ZN(n298) );
  XNOR2_X1 U338 ( .A(n298), .B(G183GAT), .ZN(n299) );
  XOR2_X1 U339 ( .A(n299), .B(KEYINPUT85), .Z(n301) );
  XNOR2_X1 U340 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n300) );
  XNOR2_X1 U341 ( .A(n301), .B(n300), .ZN(n360) );
  XNOR2_X1 U342 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n302) );
  XNOR2_X1 U343 ( .A(n302), .B(KEYINPUT82), .ZN(n319) );
  XOR2_X1 U344 ( .A(n319), .B(KEYINPUT83), .Z(n304) );
  NAND2_X1 U345 ( .A1(G227GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U346 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U347 ( .A(n360), .B(n305), .ZN(n306) );
  XNOR2_X1 U348 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U349 ( .A(n309), .B(n308), .ZN(n520) );
  XOR2_X1 U350 ( .A(G1GAT), .B(G127GAT), .Z(n399) );
  XOR2_X1 U351 ( .A(G85GAT), .B(n399), .Z(n311) );
  XOR2_X1 U352 ( .A(G29GAT), .B(G134GAT), .Z(n429) );
  XNOR2_X1 U353 ( .A(G162GAT), .B(n429), .ZN(n310) );
  XNOR2_X1 U354 ( .A(n311), .B(n310), .ZN(n323) );
  XOR2_X1 U355 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n313) );
  XNOR2_X1 U356 ( .A(KEYINPUT96), .B(KEYINPUT6), .ZN(n312) );
  XNOR2_X1 U357 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U358 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n315) );
  XNOR2_X1 U359 ( .A(KEYINPUT95), .B(KEYINPUT1), .ZN(n314) );
  XNOR2_X1 U360 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U361 ( .A(n317), .B(n316), .Z(n321) );
  XNOR2_X1 U362 ( .A(G120GAT), .B(G148GAT), .ZN(n318) );
  XNOR2_X1 U363 ( .A(n318), .B(G57GAT), .ZN(n385) );
  XNOR2_X1 U364 ( .A(n319), .B(n385), .ZN(n320) );
  XNOR2_X1 U365 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U366 ( .A(n323), .B(n322), .Z(n325) );
  NAND2_X1 U367 ( .A1(G225GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U368 ( .A(n325), .B(n324), .ZN(n330) );
  XOR2_X1 U369 ( .A(KEYINPUT2), .B(KEYINPUT91), .Z(n327) );
  XNOR2_X1 U370 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n326) );
  XNOR2_X1 U371 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U372 ( .A(G141GAT), .B(n328), .Z(n340) );
  INV_X1 U373 ( .A(n340), .ZN(n329) );
  XNOR2_X1 U374 ( .A(n330), .B(n329), .ZN(n463) );
  XNOR2_X1 U375 ( .A(KEYINPUT97), .B(n463), .ZN(n507) );
  INV_X1 U376 ( .A(n507), .ZN(n559) );
  XOR2_X1 U377 ( .A(G50GAT), .B(G162GAT), .Z(n430) );
  XOR2_X1 U378 ( .A(KEYINPUT24), .B(KEYINPUT92), .Z(n332) );
  XNOR2_X1 U379 ( .A(G218GAT), .B(G106GAT), .ZN(n331) );
  XNOR2_X1 U380 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U381 ( .A(n430), .B(n333), .Z(n335) );
  NAND2_X1 U382 ( .A1(G228GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U383 ( .A(n335), .B(n334), .ZN(n337) );
  XNOR2_X1 U384 ( .A(G78GAT), .B(KEYINPUT72), .ZN(n336) );
  XNOR2_X1 U385 ( .A(n336), .B(G204GAT), .ZN(n380) );
  XOR2_X1 U386 ( .A(n337), .B(n380), .Z(n339) );
  XNOR2_X1 U387 ( .A(KEYINPUT87), .B(KEYINPUT88), .ZN(n338) );
  XNOR2_X1 U388 ( .A(n339), .B(n338), .ZN(n344) );
  XOR2_X1 U389 ( .A(G148GAT), .B(KEYINPUT23), .Z(n342) );
  XNOR2_X1 U390 ( .A(n340), .B(KEYINPUT22), .ZN(n341) );
  XNOR2_X1 U391 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U392 ( .A(n344), .B(n343), .Z(n349) );
  XOR2_X1 U393 ( .A(KEYINPUT21), .B(KEYINPUT90), .Z(n346) );
  XNOR2_X1 U394 ( .A(KEYINPUT89), .B(G211GAT), .ZN(n345) );
  XNOR2_X1 U395 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U396 ( .A(G197GAT), .B(n347), .Z(n356) );
  XNOR2_X1 U397 ( .A(G22GAT), .B(n356), .ZN(n348) );
  XNOR2_X1 U398 ( .A(n349), .B(n348), .ZN(n459) );
  AND2_X1 U399 ( .A1(n559), .A2(n459), .ZN(n445) );
  XOR2_X1 U400 ( .A(G169GAT), .B(G8GAT), .Z(n367) );
  XNOR2_X1 U401 ( .A(G36GAT), .B(G190GAT), .ZN(n350) );
  XNOR2_X1 U402 ( .A(n350), .B(G218GAT), .ZN(n427) );
  XNOR2_X1 U403 ( .A(n367), .B(n427), .ZN(n351) );
  XOR2_X1 U404 ( .A(G176GAT), .B(G64GAT), .Z(n389) );
  XNOR2_X1 U405 ( .A(n351), .B(n389), .ZN(n355) );
  XOR2_X1 U406 ( .A(G92GAT), .B(KEYINPUT98), .Z(n353) );
  NAND2_X1 U407 ( .A1(G226GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U408 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U409 ( .A(n355), .B(n354), .Z(n358) );
  XNOR2_X1 U410 ( .A(n356), .B(G204GAT), .ZN(n357) );
  XNOR2_X1 U411 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U412 ( .A(n360), .B(n359), .ZN(n457) );
  XOR2_X1 U413 ( .A(KEYINPUT113), .B(KEYINPUT46), .Z(n395) );
  XOR2_X1 U414 ( .A(KEYINPUT69), .B(G1GAT), .Z(n362) );
  XNOR2_X1 U415 ( .A(G141GAT), .B(G197GAT), .ZN(n361) );
  XNOR2_X1 U416 ( .A(n362), .B(n361), .ZN(n366) );
  XOR2_X1 U417 ( .A(KEYINPUT68), .B(KEYINPUT70), .Z(n364) );
  XNOR2_X1 U418 ( .A(KEYINPUT30), .B(KEYINPUT67), .ZN(n363) );
  XNOR2_X1 U419 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U420 ( .A(n366), .B(n365), .ZN(n378) );
  XOR2_X1 U421 ( .A(G113GAT), .B(G36GAT), .Z(n369) );
  XOR2_X1 U422 ( .A(G15GAT), .B(G22GAT), .Z(n402) );
  XNOR2_X1 U423 ( .A(n367), .B(n402), .ZN(n368) );
  XNOR2_X1 U424 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U425 ( .A(n370), .B(G50GAT), .Z(n376) );
  XNOR2_X1 U426 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n371) );
  XNOR2_X1 U427 ( .A(n371), .B(KEYINPUT7), .ZN(n424) );
  XOR2_X1 U428 ( .A(n424), .B(KEYINPUT29), .Z(n373) );
  NAND2_X1 U429 ( .A1(G229GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U430 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U431 ( .A(n374), .B(G29GAT), .ZN(n375) );
  XNOR2_X1 U432 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U433 ( .A(n378), .B(n377), .ZN(n562) );
  XNOR2_X1 U434 ( .A(G99GAT), .B(G106GAT), .ZN(n379) );
  XNOR2_X1 U435 ( .A(n289), .B(n379), .ZN(n423) );
  XNOR2_X1 U436 ( .A(n380), .B(n423), .ZN(n393) );
  XOR2_X1 U437 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n382) );
  NAND2_X1 U438 ( .A1(G230GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U439 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U440 ( .A(n383), .B(KEYINPUT33), .Z(n387) );
  XNOR2_X1 U441 ( .A(G71GAT), .B(KEYINPUT71), .ZN(n384) );
  XNOR2_X1 U442 ( .A(n384), .B(KEYINPUT13), .ZN(n403) );
  XNOR2_X1 U443 ( .A(n385), .B(n403), .ZN(n386) );
  XNOR2_X1 U444 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U445 ( .A(n388), .B(KEYINPUT74), .ZN(n391) );
  XOR2_X1 U446 ( .A(n389), .B(KEYINPUT73), .Z(n390) );
  XNOR2_X1 U447 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U448 ( .A(n393), .B(n392), .ZN(n568) );
  XNOR2_X1 U449 ( .A(n568), .B(KEYINPUT41), .ZN(n540) );
  NAND2_X1 U450 ( .A1(n562), .A2(n540), .ZN(n394) );
  XNOR2_X1 U451 ( .A(n395), .B(n394), .ZN(n416) );
  XOR2_X1 U452 ( .A(G155GAT), .B(G78GAT), .Z(n397) );
  XNOR2_X1 U453 ( .A(G183GAT), .B(G211GAT), .ZN(n396) );
  XNOR2_X1 U454 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U455 ( .A(n398), .B(G64GAT), .Z(n401) );
  XNOR2_X1 U456 ( .A(G8GAT), .B(n399), .ZN(n400) );
  XNOR2_X1 U457 ( .A(n401), .B(n400), .ZN(n407) );
  XOR2_X1 U458 ( .A(n403), .B(n402), .Z(n405) );
  NAND2_X1 U459 ( .A1(G231GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U460 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U461 ( .A(n407), .B(n406), .Z(n415) );
  XOR2_X1 U462 ( .A(KEYINPUT81), .B(KEYINPUT79), .Z(n409) );
  XNOR2_X1 U463 ( .A(G57GAT), .B(KEYINPUT80), .ZN(n408) );
  XNOR2_X1 U464 ( .A(n409), .B(n408), .ZN(n413) );
  XOR2_X1 U465 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n411) );
  XNOR2_X1 U466 ( .A(KEYINPUT78), .B(KEYINPUT15), .ZN(n410) );
  XNOR2_X1 U467 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U468 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U469 ( .A(n415), .B(n414), .ZN(n573) );
  INV_X1 U470 ( .A(n573), .ZN(n480) );
  AND2_X1 U471 ( .A1(n416), .A2(n480), .ZN(n417) );
  XNOR2_X1 U472 ( .A(KEYINPUT114), .B(n417), .ZN(n435) );
  XOR2_X1 U473 ( .A(KEYINPUT64), .B(KEYINPUT9), .Z(n419) );
  XNOR2_X1 U474 ( .A(KEYINPUT76), .B(KEYINPUT11), .ZN(n418) );
  XNOR2_X1 U475 ( .A(n419), .B(n418), .ZN(n434) );
  XNOR2_X1 U476 ( .A(KEYINPUT75), .B(KEYINPUT66), .ZN(n421) );
  AND2_X1 U477 ( .A1(G232GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U478 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n422), .B(KEYINPUT10), .ZN(n426) );
  XNOR2_X1 U480 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U481 ( .A(n426), .B(n425), .ZN(n428) );
  XNOR2_X1 U482 ( .A(n428), .B(n427), .ZN(n432) );
  XNOR2_X1 U483 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U484 ( .A(n432), .B(n431), .ZN(n433) );
  NAND2_X1 U485 ( .A1(n435), .A2(n548), .ZN(n436) );
  XNOR2_X1 U486 ( .A(n436), .B(KEYINPUT47), .ZN(n442) );
  XNOR2_X1 U487 ( .A(KEYINPUT77), .B(n548), .ZN(n554) );
  XNOR2_X1 U488 ( .A(KEYINPUT36), .B(n554), .ZN(n575) );
  NAND2_X1 U489 ( .A1(n575), .A2(n573), .ZN(n438) );
  XNOR2_X1 U490 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n437) );
  XNOR2_X1 U491 ( .A(n438), .B(n437), .ZN(n439) );
  NAND2_X1 U492 ( .A1(n439), .A2(n568), .ZN(n440) );
  NOR2_X1 U493 ( .A1(n440), .A2(n562), .ZN(n441) );
  NOR2_X1 U494 ( .A1(n442), .A2(n441), .ZN(n443) );
  XNOR2_X1 U495 ( .A(n443), .B(KEYINPUT48), .ZN(n519) );
  NOR2_X1 U496 ( .A1(n457), .A2(n519), .ZN(n444) );
  XNOR2_X1 U497 ( .A(n444), .B(KEYINPUT54), .ZN(n558) );
  NAND2_X1 U498 ( .A1(n445), .A2(n558), .ZN(n446) );
  XNOR2_X1 U499 ( .A(n446), .B(KEYINPUT121), .ZN(n447) );
  XNOR2_X1 U500 ( .A(n447), .B(KEYINPUT55), .ZN(n448) );
  XOR2_X1 U501 ( .A(KEYINPUT107), .B(n540), .Z(n525) );
  NAND2_X1 U502 ( .A1(n555), .A2(n525), .ZN(n451) );
  XOR2_X1 U503 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n449) );
  XOR2_X1 U504 ( .A(KEYINPUT101), .B(KEYINPUT34), .Z(n469) );
  NAND2_X1 U505 ( .A1(n562), .A2(n568), .ZN(n484) );
  NOR2_X1 U506 ( .A1(n554), .A2(n480), .ZN(n452) );
  XNOR2_X1 U507 ( .A(n452), .B(KEYINPUT16), .ZN(n467) );
  XOR2_X1 U508 ( .A(KEYINPUT27), .B(n457), .Z(n456) );
  NAND2_X1 U509 ( .A1(n456), .A2(n507), .ZN(n453) );
  XOR2_X1 U510 ( .A(KEYINPUT99), .B(n453), .Z(n535) );
  NOR2_X1 U511 ( .A1(n515), .A2(n535), .ZN(n522) );
  XNOR2_X1 U512 ( .A(KEYINPUT100), .B(n522), .ZN(n454) );
  NAND2_X1 U513 ( .A1(n454), .A2(n520), .ZN(n466) );
  INV_X1 U514 ( .A(n520), .ZN(n512) );
  NOR2_X1 U515 ( .A1(n459), .A2(n512), .ZN(n455) );
  XNOR2_X1 U516 ( .A(n455), .B(KEYINPUT26), .ZN(n560) );
  NAND2_X1 U517 ( .A1(n456), .A2(n560), .ZN(n462) );
  INV_X1 U518 ( .A(n457), .ZN(n509) );
  NAND2_X1 U519 ( .A1(n512), .A2(n509), .ZN(n458) );
  NAND2_X1 U520 ( .A1(n459), .A2(n458), .ZN(n460) );
  XOR2_X1 U521 ( .A(KEYINPUT25), .B(n460), .Z(n461) );
  NAND2_X1 U522 ( .A1(n462), .A2(n461), .ZN(n464) );
  NAND2_X1 U523 ( .A1(n464), .A2(n463), .ZN(n465) );
  NAND2_X1 U524 ( .A1(n466), .A2(n465), .ZN(n479) );
  NAND2_X1 U525 ( .A1(n467), .A2(n479), .ZN(n494) );
  NOR2_X1 U526 ( .A1(n484), .A2(n494), .ZN(n477) );
  NAND2_X1 U527 ( .A1(n477), .A2(n507), .ZN(n468) );
  XNOR2_X1 U528 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U529 ( .A(G1GAT), .B(n470), .ZN(G1324GAT) );
  XOR2_X1 U530 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n472) );
  NAND2_X1 U531 ( .A1(n477), .A2(n509), .ZN(n471) );
  XNOR2_X1 U532 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U533 ( .A(G8GAT), .B(n473), .ZN(G1325GAT) );
  XOR2_X1 U534 ( .A(KEYINPUT104), .B(KEYINPUT35), .Z(n475) );
  NAND2_X1 U535 ( .A1(n477), .A2(n512), .ZN(n474) );
  XNOR2_X1 U536 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U537 ( .A(G15GAT), .B(n476), .ZN(G1326GAT) );
  NAND2_X1 U538 ( .A1(n477), .A2(n515), .ZN(n478) );
  XNOR2_X1 U539 ( .A(n478), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U540 ( .A(G29GAT), .B(KEYINPUT39), .Z(n488) );
  NAND2_X1 U541 ( .A1(n480), .A2(n479), .ZN(n481) );
  XNOR2_X1 U542 ( .A(KEYINPUT105), .B(n481), .ZN(n482) );
  NAND2_X1 U543 ( .A1(n482), .A2(n575), .ZN(n483) );
  XOR2_X1 U544 ( .A(KEYINPUT37), .B(n483), .Z(n504) );
  NOR2_X1 U545 ( .A1(n504), .A2(n484), .ZN(n486) );
  XNOR2_X1 U546 ( .A(KEYINPUT106), .B(KEYINPUT38), .ZN(n485) );
  XNOR2_X1 U547 ( .A(n486), .B(n485), .ZN(n492) );
  NAND2_X1 U548 ( .A1(n492), .A2(n507), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n488), .B(n487), .ZN(G1328GAT) );
  NAND2_X1 U550 ( .A1(n492), .A2(n509), .ZN(n489) );
  XNOR2_X1 U551 ( .A(n489), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U552 ( .A1(n492), .A2(n512), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n490), .B(KEYINPUT40), .ZN(n491) );
  XNOR2_X1 U554 ( .A(G43GAT), .B(n491), .ZN(G1330GAT) );
  NAND2_X1 U555 ( .A1(n492), .A2(n515), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n493), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U557 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n496) );
  INV_X1 U558 ( .A(n562), .ZN(n537) );
  NAND2_X1 U559 ( .A1(n537), .A2(n525), .ZN(n505) );
  NOR2_X1 U560 ( .A1(n505), .A2(n494), .ZN(n501) );
  NAND2_X1 U561 ( .A1(n501), .A2(n507), .ZN(n495) );
  XNOR2_X1 U562 ( .A(n496), .B(n495), .ZN(G1332GAT) );
  NAND2_X1 U563 ( .A1(n501), .A2(n509), .ZN(n497) );
  XNOR2_X1 U564 ( .A(n497), .B(KEYINPUT108), .ZN(n498) );
  XNOR2_X1 U565 ( .A(G64GAT), .B(n498), .ZN(G1333GAT) );
  XOR2_X1 U566 ( .A(G71GAT), .B(KEYINPUT109), .Z(n500) );
  NAND2_X1 U567 ( .A1(n501), .A2(n512), .ZN(n499) );
  XNOR2_X1 U568 ( .A(n500), .B(n499), .ZN(G1334GAT) );
  XOR2_X1 U569 ( .A(G78GAT), .B(KEYINPUT43), .Z(n503) );
  NAND2_X1 U570 ( .A1(n501), .A2(n515), .ZN(n502) );
  XNOR2_X1 U571 ( .A(n503), .B(n502), .ZN(G1335GAT) );
  NOR2_X1 U572 ( .A1(n505), .A2(n504), .ZN(n506) );
  XNOR2_X1 U573 ( .A(n506), .B(KEYINPUT110), .ZN(n516) );
  NAND2_X1 U574 ( .A1(n516), .A2(n507), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n508), .B(G85GAT), .ZN(G1336GAT) );
  XOR2_X1 U576 ( .A(G92GAT), .B(KEYINPUT111), .Z(n511) );
  NAND2_X1 U577 ( .A1(n509), .A2(n516), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n511), .B(n510), .ZN(G1337GAT) );
  NAND2_X1 U579 ( .A1(n516), .A2(n512), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n513), .B(KEYINPUT112), .ZN(n514) );
  XNOR2_X1 U581 ( .A(G99GAT), .B(n514), .ZN(G1338GAT) );
  NAND2_X1 U582 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n517), .B(KEYINPUT44), .ZN(n518) );
  XNOR2_X1 U584 ( .A(G106GAT), .B(n518), .ZN(G1339GAT) );
  NOR2_X1 U585 ( .A1(n520), .A2(n519), .ZN(n521) );
  NAND2_X1 U586 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U587 ( .A(KEYINPUT115), .B(n523), .ZN(n532) );
  NAND2_X1 U588 ( .A1(n532), .A2(n562), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n524), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U590 ( .A(G120GAT), .B(KEYINPUT49), .Z(n527) );
  NAND2_X1 U591 ( .A1(n532), .A2(n525), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n527), .B(n526), .ZN(G1341GAT) );
  XNOR2_X1 U593 ( .A(G127GAT), .B(KEYINPUT117), .ZN(n531) );
  XOR2_X1 U594 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n529) );
  NAND2_X1 U595 ( .A1(n532), .A2(n573), .ZN(n528) );
  XNOR2_X1 U596 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U597 ( .A(n531), .B(n530), .ZN(G1342GAT) );
  XOR2_X1 U598 ( .A(G134GAT), .B(KEYINPUT51), .Z(n534) );
  NAND2_X1 U599 ( .A1(n532), .A2(n554), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(G1343GAT) );
  NOR2_X1 U601 ( .A1(n519), .A2(n535), .ZN(n536) );
  NAND2_X1 U602 ( .A1(n536), .A2(n560), .ZN(n547) );
  NOR2_X1 U603 ( .A1(n537), .A2(n547), .ZN(n538) );
  XOR2_X1 U604 ( .A(KEYINPUT118), .B(n538), .Z(n539) );
  XNOR2_X1 U605 ( .A(G141GAT), .B(n539), .ZN(G1344GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n542) );
  INV_X1 U607 ( .A(n547), .ZN(n544) );
  NAND2_X1 U608 ( .A1(n544), .A2(n540), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(n543), .ZN(G1345GAT) );
  XOR2_X1 U611 ( .A(G155GAT), .B(KEYINPUT119), .Z(n546) );
  NAND2_X1 U612 ( .A1(n544), .A2(n573), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(G1346GAT) );
  NOR2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U615 ( .A(KEYINPUT120), .B(n549), .Z(n550) );
  XNOR2_X1 U616 ( .A(G162GAT), .B(n550), .ZN(G1347GAT) );
  NAND2_X1 U617 ( .A1(n555), .A2(n562), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n551), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U619 ( .A1(n555), .A2(n573), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n552), .B(KEYINPUT122), .ZN(n553) );
  XNOR2_X1 U621 ( .A(G183GAT), .B(n553), .ZN(G1350GAT) );
  NAND2_X1 U622 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(KEYINPUT58), .ZN(n557) );
  XNOR2_X1 U624 ( .A(G190GAT), .B(n557), .ZN(G1351GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT124), .B(KEYINPUT60), .Z(n564) );
  AND2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n561) );
  AND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n576) );
  NAND2_X1 U628 ( .A1(n576), .A2(n562), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n564), .B(n563), .ZN(n565) );
  XOR2_X1 U630 ( .A(n565), .B(KEYINPUT123), .Z(n567) );
  XNOR2_X1 U631 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(G1352GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n571) );
  INV_X1 U634 ( .A(n568), .ZN(n569) );
  NAND2_X1 U635 ( .A1(n576), .A2(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XOR2_X1 U637 ( .A(G204GAT), .B(n572), .Z(G1353GAT) );
  NAND2_X1 U638 ( .A1(n576), .A2(n573), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n578) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(n579) );
  XOR2_X1 U643 ( .A(G218GAT), .B(n579), .Z(G1355GAT) );
endmodule

