

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737;

  NOR2_X1 U363 ( .A1(G953), .A2(KEYINPUT83), .ZN(n443) );
  NOR2_X1 U364 ( .A1(G237), .A2(G953), .ZN(n517) );
  XNOR2_X1 U365 ( .A(n441), .B(G110), .ZN(n440) );
  NAND2_X1 U366 ( .A1(n366), .A2(n363), .ZN(n652) );
  NOR2_X2 U367 ( .A1(n428), .A2(KEYINPUT44), .ZN(n606) );
  NOR2_X2 U368 ( .A1(n557), .A2(n556), .ZN(n455) );
  NAND2_X2 U369 ( .A1(n400), .A2(n353), .ZN(n590) );
  NOR2_X2 U370 ( .A1(n546), .A2(n545), .ZN(n548) );
  NAND2_X2 U371 ( .A1(n407), .A2(n406), .ZN(n612) );
  XNOR2_X2 U372 ( .A(n485), .B(n486), .ZN(n720) );
  XNOR2_X2 U373 ( .A(n584), .B(KEYINPUT33), .ZN(n680) );
  AND2_X1 U374 ( .A1(n654), .A2(n394), .ZN(n533) );
  NOR2_X1 U375 ( .A1(n615), .A2(G902), .ZN(n397) );
  NOR2_X1 U376 ( .A1(n649), .A2(n448), .ZN(n447) );
  AND2_X1 U377 ( .A1(n385), .A2(n384), .ZN(n383) );
  NOR2_X1 U378 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U379 ( .A(n533), .B(KEYINPUT98), .ZN(n595) );
  BUF_X1 U380 ( .A(n599), .Z(n391) );
  AND2_X1 U381 ( .A1(n552), .A2(n542), .ZN(n559) );
  AND2_X1 U382 ( .A1(n368), .A2(n367), .ZN(n366) );
  OR2_X1 U383 ( .A1(n449), .A2(KEYINPUT71), .ZN(n346) );
  XNOR2_X1 U384 ( .A(n397), .B(n396), .ZN(n394) );
  XNOR2_X1 U385 ( .A(n489), .B(n452), .ZN(n451) );
  XNOR2_X1 U386 ( .A(n481), .B(n446), .ZN(n502) );
  XNOR2_X1 U387 ( .A(n412), .B(n469), .ZN(n523) );
  XNOR2_X1 U388 ( .A(n472), .B(G134), .ZN(n501) );
  XNOR2_X1 U389 ( .A(n468), .B(n462), .ZN(n412) );
  XOR2_X1 U390 ( .A(G146), .B(G125), .Z(n484) );
  XNOR2_X1 U391 ( .A(G116), .B(G119), .ZN(n468) );
  XNOR2_X1 U392 ( .A(G902), .B(KEYINPUT15), .ZN(n610) );
  XNOR2_X1 U393 ( .A(KEYINPUT73), .B(KEYINPUT3), .ZN(n462) );
  XOR2_X1 U394 ( .A(G113), .B(KEYINPUT72), .Z(n469) );
  BUF_X1 U395 ( .A(n539), .Z(n343) );
  BUF_X1 U396 ( .A(n731), .Z(n344) );
  BUF_X1 U397 ( .A(n453), .Z(n345) );
  OR2_X2 U398 ( .A1(n587), .A2(n588), .ZN(n431) );
  XNOR2_X2 U399 ( .A(KEYINPUT32), .B(n590), .ZN(n734) );
  NAND2_X1 U400 ( .A1(n640), .A2(n594), .ZN(n544) );
  OR2_X1 U401 ( .A1(n704), .A2(n364), .ZN(n363) );
  NAND2_X1 U402 ( .A1(n451), .A2(n365), .ZN(n364) );
  INV_X1 U403 ( .A(G902), .ZN(n365) );
  NAND2_X1 U404 ( .A1(n370), .A2(G902), .ZN(n367) );
  INV_X1 U405 ( .A(n451), .ZN(n370) );
  XNOR2_X1 U406 ( .A(n480), .B(KEYINPUT94), .ZN(n665) );
  XNOR2_X1 U407 ( .A(n720), .B(n427), .ZN(n426) );
  INV_X1 U408 ( .A(n552), .ZN(n425) );
  INV_X1 U409 ( .A(KEYINPUT81), .ZN(n409) );
  XOR2_X1 U410 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n515) );
  INV_X1 U411 ( .A(KEYINPUT90), .ZN(n416) );
  NOR2_X1 U412 ( .A1(n437), .A2(n436), .ZN(n435) );
  INV_X1 U413 ( .A(n609), .ZN(n436) );
  INV_X1 U414 ( .A(n447), .ZN(n437) );
  XNOR2_X1 U415 ( .A(n397), .B(n390), .ZN(n389) );
  NAND2_X1 U416 ( .A1(n360), .A2(n652), .ZN(n359) );
  NOR2_X1 U417 ( .A1(n361), .A2(n369), .ZN(n360) );
  XNOR2_X1 U418 ( .A(n376), .B(n375), .ZN(n374) );
  XNOR2_X1 U419 ( .A(G119), .B(G137), .ZN(n375) );
  XNOR2_X1 U420 ( .A(n377), .B(G110), .ZN(n376) );
  INV_X1 U421 ( .A(G128), .ZN(n377) );
  XNOR2_X1 U422 ( .A(n373), .B(n372), .ZN(n371) );
  XNOR2_X1 U423 ( .A(KEYINPUT23), .B(KEYINPUT97), .ZN(n373) );
  XNOR2_X1 U424 ( .A(KEYINPUT24), .B(KEYINPUT82), .ZN(n372) );
  NAND2_X1 U425 ( .A1(n445), .A2(n444), .ZN(n446) );
  NAND2_X1 U426 ( .A1(n443), .A2(G234), .ZN(n444) );
  XOR2_X1 U427 ( .A(KEYINPUT70), .B(KEYINPUT10), .Z(n486) );
  XOR2_X1 U428 ( .A(KEYINPUT9), .B(G122), .Z(n499) );
  XNOR2_X1 U429 ( .A(G107), .B(G116), .ZN(n498) );
  XNOR2_X1 U430 ( .A(n471), .B(n713), .ZN(n690) );
  NAND2_X1 U431 ( .A1(n391), .A2(n382), .ZN(n381) );
  NAND2_X1 U432 ( .A1(n380), .A2(n595), .ZN(n557) );
  AND2_X1 U433 ( .A1(n532), .A2(n531), .ZN(n380) );
  XNOR2_X1 U434 ( .A(n520), .B(n521), .ZN(n542) );
  XNOR2_X1 U435 ( .A(KEYINPUT66), .B(KEYINPUT22), .ZN(n580) );
  INV_X2 U436 ( .A(G953), .ZN(n726) );
  AND2_X1 U437 ( .A1(n531), .A2(n450), .ZN(n449) );
  INV_X1 U438 ( .A(n651), .ZN(n450) );
  INV_X1 U439 ( .A(KEYINPUT25), .ZN(n452) );
  XNOR2_X1 U440 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n421) );
  OR2_X1 U441 ( .A1(G902), .A2(G237), .ZN(n479) );
  INV_X1 U442 ( .A(n449), .ZN(n361) );
  NAND2_X1 U443 ( .A1(n348), .A2(n366), .ZN(n362) );
  INV_X1 U444 ( .A(G469), .ZN(n396) );
  INV_X1 U445 ( .A(G101), .ZN(n461) );
  INV_X1 U446 ( .A(n648), .ZN(n448) );
  XNOR2_X1 U447 ( .A(n501), .B(n474), .ZN(n719) );
  NAND2_X1 U448 ( .A1(n442), .A2(KEYINPUT83), .ZN(n445) );
  NAND2_X1 U449 ( .A1(n726), .A2(G234), .ZN(n442) );
  XNOR2_X1 U450 ( .A(n516), .B(n518), .ZN(n427) );
  XNOR2_X1 U451 ( .A(KEYINPUT12), .B(KEYINPUT11), .ZN(n514) );
  XOR2_X1 U452 ( .A(G113), .B(G131), .Z(n510) );
  XOR2_X1 U453 ( .A(KEYINPUT96), .B(G140), .Z(n477) );
  XNOR2_X1 U454 ( .A(n719), .B(G146), .ZN(n522) );
  XNOR2_X1 U455 ( .A(n484), .B(n418), .ZN(n466) );
  XNOR2_X1 U456 ( .A(n420), .B(n419), .ZN(n418) );
  XNOR2_X1 U457 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n420) );
  NAND2_X1 U458 ( .A1(n726), .A2(G224), .ZN(n419) );
  XNOR2_X1 U459 ( .A(n550), .B(KEYINPUT112), .ZN(n669) );
  INV_X1 U460 ( .A(KEYINPUT34), .ZN(n386) );
  INV_X1 U461 ( .A(n542), .ZN(n551) );
  XNOR2_X1 U462 ( .A(n522), .B(n458), .ZN(n623) );
  XNOR2_X1 U463 ( .A(n523), .B(n459), .ZN(n458) );
  XNOR2_X1 U464 ( .A(n347), .B(n460), .ZN(n459) );
  XNOR2_X1 U465 ( .A(n461), .B(KEYINPUT5), .ZN(n460) );
  NAND2_X1 U466 ( .A1(n433), .A2(n434), .ZN(n432) );
  NAND2_X1 U467 ( .A1(n609), .A2(KEYINPUT2), .ZN(n434) );
  NOR2_X1 U468 ( .A1(n583), .A2(n598), .ZN(n584) );
  XNOR2_X1 U469 ( .A(n378), .B(KEYINPUT41), .ZN(n650) );
  NOR2_X1 U470 ( .A1(n669), .A2(n667), .ZN(n378) );
  AND2_X1 U471 ( .A1(n642), .A2(n404), .ZN(n526) );
  XNOR2_X1 U472 ( .A(n439), .B(G101), .ZN(n438) );
  INV_X1 U473 ( .A(KEYINPUT93), .ZN(n439) );
  XNOR2_X1 U474 ( .A(G122), .B(KEYINPUT16), .ZN(n470) );
  XNOR2_X1 U475 ( .A(n374), .B(n371), .ZN(n483) );
  XOR2_X1 U476 ( .A(n506), .B(n505), .Z(n619) );
  XNOR2_X1 U477 ( .A(n697), .B(n696), .ZN(n698) );
  XNOR2_X1 U478 ( .A(KEYINPUT92), .B(n616), .ZN(n706) );
  XNOR2_X1 U479 ( .A(n387), .B(n355), .ZN(n731) );
  NOR2_X2 U480 ( .A1(n553), .A2(n429), .ZN(n640) );
  NOR2_X1 U481 ( .A1(n557), .A2(n379), .ZN(n534) );
  AND2_X1 U482 ( .A1(n582), .A2(n402), .ZN(n635) );
  NOR2_X1 U483 ( .A1(n398), .A2(n591), .ZN(n402) );
  INV_X1 U484 ( .A(n591), .ZN(n430) );
  AND2_X1 U485 ( .A1(n524), .A2(G210), .ZN(n347) );
  AND2_X1 U486 ( .A1(n363), .A2(n369), .ZN(n348) );
  XOR2_X1 U487 ( .A(KEYINPUT6), .B(KEYINPUT106), .Z(n349) );
  XNOR2_X1 U488 ( .A(n657), .B(n349), .ZN(n583) );
  AND2_X1 U489 ( .A1(n346), .A2(n362), .ZN(n350) );
  AND2_X1 U490 ( .A1(n542), .A2(n425), .ZN(n351) );
  AND2_X1 U491 ( .A1(G210), .A2(n479), .ZN(n352) );
  AND2_X1 U492 ( .A1(n589), .A2(n583), .ZN(n353) );
  XOR2_X1 U493 ( .A(n577), .B(KEYINPUT91), .Z(n354) );
  XOR2_X1 U494 ( .A(n586), .B(KEYINPUT86), .Z(n355) );
  INV_X1 U495 ( .A(KEYINPUT71), .ZN(n369) );
  OR2_X1 U496 ( .A1(KEYINPUT2), .A2(n611), .ZN(n356) );
  XOR2_X1 U497 ( .A(KEYINPUT48), .B(KEYINPUT88), .Z(n357) );
  NAND2_X1 U498 ( .A1(n358), .A2(n730), .ZN(n410) );
  NAND2_X1 U499 ( .A1(n544), .A2(KEYINPUT47), .ZN(n358) );
  NAND2_X1 U500 ( .A1(n350), .A2(n359), .ZN(n535) );
  NAND2_X1 U501 ( .A1(n704), .A2(n370), .ZN(n368) );
  NOR2_X2 U502 ( .A1(n650), .A2(n553), .ZN(n555) );
  NAND2_X1 U503 ( .A1(n351), .A2(n343), .ZN(n379) );
  XNOR2_X2 U504 ( .A(n525), .B(G472), .ZN(n657) );
  NAND2_X1 U505 ( .A1(n383), .A2(n381), .ZN(n388) );
  NOR2_X1 U506 ( .A1(n680), .A2(n386), .ZN(n382) );
  NAND2_X1 U507 ( .A1(n680), .A2(n386), .ZN(n384) );
  NAND2_X1 U508 ( .A1(n585), .A2(n386), .ZN(n385) );
  NAND2_X1 U509 ( .A1(n388), .A2(n351), .ZN(n387) );
  NAND2_X1 U510 ( .A1(n654), .A2(n389), .ZN(n598) );
  XNOR2_X1 U511 ( .A(n396), .B(KEYINPUT1), .ZN(n390) );
  XNOR2_X1 U512 ( .A(G122), .B(n401), .ZN(n509) );
  BUF_X1 U513 ( .A(G104), .Z(n401) );
  NAND2_X1 U514 ( .A1(n424), .A2(n447), .ZN(n724) );
  NOR2_X1 U515 ( .A1(n535), .A2(n583), .ZN(n404) );
  BUF_X1 U516 ( .A(n685), .Z(n392) );
  BUF_X1 U517 ( .A(n709), .Z(n393) );
  XNOR2_X1 U518 ( .A(n539), .B(n549), .ZN(n664) );
  XNOR2_X1 U519 ( .A(n714), .B(KEYINPUT74), .ZN(n395) );
  XNOR2_X1 U520 ( .A(n714), .B(KEYINPUT74), .ZN(n475) );
  XNOR2_X2 U521 ( .A(n413), .B(n541), .ZN(n576) );
  NAND2_X2 U522 ( .A1(n576), .A2(n575), .ZN(n578) );
  XNOR2_X1 U523 ( .A(n422), .B(n421), .ZN(n561) );
  NAND2_X1 U524 ( .A1(n736), .A2(n737), .ZN(n422) );
  XNOR2_X1 U525 ( .A(n487), .B(n720), .ZN(n704) );
  XNOR2_X1 U526 ( .A(n623), .B(n622), .ZN(n624) );
  NOR2_X1 U527 ( .A1(n587), .A2(n597), .ZN(n582) );
  XNOR2_X1 U528 ( .A(n410), .B(n409), .ZN(n546) );
  XNOR2_X1 U529 ( .A(n394), .B(KEYINPUT1), .ZN(n398) );
  XNOR2_X1 U530 ( .A(n408), .B(n522), .ZN(n615) );
  XNOR2_X1 U531 ( .A(n475), .B(n478), .ZN(n408) );
  XNOR2_X1 U532 ( .A(n455), .B(n558), .ZN(n570) );
  BUF_X1 U533 ( .A(n576), .Z(n399) );
  INV_X1 U534 ( .A(KEYINPUT2), .ZN(n457) );
  INV_X1 U535 ( .A(n587), .ZN(n400) );
  XNOR2_X2 U536 ( .A(n581), .B(n580), .ZN(n587) );
  NAND2_X1 U537 ( .A1(n607), .A2(n414), .ZN(n403) );
  XNOR2_X2 U538 ( .A(n403), .B(n608), .ZN(n709) );
  XNOR2_X2 U539 ( .A(n569), .B(n357), .ZN(n424) );
  XNOR2_X1 U540 ( .A(n519), .B(n426), .ZN(n697) );
  XNOR2_X1 U541 ( .A(n613), .B(n405), .ZN(n617) );
  XNOR2_X1 U542 ( .A(n615), .B(n614), .ZN(n405) );
  NAND2_X1 U543 ( .A1(n685), .A2(n356), .ZN(n406) );
  NAND2_X1 U544 ( .A1(n411), .A2(KEYINPUT84), .ZN(n407) );
  NAND2_X1 U545 ( .A1(n605), .A2(n604), .ZN(n417) );
  XNOR2_X2 U546 ( .A(n440), .B(n438), .ZN(n714) );
  NAND2_X1 U547 ( .A1(n456), .A2(n432), .ZN(n411) );
  NAND2_X1 U548 ( .A1(n539), .A2(n665), .ZN(n413) );
  INV_X1 U549 ( .A(n599), .ZN(n585) );
  NAND2_X1 U550 ( .A1(n599), .A2(n579), .ZN(n581) );
  XNOR2_X2 U551 ( .A(n578), .B(n354), .ZN(n599) );
  NAND2_X1 U552 ( .A1(n709), .A2(n457), .ZN(n456) );
  XNOR2_X1 U553 ( .A(n606), .B(KEYINPUT75), .ZN(n414) );
  NOR2_X2 U554 ( .A1(n709), .A2(n724), .ZN(n685) );
  NAND2_X1 U555 ( .A1(n415), .A2(n734), .ZN(n428) );
  NOR2_X1 U556 ( .A1(n731), .A2(n635), .ZN(n415) );
  XNOR2_X1 U557 ( .A(n417), .B(n416), .ZN(n607) );
  XNOR2_X2 U558 ( .A(n555), .B(n554), .ZN(n736) );
  INV_X1 U559 ( .A(n343), .ZN(n564) );
  XNOR2_X2 U560 ( .A(n423), .B(n352), .ZN(n539) );
  NAND2_X1 U561 ( .A1(n690), .A2(n610), .ZN(n423) );
  NAND2_X1 U562 ( .A1(n424), .A2(n435), .ZN(n433) );
  NAND2_X1 U563 ( .A1(n428), .A2(KEYINPUT44), .ZN(n605) );
  INV_X1 U564 ( .A(n399), .ZN(n429) );
  NOR2_X1 U565 ( .A1(n431), .A2(n430), .ZN(n592) );
  XNOR2_X2 U566 ( .A(G107), .B(G104), .ZN(n441) );
  NAND2_X1 U567 ( .A1(n453), .A2(G478), .ZN(n618) );
  NAND2_X1 U568 ( .A1(n453), .A2(G472), .ZN(n625) );
  NAND2_X1 U569 ( .A1(n453), .A2(G210), .ZN(n692) );
  NAND2_X1 U570 ( .A1(n453), .A2(G475), .ZN(n699) );
  NAND2_X1 U571 ( .A1(n345), .A2(G469), .ZN(n613) );
  NAND2_X1 U572 ( .A1(n345), .A2(G217), .ZN(n703) );
  XNOR2_X2 U573 ( .A(n612), .B(KEYINPUT65), .ZN(n453) );
  XNOR2_X2 U574 ( .A(n454), .B(n560), .ZN(n737) );
  NAND2_X1 U575 ( .A1(n570), .A2(n559), .ZN(n454) );
  NOR2_X2 U576 ( .A1(n651), .A2(n652), .ZN(n654) );
  XOR2_X2 U577 ( .A(KEYINPUT107), .B(n559), .Z(n642) );
  XNOR2_X1 U578 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n463) );
  INV_X1 U579 ( .A(KEYINPUT76), .ZN(n547) );
  INV_X1 U580 ( .A(n629), .ZN(n603) );
  NOR2_X1 U581 ( .A1(n603), .A2(n602), .ZN(n604) );
  BUF_X1 U582 ( .A(n650), .Z(n681) );
  XNOR2_X1 U583 ( .A(n690), .B(n463), .ZN(n691) );
  INV_X1 U584 ( .A(KEYINPUT63), .ZN(n627) );
  XOR2_X1 U585 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n614) );
  XNOR2_X2 U586 ( .A(G143), .B(G128), .ZN(n472) );
  INV_X1 U587 ( .A(n472), .ZN(n464) );
  XNOR2_X1 U588 ( .A(n464), .B(KEYINPUT4), .ZN(n465) );
  XNOR2_X1 U589 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U590 ( .A(n395), .B(n467), .ZN(n471) );
  XOR2_X1 U591 ( .A(n470), .B(n523), .Z(n713) );
  XNOR2_X1 U592 ( .A(G131), .B(KEYINPUT4), .ZN(n473) );
  XNOR2_X1 U593 ( .A(n473), .B(G137), .ZN(n474) );
  NAND2_X1 U594 ( .A1(G227), .A2(n726), .ZN(n476) );
  XNOR2_X1 U595 ( .A(n477), .B(n476), .ZN(n478) );
  NAND2_X1 U596 ( .A1(n479), .A2(G214), .ZN(n480) );
  XOR2_X1 U597 ( .A(KEYINPUT8), .B(KEYINPUT69), .Z(n481) );
  NAND2_X1 U598 ( .A1(G221), .A2(n502), .ZN(n482) );
  XNOR2_X1 U599 ( .A(n483), .B(n482), .ZN(n487) );
  XNOR2_X1 U600 ( .A(G140), .B(n484), .ZN(n485) );
  NAND2_X1 U601 ( .A1(n610), .A2(G234), .ZN(n488) );
  XNOR2_X1 U602 ( .A(n488), .B(KEYINPUT20), .ZN(n496) );
  NAND2_X1 U603 ( .A1(G217), .A2(n496), .ZN(n489) );
  NAND2_X1 U604 ( .A1(G237), .A2(G234), .ZN(n490) );
  XNOR2_X1 U605 ( .A(n490), .B(KEYINPUT14), .ZN(n492) );
  NAND2_X1 U606 ( .A1(G902), .A2(n492), .ZN(n571) );
  NOR2_X1 U607 ( .A1(G900), .A2(n571), .ZN(n491) );
  NAND2_X1 U608 ( .A1(n491), .A2(G953), .ZN(n494) );
  NAND2_X1 U609 ( .A1(G952), .A2(n492), .ZN(n678) );
  NOR2_X1 U610 ( .A1(n678), .A2(G953), .ZN(n493) );
  XNOR2_X1 U611 ( .A(n493), .B(KEYINPUT95), .ZN(n573) );
  NAND2_X1 U612 ( .A1(n494), .A2(n573), .ZN(n495) );
  XNOR2_X1 U613 ( .A(n495), .B(KEYINPUT80), .ZN(n531) );
  NAND2_X1 U614 ( .A1(G221), .A2(n496), .ZN(n497) );
  XNOR2_X1 U615 ( .A(KEYINPUT21), .B(n497), .ZN(n651) );
  XNOR2_X1 U616 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U617 ( .A(n501), .B(n500), .ZN(n506) );
  XOR2_X1 U618 ( .A(KEYINPUT103), .B(KEYINPUT7), .Z(n504) );
  NAND2_X1 U619 ( .A1(G217), .A2(n502), .ZN(n503) );
  XNOR2_X1 U620 ( .A(n504), .B(n503), .ZN(n505) );
  NOR2_X1 U621 ( .A1(G902), .A2(n619), .ZN(n508) );
  XNOR2_X1 U622 ( .A(G478), .B(KEYINPUT104), .ZN(n507) );
  XNOR2_X1 U623 ( .A(n508), .B(n507), .ZN(n552) );
  XNOR2_X1 U624 ( .A(KEYINPUT13), .B(G475), .ZN(n521) );
  XNOR2_X1 U625 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U626 ( .A(n511), .B(KEYINPUT99), .Z(n513) );
  XNOR2_X1 U627 ( .A(G143), .B(KEYINPUT102), .ZN(n512) );
  XNOR2_X1 U628 ( .A(n513), .B(n512), .ZN(n519) );
  XNOR2_X1 U629 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U630 ( .A(n517), .B(KEYINPUT78), .ZN(n524) );
  NAND2_X1 U631 ( .A1(G214), .A2(n524), .ZN(n518) );
  NOR2_X1 U632 ( .A1(G902), .A2(n697), .ZN(n520) );
  NOR2_X1 U633 ( .A1(n623), .A2(G902), .ZN(n525) );
  INV_X1 U634 ( .A(n583), .ZN(n588) );
  NAND2_X1 U635 ( .A1(n665), .A2(n526), .ZN(n563) );
  NOR2_X1 U636 ( .A1(n398), .A2(n563), .ZN(n527) );
  XNOR2_X1 U637 ( .A(n527), .B(KEYINPUT43), .ZN(n528) );
  NOR2_X1 U638 ( .A1(n343), .A2(n528), .ZN(n649) );
  XOR2_X1 U639 ( .A(KEYINPUT30), .B(KEYINPUT108), .Z(n530) );
  INV_X1 U640 ( .A(n657), .ZN(n597) );
  NAND2_X1 U641 ( .A1(n597), .A2(n665), .ZN(n529) );
  XNOR2_X1 U642 ( .A(n530), .B(n529), .ZN(n532) );
  XNOR2_X1 U643 ( .A(n534), .B(KEYINPUT109), .ZN(n730) );
  NOR2_X1 U644 ( .A1(n535), .A2(n657), .ZN(n537) );
  XNOR2_X1 U645 ( .A(KEYINPUT110), .B(KEYINPUT28), .ZN(n536) );
  XNOR2_X1 U646 ( .A(n537), .B(n536), .ZN(n538) );
  NAND2_X1 U647 ( .A1(n394), .A2(n538), .ZN(n553) );
  XNOR2_X1 U648 ( .A(KEYINPUT79), .B(KEYINPUT19), .ZN(n540) );
  XNOR2_X1 U649 ( .A(n540), .B(KEYINPUT67), .ZN(n541) );
  NOR2_X1 U650 ( .A1(n552), .A2(n542), .ZN(n645) );
  NOR2_X1 U651 ( .A1(n645), .A2(n559), .ZN(n543) );
  XNOR2_X1 U652 ( .A(n543), .B(KEYINPUT105), .ZN(n594) );
  NOR2_X1 U653 ( .A1(KEYINPUT47), .A2(n544), .ZN(n545) );
  XNOR2_X1 U654 ( .A(n548), .B(n547), .ZN(n562) );
  XNOR2_X1 U655 ( .A(KEYINPUT38), .B(KEYINPUT77), .ZN(n549) );
  NAND2_X1 U656 ( .A1(n664), .A2(n665), .ZN(n550) );
  NAND2_X1 U657 ( .A1(n552), .A2(n551), .ZN(n667) );
  XNOR2_X1 U658 ( .A(KEYINPUT113), .B(KEYINPUT42), .ZN(n554) );
  XOR2_X1 U659 ( .A(KEYINPUT111), .B(KEYINPUT40), .Z(n560) );
  INV_X1 U660 ( .A(n664), .ZN(n556) );
  XNOR2_X1 U661 ( .A(KEYINPUT89), .B(KEYINPUT39), .ZN(n558) );
  NOR2_X1 U662 ( .A1(n562), .A2(n561), .ZN(n568) );
  XNOR2_X1 U663 ( .A(KEYINPUT36), .B(n565), .ZN(n566) );
  NAND2_X1 U664 ( .A1(n566), .A2(n398), .ZN(n567) );
  XNOR2_X1 U665 ( .A(n567), .B(KEYINPUT114), .ZN(n732) );
  NAND2_X1 U666 ( .A1(n568), .A2(n732), .ZN(n569) );
  NAND2_X1 U667 ( .A1(n570), .A2(n645), .ZN(n648) );
  NOR2_X1 U668 ( .A1(G898), .A2(n726), .ZN(n716) );
  INV_X1 U669 ( .A(n571), .ZN(n572) );
  NAND2_X1 U670 ( .A1(n716), .A2(n572), .ZN(n574) );
  NAND2_X1 U671 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U672 ( .A(KEYINPUT68), .B(KEYINPUT0), .Z(n577) );
  NOR2_X1 U673 ( .A1(n667), .A2(n651), .ZN(n579) );
  INV_X1 U674 ( .A(KEYINPUT35), .ZN(n586) );
  INV_X1 U675 ( .A(n652), .ZN(n591) );
  INV_X1 U676 ( .A(n398), .ZN(n593) );
  NOR2_X1 U677 ( .A1(n591), .A2(n593), .ZN(n589) );
  NAND2_X1 U678 ( .A1(n593), .A2(n592), .ZN(n629) );
  INV_X1 U679 ( .A(n594), .ZN(n668) );
  NAND2_X1 U680 ( .A1(n391), .A2(n595), .ZN(n596) );
  NOR2_X1 U681 ( .A1(n597), .A2(n596), .ZN(n631) );
  NOR2_X1 U682 ( .A1(n657), .A2(n598), .ZN(n661) );
  NAND2_X1 U683 ( .A1(n661), .A2(n391), .ZN(n600) );
  XNOR2_X1 U684 ( .A(n600), .B(KEYINPUT31), .ZN(n646) );
  NOR2_X1 U685 ( .A1(n631), .A2(n646), .ZN(n601) );
  NOR2_X1 U686 ( .A1(n668), .A2(n601), .ZN(n602) );
  XNOR2_X1 U687 ( .A(KEYINPUT85), .B(KEYINPUT45), .ZN(n608) );
  INV_X1 U688 ( .A(n610), .ZN(n609) );
  NOR2_X1 U689 ( .A1(KEYINPUT84), .A2(n610), .ZN(n611) );
  NOR2_X1 U690 ( .A1(G952), .A2(n726), .ZN(n616) );
  NOR2_X1 U691 ( .A1(n617), .A2(n706), .ZN(G54) );
  XNOR2_X1 U692 ( .A(n618), .B(n619), .ZN(n620) );
  NOR2_X2 U693 ( .A1(n620), .A2(n706), .ZN(n621) );
  XNOR2_X1 U694 ( .A(n621), .B(KEYINPUT124), .ZN(G63) );
  XOR2_X1 U695 ( .A(KEYINPUT62), .B(KEYINPUT115), .Z(n622) );
  XNOR2_X1 U696 ( .A(n625), .B(n624), .ZN(n626) );
  NOR2_X2 U697 ( .A1(n626), .A2(n706), .ZN(n628) );
  XNOR2_X1 U698 ( .A(n628), .B(n627), .ZN(G57) );
  XNOR2_X1 U699 ( .A(G101), .B(n629), .ZN(G3) );
  NAND2_X1 U700 ( .A1(n631), .A2(n642), .ZN(n630) );
  XNOR2_X1 U701 ( .A(n630), .B(n401), .ZN(G6) );
  XOR2_X1 U702 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n633) );
  NAND2_X1 U703 ( .A1(n631), .A2(n645), .ZN(n632) );
  XNOR2_X1 U704 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U705 ( .A(G107), .B(n634), .ZN(G9) );
  XOR2_X1 U706 ( .A(n635), .B(G110), .Z(G12) );
  XOR2_X1 U707 ( .A(KEYINPUT117), .B(KEYINPUT29), .Z(n637) );
  NAND2_X1 U708 ( .A1(n640), .A2(n645), .ZN(n636) );
  XNOR2_X1 U709 ( .A(n637), .B(n636), .ZN(n639) );
  XOR2_X1 U710 ( .A(G128), .B(KEYINPUT116), .Z(n638) );
  XNOR2_X1 U711 ( .A(n639), .B(n638), .ZN(G30) );
  NAND2_X1 U712 ( .A1(n640), .A2(n642), .ZN(n641) );
  XNOR2_X1 U713 ( .A(n641), .B(G146), .ZN(G48) );
  NAND2_X1 U714 ( .A1(n646), .A2(n642), .ZN(n643) );
  XNOR2_X1 U715 ( .A(n643), .B(KEYINPUT118), .ZN(n644) );
  XNOR2_X1 U716 ( .A(G113), .B(n644), .ZN(G15) );
  NAND2_X1 U717 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U718 ( .A(n647), .B(G116), .ZN(G18) );
  XNOR2_X1 U719 ( .A(G134), .B(n648), .ZN(G36) );
  XOR2_X1 U720 ( .A(G140), .B(n649), .Z(G42) );
  NAND2_X1 U721 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U722 ( .A(n653), .B(KEYINPUT49), .ZN(n659) );
  NOR2_X1 U723 ( .A1(n654), .A2(n398), .ZN(n655) );
  XOR2_X1 U724 ( .A(KEYINPUT50), .B(n655), .Z(n656) );
  NAND2_X1 U725 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U726 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U727 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U728 ( .A(KEYINPUT51), .B(n662), .Z(n663) );
  NOR2_X1 U729 ( .A1(n681), .A2(n663), .ZN(n674) );
  NOR2_X1 U730 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U731 ( .A1(n667), .A2(n666), .ZN(n671) );
  NOR2_X1 U732 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U733 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U734 ( .A1(n672), .A2(n680), .ZN(n673) );
  NOR2_X1 U735 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U736 ( .A(n675), .B(KEYINPUT52), .Z(n676) );
  XNOR2_X1 U737 ( .A(KEYINPUT119), .B(n676), .ZN(n677) );
  NOR2_X1 U738 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U739 ( .A(n679), .B(KEYINPUT120), .ZN(n683) );
  NOR2_X1 U740 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U741 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U742 ( .A(KEYINPUT121), .B(n684), .Z(n687) );
  XNOR2_X1 U743 ( .A(KEYINPUT2), .B(n392), .ZN(n686) );
  NAND2_X1 U744 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U745 ( .A1(n688), .A2(G953), .ZN(n689) );
  XNOR2_X1 U746 ( .A(n689), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U747 ( .A(n692), .B(n691), .ZN(n693) );
  NOR2_X2 U748 ( .A1(n693), .A2(n706), .ZN(n695) );
  XOR2_X1 U749 ( .A(KEYINPUT87), .B(KEYINPUT56), .Z(n694) );
  XNOR2_X1 U750 ( .A(n695), .B(n694), .ZN(G51) );
  XOR2_X1 U751 ( .A(KEYINPUT122), .B(KEYINPUT59), .Z(n696) );
  XNOR2_X1 U752 ( .A(n699), .B(n698), .ZN(n700) );
  NOR2_X2 U753 ( .A1(n700), .A2(n706), .ZN(n702) );
  XOR2_X1 U754 ( .A(KEYINPUT60), .B(KEYINPUT123), .Z(n701) );
  XNOR2_X1 U755 ( .A(n702), .B(n701), .ZN(G60) );
  XNOR2_X1 U756 ( .A(n704), .B(n703), .ZN(n705) );
  NOR2_X1 U757 ( .A1(n706), .A2(n705), .ZN(G66) );
  NAND2_X1 U758 ( .A1(G953), .A2(G224), .ZN(n707) );
  XNOR2_X1 U759 ( .A(KEYINPUT61), .B(n707), .ZN(n708) );
  AND2_X1 U760 ( .A1(n708), .A2(G898), .ZN(n711) );
  NOR2_X1 U761 ( .A1(G953), .A2(n393), .ZN(n710) );
  NOR2_X1 U762 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U763 ( .A(n712), .B(KEYINPUT125), .ZN(n718) );
  XOR2_X1 U764 ( .A(n714), .B(n713), .Z(n715) );
  NOR2_X1 U765 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U766 ( .A(n718), .B(n717), .ZN(G69) );
  XOR2_X1 U767 ( .A(n719), .B(n720), .Z(n725) );
  XNOR2_X1 U768 ( .A(G227), .B(n725), .ZN(n721) );
  NAND2_X1 U769 ( .A1(n721), .A2(G900), .ZN(n722) );
  NAND2_X1 U770 ( .A1(G953), .A2(n722), .ZN(n723) );
  XNOR2_X1 U771 ( .A(n723), .B(KEYINPUT126), .ZN(n729) );
  XNOR2_X1 U772 ( .A(n725), .B(n724), .ZN(n727) );
  NAND2_X1 U773 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U774 ( .A1(n729), .A2(n728), .ZN(G72) );
  XNOR2_X1 U775 ( .A(G143), .B(n730), .ZN(G45) );
  XOR2_X1 U776 ( .A(n344), .B(G122), .Z(G24) );
  XOR2_X1 U777 ( .A(G125), .B(n732), .Z(n733) );
  XNOR2_X1 U778 ( .A(KEYINPUT37), .B(n733), .ZN(G27) );
  XOR2_X1 U779 ( .A(G119), .B(n734), .Z(n735) );
  XNOR2_X1 U780 ( .A(KEYINPUT127), .B(n735), .ZN(G21) );
  XNOR2_X1 U781 ( .A(G137), .B(n736), .ZN(G39) );
  XNOR2_X1 U782 ( .A(G131), .B(n737), .ZN(G33) );
endmodule

