//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 1 0 0 1 0 1 1 0 0 1 1 1 0 1 1 0 1 1 0 0 1 1 0 1 0 0 0 1 1 0 1 1 1 0 0 1 0 0 1 1 0 1 1 0 0 0 1 1 1 0 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1280, new_n1281, new_n1282, new_n1283, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1331, new_n1332, new_n1333, new_n1334;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n201), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT64), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT65), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n226), .B1(new_n222), .B2(new_n223), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n209), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n212), .B1(new_n215), .B2(new_n217), .C1(new_n228), .C2(KEYINPUT1), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT66), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n202), .A2(G68), .ZN(new_n243));
  INV_X1    g0043(.A(G68), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(G50), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n242), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G274), .ZN(new_n250));
  AND2_X1   g0050(.A1(G1), .A2(G13), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G33), .A2(G41), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G238), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n251), .A2(new_n252), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n254), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n256), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G226), .ZN(new_n261));
  INV_X1    g0061(.A(G1698), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G232), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G1698), .ZN(new_n265));
  AND2_X1   g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NOR2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n263), .B(new_n265), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G97), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n258), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(KEYINPUT13), .B1(new_n260), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n268), .A2(new_n269), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT13), .ZN(new_n275));
  INV_X1    g0075(.A(G41), .ZN(new_n276));
  INV_X1    g0076(.A(G45), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n206), .A2(new_n278), .B1(new_n251), .B2(new_n252), .ZN(new_n279));
  AOI22_X1  g0079(.A1(new_n279), .A2(G238), .B1(new_n253), .B2(new_n255), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n274), .A2(new_n275), .A3(new_n280), .ZN(new_n281));
  AND3_X1   g0081(.A1(new_n271), .A2(G179), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT71), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n271), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n274), .A2(new_n280), .A3(KEYINPUT71), .A4(new_n275), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n284), .A2(G169), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n282), .B1(new_n286), .B2(KEYINPUT14), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT14), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n284), .A2(new_n288), .A3(G169), .A4(new_n285), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n213), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G20), .A2(G33), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  OAI22_X1  g0094(.A1(new_n294), .A2(new_n202), .B1(new_n207), .B2(G68), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n207), .A2(G33), .ZN(new_n296));
  INV_X1    g0096(.A(G77), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n292), .B1(new_n295), .B2(new_n298), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n299), .A2(KEYINPUT72), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(KEYINPUT72), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT11), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT11), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n300), .A2(new_n304), .A3(new_n301), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n306), .A2(G68), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n307), .B(KEYINPUT12), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT67), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n309), .B1(new_n207), .B2(G1), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n206), .A2(KEYINPUT67), .A3(G20), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G68), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n306), .A2(new_n213), .A3(new_n291), .ZN(new_n314));
  OR3_X1    g0114(.A1(new_n313), .A2(KEYINPUT73), .A3(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT73), .B1(new_n313), .B2(new_n314), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n308), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n303), .A2(new_n305), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n290), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n271), .A2(new_n281), .A3(G190), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n303), .A2(new_n305), .A3(new_n320), .A4(new_n317), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n284), .A2(G200), .A3(new_n285), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  OR2_X1    g0126(.A1(KEYINPUT3), .A2(G33), .ZN(new_n327));
  NAND2_X1  g0127(.A1(KEYINPUT3), .A2(G33), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n329), .A2(G222), .A3(new_n262), .ZN(new_n330));
  OAI211_X1 g0130(.A(G223), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n266), .A2(new_n267), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(G77), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n330), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n273), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n256), .B1(new_n259), .B2(new_n261), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G169), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n203), .A2(G20), .ZN(new_n341));
  INV_X1    g0141(.A(G150), .ZN(new_n342));
  XNOR2_X1  g0142(.A(KEYINPUT8), .B(G58), .ZN(new_n343));
  OAI221_X1 g0143(.A(new_n341), .B1(new_n342), .B2(new_n294), .C1(new_n296), .C2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n306), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n344), .A2(new_n292), .B1(new_n202), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n312), .A2(G50), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT68), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n314), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n312), .A2(KEYINPUT68), .A3(G50), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n346), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n336), .B1(new_n273), .B2(new_n334), .ZN(new_n354));
  INV_X1    g0154(.A(G179), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n340), .A2(new_n353), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT9), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n343), .A2(new_n296), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n207), .B1(new_n201), .B2(new_n202), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n294), .A2(new_n342), .ZN(new_n362));
  NOR3_X1   g0162(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n292), .ZN(new_n364));
  OAI22_X1  g0164(.A1(new_n363), .A2(new_n364), .B1(G50), .B2(new_n306), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n359), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(KEYINPUT10), .B1(new_n354), .B2(G190), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n346), .A2(KEYINPUT9), .A3(new_n352), .ZN(new_n369));
  AND3_X1   g0169(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT70), .ZN(new_n371));
  INV_X1    g0171(.A(G200), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n371), .B1(new_n354), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n338), .A2(KEYINPUT70), .A3(G200), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n370), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n354), .A2(G190), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n338), .A2(G200), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n367), .A2(new_n369), .A3(new_n377), .A4(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT10), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n358), .B1(new_n376), .B2(new_n380), .ZN(new_n381));
  XOR2_X1   g0181(.A(KEYINPUT8), .B(G58), .Z(new_n382));
  AOI22_X1  g0182(.A1(new_n382), .A2(new_n293), .B1(G20), .B2(G77), .ZN(new_n383));
  XNOR2_X1  g0183(.A(KEYINPUT15), .B(G87), .ZN(new_n384));
  OR2_X1    g0184(.A1(new_n384), .A2(new_n296), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n364), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n312), .A2(G77), .ZN(new_n387));
  OAI22_X1  g0187(.A1(new_n387), .A2(new_n314), .B1(G77), .B2(new_n306), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(G244), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n256), .B1(new_n259), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n329), .A2(G238), .A3(G1698), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n329), .A2(G232), .A3(new_n262), .ZN(new_n394));
  INV_X1    g0194(.A(G107), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n393), .B(new_n394), .C1(new_n395), .C2(new_n329), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n392), .B1(new_n396), .B2(new_n273), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n390), .B1(G169), .B2(new_n397), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n397), .A2(new_n355), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n389), .B1(new_n397), .B2(new_n372), .ZN(new_n401));
  OR2_X1    g0201(.A1(new_n401), .A2(KEYINPUT69), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n401), .A2(KEYINPUT69), .B1(G190), .B2(new_n397), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n400), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n381), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n343), .B1(new_n310), .B2(new_n311), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n406), .A2(new_n350), .B1(new_n345), .B2(new_n343), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT7), .B1(new_n332), .B2(new_n207), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT7), .ZN(new_n410));
  NOR4_X1   g0210(.A1(new_n266), .A2(new_n267), .A3(new_n410), .A4(G20), .ZN(new_n411));
  OAI21_X1  g0211(.A(G68), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(G58), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n413), .A2(new_n244), .ZN(new_n414));
  OAI21_X1  g0214(.A(G20), .B1(new_n414), .B2(new_n201), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n293), .A2(G159), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n412), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT16), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n364), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n412), .A2(KEYINPUT16), .A3(new_n418), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n408), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OR2_X1    g0223(.A1(G223), .A2(G1698), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n261), .A2(G1698), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n424), .B(new_n425), .C1(new_n266), .C2(new_n267), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G33), .A2(G87), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n273), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n279), .A2(G232), .B1(new_n253), .B2(new_n255), .ZN(new_n430));
  AOI21_X1  g0230(.A(G169), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n258), .A2(G232), .A3(new_n254), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n256), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n258), .B1(new_n426), .B2(new_n427), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(KEYINPUT74), .B1(new_n436), .B2(new_n355), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n429), .A2(new_n430), .A3(KEYINPUT74), .A4(new_n355), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n432), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT18), .B1(new_n423), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n327), .A2(new_n207), .A3(new_n328), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n410), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n327), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n328), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n244), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n420), .B1(new_n445), .B2(new_n417), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n446), .A2(new_n422), .A3(new_n292), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n407), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n429), .A2(new_n355), .A3(new_n430), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT74), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n431), .B1(new_n451), .B2(new_n438), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT18), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n448), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(G190), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n436), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n372), .B1(new_n434), .B2(new_n435), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n447), .A2(new_n458), .A3(new_n407), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT17), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n447), .A2(new_n458), .A3(KEYINPUT17), .A4(new_n407), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n441), .A2(new_n454), .A3(new_n461), .A4(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n326), .A2(new_n405), .A3(KEYINPUT75), .A4(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT75), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n464), .A2(new_n381), .A3(new_n404), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n466), .B1(new_n467), .B2(new_n325), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G283), .ZN(new_n470));
  INV_X1    g0270(.A(G97), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n470), .B(new_n207), .C1(G33), .C2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(G116), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G20), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n472), .A2(new_n292), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT20), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n472), .A2(KEYINPUT20), .A3(new_n292), .A4(new_n474), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n306), .A2(G116), .ZN(new_n480));
  INV_X1    g0280(.A(G33), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n481), .A2(G1), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n314), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n480), .B1(new_n483), .B2(G116), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n479), .A2(new_n484), .ZN(new_n485));
  OAI211_X1 g0285(.A(G257), .B(new_n262), .C1(new_n266), .C2(new_n267), .ZN(new_n486));
  OAI211_X1 g0286(.A(G264), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n487));
  XOR2_X1   g0287(.A(KEYINPUT81), .B(G303), .Z(new_n488));
  OAI211_X1 g0288(.A(new_n486), .B(new_n487), .C1(new_n488), .C2(new_n329), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n355), .B1(new_n489), .B2(new_n273), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n485), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n277), .A2(G1), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT77), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n494), .A2(new_n276), .A3(KEYINPUT5), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT5), .ZN(new_n496));
  AOI21_X1  g0296(.A(KEYINPUT77), .B1(new_n496), .B2(G41), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n496), .A2(G41), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n493), .B(new_n495), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n499), .A2(KEYINPUT80), .A3(G270), .A4(new_n258), .ZN(new_n500));
  AND2_X1   g0300(.A1(new_n495), .A2(new_n493), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n494), .B1(new_n276), .B2(KEYINPUT5), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(new_n496), .B2(G41), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n501), .A2(new_n503), .A3(new_n253), .ZN(new_n504));
  AND2_X1   g0304(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n499), .A2(G270), .A3(new_n258), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT80), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n492), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n489), .A2(new_n273), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n508), .A2(new_n511), .A3(new_n504), .A4(new_n500), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n339), .B1(new_n479), .B2(new_n484), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT21), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n514), .B1(new_n512), .B2(new_n513), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n510), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n512), .A2(G200), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n485), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n512), .A2(new_n455), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(KEYINPUT82), .B1(new_n517), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n512), .A2(new_n513), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(KEYINPUT21), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT82), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n518), .B(new_n485), .C1(new_n455), .C2(new_n512), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n526), .A2(new_n527), .A3(new_n528), .A4(new_n510), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n522), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n273), .B1(new_n501), .B2(new_n503), .ZN(new_n531));
  OAI211_X1 g0331(.A(G257), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n532));
  OAI211_X1 g0332(.A(G250), .B(new_n262), .C1(new_n266), .C2(new_n267), .ZN(new_n533));
  INV_X1    g0333(.A(G294), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n532), .B(new_n533), .C1(new_n481), .C2(new_n534), .ZN(new_n535));
  AOI22_X1  g0335(.A1(G264), .A2(new_n531), .B1(new_n535), .B2(new_n273), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n536), .A2(new_n355), .A3(new_n504), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(new_n273), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n499), .A2(G264), .A3(new_n258), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n538), .A2(new_n504), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n339), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT23), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n544), .A2(new_n395), .A3(G20), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT83), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G33), .A2(G116), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n547), .B1(new_n548), .B2(G20), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n207), .A2(KEYINPUT83), .A3(G33), .A4(G116), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n546), .A2(KEYINPUT84), .A3(new_n549), .A4(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n549), .A2(new_n550), .A3(new_n545), .A4(new_n543), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT84), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n207), .B(G87), .C1(new_n266), .C2(new_n267), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(KEYINPUT22), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT22), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n329), .A2(new_n558), .A3(new_n207), .A4(G87), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n557), .A2(new_n559), .B1(KEYINPUT85), .B2(KEYINPUT24), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(KEYINPUT85), .A2(KEYINPUT24), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n555), .A2(new_n560), .A3(new_n562), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n364), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OR2_X1    g0366(.A1(new_n314), .A2(new_n482), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n567), .A2(new_n395), .ZN(new_n568));
  XOR2_X1   g0368(.A(KEYINPUT86), .B(KEYINPUT25), .Z(new_n569));
  NOR2_X1   g0369(.A1(new_n306), .A2(G107), .ZN(new_n570));
  XNOR2_X1  g0370(.A(new_n569), .B(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n542), .B1(new_n566), .B2(new_n573), .ZN(new_n574));
  AND3_X1   g0374(.A1(new_n555), .A2(new_n560), .A3(new_n562), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n562), .B1(new_n555), .B2(new_n560), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n292), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n540), .A2(new_n372), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n538), .A2(new_n455), .A3(new_n504), .A4(new_n539), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n577), .A2(new_n572), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n574), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g0382(.A(G97), .B(G107), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT6), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n584), .A2(new_n471), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n583), .A2(new_n584), .B1(new_n395), .B2(new_n585), .ZN(new_n586));
  OAI22_X1  g0386(.A1(new_n586), .A2(new_n207), .B1(new_n297), .B2(new_n294), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n395), .B1(new_n443), .B2(new_n444), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n292), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n306), .A2(G97), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(new_n567), .B2(new_n471), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(G244), .B(new_n262), .C1(new_n266), .C2(new_n267), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT76), .ZN(new_n596));
  OR2_X1    g0396(.A1(new_n596), .A2(KEYINPUT4), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n329), .A2(G244), .A3(new_n262), .A4(new_n597), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n329), .A2(G250), .A3(G1698), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n599), .A2(new_n600), .A3(new_n470), .A4(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n273), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n499), .A2(G257), .A3(new_n258), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n604), .A2(new_n504), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n603), .A2(new_n605), .A3(new_n355), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(new_n504), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n607), .B1(new_n273), .B2(new_n602), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n594), .B(new_n606), .C1(G169), .C2(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(G107), .B1(new_n409), .B2(new_n411), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n294), .A2(new_n297), .ZN(new_n611));
  AND2_X1   g0411(.A1(G97), .A2(G107), .ZN(new_n612));
  NOR2_X1   g0412(.A1(G97), .A2(G107), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n584), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n395), .A2(KEYINPUT6), .A3(G97), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n611), .B1(new_n616), .B2(G20), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n610), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n592), .B1(new_n618), .B2(new_n292), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n603), .A2(new_n605), .A3(G190), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n619), .B(new_n620), .C1(new_n608), .C2(new_n372), .ZN(new_n621));
  OAI211_X1 g0421(.A(G238), .B(new_n262), .C1(new_n266), .C2(new_n267), .ZN(new_n622));
  OAI211_X1 g0422(.A(G244), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n622), .A2(new_n623), .A3(new_n548), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n273), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n253), .A2(new_n493), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT78), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n627), .A2(new_n206), .A3(G45), .ZN(new_n628));
  OAI21_X1  g0428(.A(KEYINPUT78), .B1(new_n277), .B2(G1), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n258), .A2(G250), .A3(new_n628), .A4(new_n629), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n372), .B1(new_n625), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT19), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n207), .B1(new_n269), .B2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(G87), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n613), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n207), .B(G68), .C1(new_n266), .C2(new_n267), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n634), .B1(new_n296), .B2(new_n471), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n641), .A2(new_n292), .B1(new_n345), .B2(new_n384), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n483), .A2(G87), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n626), .A2(new_n630), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n645), .B1(new_n273), .B2(new_n624), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(G190), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n633), .A2(new_n644), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n625), .A2(new_n631), .ZN(new_n649));
  OR3_X1    g0449(.A1(new_n314), .A2(new_n384), .A3(new_n482), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n649), .A2(new_n339), .B1(new_n642), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT79), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n649), .B2(G179), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n646), .A2(KEYINPUT79), .A3(new_n355), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n651), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n609), .A2(new_n621), .A3(new_n648), .A4(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n582), .A2(new_n656), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n469), .A2(new_n530), .A3(new_n657), .ZN(G372));
  NAND2_X1  g0458(.A1(new_n655), .A2(new_n648), .ZN(new_n659));
  OAI21_X1  g0459(.A(KEYINPUT26), .B1(new_n659), .B2(new_n609), .ZN(new_n660));
  INV_X1    g0460(.A(new_n609), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT26), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n625), .A2(new_n631), .A3(G190), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n663), .A2(new_n632), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n646), .A2(new_n355), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n664), .A2(new_n644), .B1(new_n651), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n661), .A2(new_n662), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n651), .A2(new_n665), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT88), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n668), .B(new_n669), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n660), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  AOI22_X1  g0471(.A1(new_n524), .A2(new_n525), .B1(new_n509), .B2(new_n492), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n574), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n581), .A2(new_n609), .A3(new_n666), .A4(new_n621), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n673), .B1(new_n674), .B2(KEYINPUT87), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT87), .ZN(new_n676));
  AND4_X1   g0476(.A1(new_n609), .A2(new_n621), .A3(new_n648), .A4(new_n668), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n676), .B1(new_n677), .B2(new_n581), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n671), .B1(new_n675), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n469), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT89), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n448), .A2(new_n453), .A3(new_n452), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n453), .B1(new_n448), .B2(new_n452), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n441), .A2(KEYINPUT89), .A3(new_n454), .ZN(new_n685));
  AOI22_X1  g0485(.A1(new_n324), .A2(new_n400), .B1(new_n290), .B2(new_n318), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n461), .A2(new_n462), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n684), .B(new_n685), .C1(new_n686), .C2(new_n687), .ZN(new_n688));
  AOI22_X1  g0488(.A1(new_n370), .A2(new_n375), .B1(new_n379), .B2(KEYINPUT10), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n358), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n680), .A2(new_n691), .ZN(G369));
  NAND3_X1  g0492(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n694));
  XOR2_X1   g0494(.A(new_n694), .B(KEYINPUT90), .Z(new_n695));
  INV_X1    g0495(.A(G213), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n696), .B1(new_n693), .B2(KEYINPUT27), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(G343), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n530), .B1(new_n485), .B2(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n485), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n517), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT91), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(G330), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n700), .B1(new_n566), .B2(new_n573), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n574), .A2(new_n709), .A3(new_n581), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n574), .B2(new_n701), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n574), .A2(new_n700), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n672), .A2(new_n700), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(new_n710), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n712), .A2(new_n713), .A3(new_n717), .ZN(G399));
  INV_X1    g0518(.A(new_n210), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(G41), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n637), .A2(G116), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n721), .A2(G1), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(new_n217), .B2(new_n721), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT28), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n674), .B1(new_n672), .B2(new_n574), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n661), .A2(new_n662), .A3(new_n648), .A4(new_n655), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n668), .A2(new_n648), .ZN(new_n728));
  OAI21_X1  g0528(.A(KEYINPUT26), .B1(new_n728), .B2(new_n609), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n727), .A2(new_n670), .A3(new_n729), .ZN(new_n730));
  OAI211_X1 g0530(.A(KEYINPUT29), .B(new_n701), .C1(new_n726), .C2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n674), .A2(KEYINPUT87), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n609), .A2(new_n621), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n733), .A2(new_n676), .A3(new_n581), .A4(new_n666), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n732), .A2(new_n734), .A3(new_n673), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n700), .B1(new_n735), .B2(new_n671), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n731), .B1(new_n736), .B2(KEYINPUT29), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n536), .A2(new_n646), .A3(new_n490), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT92), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT30), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n738), .A2(new_n509), .A3(new_n608), .A4(new_n741), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n603), .A2(new_n505), .A3(new_n508), .A4(new_n605), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n536), .A2(new_n646), .A3(new_n490), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n739), .B(new_n740), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n646), .A2(G179), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT93), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n746), .A2(new_n747), .A3(new_n512), .ZN(new_n748));
  AOI22_X1  g0548(.A1(new_n504), .A2(new_n536), .B1(new_n603), .B2(new_n605), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n747), .B1(new_n746), .B2(new_n512), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n742), .B(new_n745), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n752), .A2(KEYINPUT31), .A3(new_n700), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(KEYINPUT94), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT94), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n752), .A2(new_n755), .A3(KEYINPUT31), .A4(new_n700), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n752), .A2(new_n700), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT31), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n754), .A2(new_n756), .A3(new_n759), .ZN(new_n760));
  AND3_X1   g0560(.A1(new_n530), .A2(new_n657), .A3(new_n701), .ZN(new_n761));
  OAI21_X1  g0561(.A(G330), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n737), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n725), .B1(new_n764), .B2(G1), .ZN(G364));
  INV_X1    g0565(.A(G13), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n206), .B1(new_n767), .B2(G45), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n720), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n708), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(G330), .B2(new_n706), .ZN(new_n772));
  INV_X1    g0572(.A(new_n770), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n210), .A2(G355), .A3(new_n329), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n719), .A2(new_n329), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n775), .B1(G45), .B2(new_n217), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n248), .A2(new_n277), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n774), .B1(G116), .B2(new_n210), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  OR3_X1    g0578(.A1(KEYINPUT95), .A2(G13), .A3(G33), .ZN(new_n779));
  OAI21_X1  g0579(.A(KEYINPUT95), .B1(G13), .B2(G33), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(G20), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n213), .B1(G20), .B2(new_n339), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n773), .B1(new_n778), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n784), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n207), .A2(G179), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n788), .A2(new_n455), .A3(G200), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n395), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n788), .A2(G190), .A3(G200), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n636), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n790), .A2(new_n792), .A3(new_n332), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n793), .B(KEYINPUT96), .Z(new_n794));
  NOR2_X1   g0594(.A1(new_n207), .A2(new_n355), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G190), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(G200), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(G58), .ZN(new_n798));
  NOR3_X1   g0598(.A1(new_n455), .A2(G179), .A3(G200), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(new_n207), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(G97), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n796), .A2(new_n372), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G50), .ZN(new_n804));
  NOR2_X1   g0604(.A1(G190), .A2(G200), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n788), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G159), .ZN(new_n807));
  OAI21_X1  g0607(.A(KEYINPUT32), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n798), .A2(new_n802), .A3(new_n804), .A4(new_n808), .ZN(new_n809));
  NOR3_X1   g0609(.A1(new_n806), .A2(KEYINPUT32), .A3(new_n807), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n795), .A2(new_n455), .A3(G200), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n795), .A2(new_n805), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n811), .A2(new_n244), .B1(new_n812), .B2(new_n297), .ZN(new_n813));
  NOR3_X1   g0613(.A1(new_n809), .A2(new_n810), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n797), .A2(G322), .ZN(new_n815));
  INV_X1    g0615(.A(G283), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n815), .B1(new_n816), .B2(new_n789), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(G294), .B2(new_n801), .ZN(new_n818));
  INV_X1    g0618(.A(new_n791), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n803), .A2(G326), .B1(new_n819), .B2(G303), .ZN(new_n820));
  INV_X1    g0620(.A(new_n811), .ZN(new_n821));
  XNOR2_X1  g0621(.A(KEYINPUT33), .B(G317), .ZN(new_n822));
  INV_X1    g0622(.A(new_n812), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n821), .A2(new_n822), .B1(new_n823), .B2(G311), .ZN(new_n824));
  INV_X1    g0624(.A(new_n806), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n329), .B1(new_n825), .B2(G329), .ZN(new_n826));
  AND3_X1   g0626(.A1(new_n820), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n794), .A2(new_n814), .B1(new_n818), .B2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n783), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n786), .B1(new_n787), .B2(new_n828), .C1(new_n706), .C2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n772), .A2(new_n830), .ZN(G396));
  NAND2_X1  g0631(.A1(new_n400), .A2(new_n701), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n402), .A2(new_n403), .B1(new_n390), .B2(new_n700), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n832), .B1(new_n833), .B2(new_n400), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n736), .B(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n770), .B1(new_n836), .B2(new_n762), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n762), .B2(new_n836), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n781), .A2(new_n784), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n773), .B1(new_n297), .B2(new_n839), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n821), .A2(G150), .B1(new_n823), .B2(G159), .ZN(new_n841));
  INV_X1    g0641(.A(new_n797), .ZN(new_n842));
  INV_X1    g0642(.A(G143), .ZN(new_n843));
  INV_X1    g0643(.A(G137), .ZN(new_n844));
  INV_X1    g0644(.A(new_n803), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n841), .B1(new_n842), .B2(new_n843), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT34), .ZN(new_n847));
  OR2_X1    g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n847), .ZN(new_n849));
  INV_X1    g0649(.A(G132), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n329), .B1(new_n806), .B2(new_n850), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n851), .B(KEYINPUT97), .Z(new_n852));
  OAI22_X1  g0652(.A1(new_n800), .A2(new_n413), .B1(new_n791), .B2(new_n202), .ZN(new_n853));
  INV_X1    g0653(.A(new_n789), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n853), .B1(G68), .B2(new_n854), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n848), .A2(new_n849), .A3(new_n852), .A4(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(G303), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n842), .A2(new_n534), .B1(new_n845), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(G107), .B2(new_n819), .ZN(new_n859));
  INV_X1    g0659(.A(G311), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n812), .A2(new_n473), .B1(new_n806), .B2(new_n860), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n329), .B(new_n861), .C1(G283), .C2(new_n821), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n789), .A2(new_n636), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n859), .A2(new_n802), .A3(new_n862), .A4(new_n864), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n856), .A2(new_n865), .ZN(new_n866));
  OAI221_X1 g0666(.A(new_n840), .B1(new_n787), .B2(new_n866), .C1(new_n835), .C2(new_n782), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n838), .A2(new_n867), .ZN(G384));
  NOR2_X1   g0668(.A1(new_n767), .A2(new_n206), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT39), .ZN(new_n870));
  INV_X1    g0670(.A(new_n687), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n684), .A2(new_n871), .A3(new_n685), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n423), .A2(new_n698), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n459), .B1(new_n423), .B2(new_n440), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT99), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT37), .ZN(new_n878));
  INV_X1    g0678(.A(new_n698), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n448), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n876), .A2(new_n877), .A3(new_n878), .A4(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT37), .B1(new_n875), .B2(new_n873), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n448), .A2(new_n452), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n883), .A2(new_n880), .A3(new_n878), .A4(new_n459), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(KEYINPUT99), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n881), .A2(new_n882), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT38), .B1(new_n874), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n882), .A2(new_n884), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n463), .A2(new_n873), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n888), .A2(new_n889), .A3(KEYINPUT38), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n870), .B1(new_n887), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n319), .A2(new_n700), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n888), .A2(new_n889), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT38), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n888), .A2(new_n889), .A3(KEYINPUT38), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n895), .A2(KEYINPUT39), .A3(new_n896), .ZN(new_n897));
  AND3_X1   g0697(.A1(new_n891), .A2(new_n892), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n895), .A2(new_n896), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n318), .A2(new_n700), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n319), .A2(new_n324), .A3(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n318), .B(new_n700), .C1(new_n290), .C2(new_n323), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI211_X1 g0703(.A(new_n700), .B(new_n834), .C1(new_n735), .C2(new_n671), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n832), .B(KEYINPUT98), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n899), .B(new_n903), .C1(new_n904), .C2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n684), .ZN(new_n908));
  INV_X1    g0708(.A(new_n685), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n698), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n898), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n469), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n691), .B1(new_n913), .B2(new_n737), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n912), .B(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(G330), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n874), .A2(new_n886), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n890), .B1(new_n917), .B2(new_n894), .ZN(new_n918));
  AND3_X1   g0718(.A1(new_n752), .A2(KEYINPUT31), .A3(new_n700), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT31), .B1(new_n752), .B2(new_n700), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n530), .A2(new_n657), .A3(new_n701), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n834), .B1(new_n901), .B2(new_n902), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(KEYINPUT40), .B1(new_n918), .B2(new_n925), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n923), .A2(new_n924), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT40), .B1(new_n895), .B2(new_n896), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n469), .A2(new_n923), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n916), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n931), .B2(new_n930), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n869), .B1(new_n915), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n915), .B2(new_n933), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n473), .B(new_n215), .C1(new_n616), .C2(KEYINPUT35), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(KEYINPUT35), .B2(new_n616), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT36), .ZN(new_n938));
  OAI21_X1  g0738(.A(G77), .B1(new_n413), .B2(new_n244), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n243), .B1(new_n217), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n940), .A2(G1), .A3(new_n766), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n935), .A2(new_n938), .A3(new_n941), .ZN(G367));
  INV_X1    g0742(.A(new_n775), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n785), .B1(new_n210), .B2(new_n384), .C1(new_n943), .C2(new_n238), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT105), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n773), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n945), .B2(new_n944), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n332), .B1(new_n812), .B2(new_n816), .ZN(new_n948));
  INV_X1    g0748(.A(G317), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n811), .A2(new_n534), .B1(new_n806), .B2(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n791), .A2(new_n473), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n948), .B(new_n950), .C1(KEYINPUT46), .C2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(KEYINPUT46), .B2(new_n951), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n845), .A2(new_n860), .B1(new_n395), .B2(new_n800), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n842), .A2(new_n488), .B1(new_n789), .B2(new_n471), .ZN(new_n955));
  NOR3_X1   g0755(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n800), .A2(new_n244), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(G150), .B2(new_n797), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT106), .ZN(new_n959));
  AOI22_X1  g0759(.A1(G50), .A2(new_n823), .B1(new_n825), .B2(G137), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n960), .B(new_n329), .C1(new_n807), .C2(new_n811), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n854), .A2(G77), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n962), .B1(new_n413), .B2(new_n791), .C1(new_n845), .C2(new_n843), .ZN(new_n963));
  NOR3_X1   g0763(.A1(new_n959), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n956), .A2(new_n964), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT47), .Z(new_n966));
  AOI21_X1  g0766(.A(new_n947), .B1(new_n966), .B2(new_n784), .ZN(new_n967));
  OR3_X1    g0767(.A1(new_n670), .A2(new_n644), .A3(new_n701), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n666), .B1(new_n644), .B2(new_n701), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n967), .B1(new_n829), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n733), .B1(new_n619), .B2(new_n701), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n661), .A2(new_n700), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n712), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n716), .A2(new_n974), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n978), .A2(KEYINPUT42), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT101), .Z(new_n980));
  OAI21_X1  g0780(.A(new_n609), .B1(new_n972), .B2(new_n574), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n978), .A2(KEYINPUT42), .B1(new_n701), .B2(new_n981), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n970), .A2(KEYINPUT100), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT43), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n970), .A2(KEYINPUT100), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n970), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n987), .B1(new_n985), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n983), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n987), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n990), .A2(KEYINPUT102), .B1(new_n983), .B2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n990), .A2(KEYINPUT102), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n977), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n992), .B(new_n976), .C1(KEYINPUT102), .C2(new_n990), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n768), .B(KEYINPUT104), .Z(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n712), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n717), .A2(new_n713), .ZN(new_n1001));
  AND3_X1   g0801(.A1(new_n1001), .A2(KEYINPUT44), .A3(new_n975), .ZN(new_n1002));
  AOI21_X1  g0802(.A(KEYINPUT44), .B1(new_n1001), .B2(new_n975), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n717), .A2(new_n713), .A3(new_n974), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT45), .ZN(new_n1006));
  OR3_X1    g0806(.A1(new_n1000), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1000), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT103), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n711), .A2(new_n714), .ZN(new_n1011));
  AND3_X1   g0811(.A1(new_n707), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n707), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n717), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  NOR3_X1   g0815(.A1(new_n1012), .A2(new_n1013), .A3(new_n717), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n764), .B1(new_n1009), .B2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n720), .B(KEYINPUT41), .Z(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n999), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n971), .B1(new_n997), .B2(new_n1021), .ZN(G387));
  INV_X1    g0822(.A(new_n1017), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n764), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1017), .A2(new_n763), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1024), .A2(new_n720), .A3(new_n1025), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n711), .A2(new_n829), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n210), .A2(new_n329), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n1028), .A2(new_n722), .B1(G107), .B2(new_n210), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n235), .A2(new_n277), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n722), .B(new_n277), .C1(new_n244), .C2(new_n297), .ZN(new_n1031));
  XOR2_X1   g0831(.A(KEYINPUT107), .B(KEYINPUT50), .Z(new_n1032));
  NOR3_X1   g0832(.A1(new_n1032), .A2(G50), .A3(new_n343), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1032), .B1(G50), .B2(new_n343), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n943), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1029), .B1(new_n1030), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n785), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n770), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n842), .A2(new_n949), .B1(new_n488), .B2(new_n812), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT108), .Z(new_n1041));
  XOR2_X1   g0841(.A(KEYINPUT109), .B(G322), .Z(new_n1042));
  OAI22_X1  g0842(.A1(new_n845), .A2(new_n1042), .B1(new_n811), .B2(new_n860), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT110), .ZN(new_n1044));
  AOI21_X1  g0844(.A(KEYINPUT48), .B1(new_n1041), .B2(new_n1044), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n800), .A2(new_n816), .B1(new_n791), .B2(new_n534), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1041), .A2(KEYINPUT48), .A3(new_n1044), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1047), .A2(KEYINPUT49), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n329), .B1(new_n825), .B2(G326), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(new_n473), .C2(new_n789), .ZN(new_n1051));
  AOI21_X1  g0851(.A(KEYINPUT49), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n800), .A2(new_n384), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1054), .B1(new_n297), .B2(new_n791), .C1(new_n202), .C2(new_n842), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n812), .A2(new_n244), .B1(new_n806), .B2(new_n342), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n332), .B(new_n1056), .C1(new_n382), .C2(new_n821), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1057), .B1(new_n471), .B2(new_n789), .C1(new_n807), .C2(new_n845), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n1051), .A2(new_n1052), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1039), .B1(new_n1059), .B2(new_n784), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n1023), .A2(new_n999), .B1(new_n1027), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1026), .A2(new_n1061), .ZN(G393));
  AND2_X1   g0862(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n999), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G311), .A2(new_n797), .B1(new_n803), .B2(G317), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT111), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n1066), .A2(KEYINPUT52), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(KEYINPUT52), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n823), .A2(G294), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1069), .B1(new_n473), .B2(new_n800), .C1(new_n488), .C2(new_n811), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT112), .Z(new_n1071));
  OAI21_X1  g0871(.A(new_n332), .B1(new_n1042), .B2(new_n806), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n790), .B(new_n1072), .C1(G283), .C2(new_n819), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1067), .A2(new_n1068), .A3(new_n1071), .A4(new_n1073), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(G150), .A2(new_n803), .B1(new_n797), .B2(G159), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT51), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n329), .B1(new_n811), .B2(new_n202), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n812), .A2(new_n343), .B1(new_n806), .B2(new_n843), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n864), .B1(new_n244), .B2(new_n791), .C1(new_n297), .C2(new_n800), .ZN(new_n1079));
  OR4_X1    g0879(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n787), .B1(new_n1074), .B2(new_n1080), .ZN(new_n1081));
  OR2_X1    g0881(.A1(new_n943), .A2(new_n242), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1038), .B1(G97), .B2(new_n719), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n773), .B(new_n1081), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n974), .B2(new_n829), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1064), .A2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1017), .A2(new_n763), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1087), .A2(new_n1063), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT113), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n721), .B1(new_n1087), .B2(new_n1063), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1086), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(G390));
  OAI211_X1 g0892(.A(G330), .B(new_n924), .C1(new_n760), .C2(new_n761), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n885), .A2(new_n882), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n1094), .A2(new_n881), .B1(new_n873), .B2(new_n872), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n896), .B1(new_n1095), .B2(KEYINPUT38), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n833), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n400), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n701), .B(new_n1099), .C1(new_n726), .C2(new_n730), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n832), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n903), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n892), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1096), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(KEYINPUT38), .B1(new_n888), .B2(new_n889), .ZN(new_n1105));
  NOR3_X1   g0905(.A1(new_n890), .A2(new_n1105), .A3(new_n870), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(new_n1096), .B2(new_n870), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n679), .A2(new_n701), .A3(new_n835), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n905), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n892), .B1(new_n1109), .B2(new_n903), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1093), .B(new_n1104), .C1(new_n1107), .C2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n906), .B1(new_n736), .B2(new_n835), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n903), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1103), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n891), .A2(new_n897), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n918), .A2(new_n892), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1114), .A2(new_n1115), .B1(new_n1116), .B2(new_n1102), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n916), .B1(new_n921), .B2(new_n922), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n924), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1111), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n469), .A2(new_n1118), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1121), .B(new_n691), .C1(new_n913), .C2(new_n737), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  AOI211_X1 g0923(.A(KEYINPUT114), .B(new_n903), .C1(new_n1118), .C2(new_n835), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT114), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n759), .A2(new_n753), .ZN(new_n1126));
  OAI211_X1 g0926(.A(G330), .B(new_n835), .C1(new_n761), .C2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1125), .B1(new_n1127), .B2(new_n1113), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n1100), .A2(new_n832), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1093), .A2(new_n1129), .ZN(new_n1130));
  NOR3_X1   g0930(.A1(new_n1124), .A2(new_n1128), .A3(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1113), .B1(new_n762), .B2(new_n834), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1112), .B1(new_n1132), .B2(new_n1119), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1123), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n721), .B1(new_n1120), .B2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n1120), .B2(new_n1134), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1115), .A2(new_n781), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n811), .A2(new_n395), .B1(new_n812), .B2(new_n471), .ZN(new_n1138));
  AND2_X1   g0938(.A1(new_n1138), .A2(KEYINPUT116), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1138), .A2(KEYINPUT116), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n789), .A2(new_n244), .B1(new_n806), .B2(new_n534), .ZN(new_n1141));
  OR3_X1    g0941(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  OR3_X1    g0942(.A1(new_n792), .A2(KEYINPUT117), .A3(new_n329), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(G77), .A2(new_n801), .B1(new_n803), .B2(G283), .ZN(new_n1144));
  OAI21_X1  g0944(.A(KEYINPUT117), .B1(new_n792), .B2(new_n329), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n797), .A2(G116), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1143), .A2(new_n1144), .A3(new_n1145), .A4(new_n1146), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n803), .A2(G128), .B1(new_n854), .B2(G50), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n1148), .B1(new_n850), .B2(new_n842), .C1(new_n807), .C2(new_n800), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n821), .A2(G137), .B1(new_n825), .B2(G125), .ZN(new_n1150));
  OR3_X1    g0950(.A1(new_n791), .A2(KEYINPUT53), .A3(new_n342), .ZN(new_n1151));
  OAI21_X1  g0951(.A(KEYINPUT53), .B1(new_n791), .B2(new_n342), .ZN(new_n1152));
  XOR2_X1   g0952(.A(KEYINPUT54), .B(G143), .Z(new_n1153));
  AOI21_X1  g0953(.A(new_n332), .B1(new_n823), .B2(new_n1153), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .A4(new_n1154), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n1142), .A2(new_n1147), .B1(new_n1149), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT118), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n787), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n1157), .B2(new_n1156), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n839), .A2(new_n343), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1137), .A2(new_n770), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  AND2_X1   g0961(.A1(new_n1136), .A2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1120), .A2(new_n998), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT115), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1162), .A2(new_n1164), .ZN(G378));
  INV_X1    g0965(.A(KEYINPUT123), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n903), .B1(new_n904), .B2(new_n906), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1167), .A2(new_n1103), .B1(new_n891), .B2(new_n897), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1093), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1113), .B1(new_n832), .B2(new_n1100), .ZN(new_n1170));
  NOR3_X1   g0970(.A1(new_n1170), .A2(new_n918), .A3(new_n892), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n1168), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1119), .B1(new_n1173), .B2(new_n1104), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1132), .A2(new_n1119), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n1109), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1127), .A2(new_n1113), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(KEYINPUT114), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1127), .A2(new_n1125), .A3(new_n1113), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1179), .A2(new_n1093), .A3(new_n1129), .A4(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1177), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1122), .B1(new_n1175), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n879), .A2(new_n353), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n689), .B2(new_n358), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n379), .A2(KEYINPUT10), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n373), .A2(new_n374), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n357), .B(new_n1184), .C1(new_n1187), .C2(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1192));
  AND3_X1   g0992(.A1(new_n1186), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1192), .B1(new_n1186), .B2(new_n1191), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(KEYINPUT122), .B1(new_n1195), .B2(KEYINPUT121), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1194), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1186), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1198), .A2(KEYINPUT122), .A3(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(G330), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1197), .B1(new_n930), .B2(new_n1202), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1196), .B(new_n1201), .C1(new_n926), .C2(new_n929), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n912), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n923), .B(new_n924), .C1(new_n887), .C2(new_n890), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n1206), .A2(KEYINPUT40), .B1(new_n927), .B2(new_n928), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1196), .B1(new_n1207), .B2(new_n1201), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT40), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n1096), .B2(new_n927), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n928), .A2(new_n923), .A3(new_n924), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1197), .B(new_n1202), .C1(new_n1210), .C2(new_n1211), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n898), .A2(new_n911), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1208), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1205), .A2(KEYINPUT57), .A3(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1166), .B1(new_n1183), .B2(new_n1215), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1208), .A2(new_n1213), .A3(new_n1212), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1213), .B1(new_n1208), .B2(new_n1212), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1123), .B1(new_n1120), .B2(new_n1134), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1219), .A2(KEYINPUT123), .A3(KEYINPUT57), .A4(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1216), .A2(new_n1221), .A3(new_n720), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(KEYINPUT124), .ZN(new_n1223));
  AOI211_X1 g1023(.A(KEYINPUT125), .B(KEYINPUT57), .C1(new_n1219), .C2(new_n1220), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT125), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1220), .A2(new_n1214), .A3(new_n1205), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT57), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1225), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1224), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT124), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1216), .A2(new_n1221), .A3(new_n1230), .A4(new_n720), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1223), .A2(new_n1229), .A3(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1195), .A2(new_n781), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(new_n332), .B2(new_n276), .ZN(new_n1235));
  AOI211_X1 g1035(.A(G41), .B(new_n329), .C1(new_n825), .C2(G283), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1236), .B1(new_n413), .B2(new_n789), .C1(new_n297), .C2(new_n791), .ZN(new_n1237));
  XOR2_X1   g1037(.A(new_n1237), .B(KEYINPUT119), .Z(new_n1238));
  OAI22_X1  g1038(.A1(new_n811), .A2(new_n471), .B1(new_n812), .B2(new_n384), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n842), .A2(new_n395), .B1(new_n845), .B2(new_n473), .ZN(new_n1240));
  NOR4_X1   g1040(.A1(new_n1238), .A2(new_n957), .A3(new_n1239), .A4(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1235), .B1(new_n1241), .B2(KEYINPUT58), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n811), .A2(new_n850), .B1(new_n812), .B2(new_n844), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(G150), .A2(new_n801), .B1(new_n803), .B2(G125), .ZN(new_n1244));
  INV_X1    g1044(.A(G128), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1244), .B1(new_n1245), .B2(new_n842), .ZN(new_n1246));
  AOI211_X1 g1046(.A(new_n1243), .B(new_n1246), .C1(new_n819), .C2(new_n1153), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT59), .ZN(new_n1248));
  OR2_X1    g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n854), .A2(G159), .ZN(new_n1251));
  AOI211_X1 g1051(.A(G33), .B(G41), .C1(new_n825), .C2(G124), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .A4(new_n1252), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1242), .B(new_n1253), .C1(KEYINPUT58), .C2(new_n1241), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n784), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n773), .B1(new_n202), .B2(new_n839), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1233), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  XOR2_X1   g1057(.A(new_n1257), .B(KEYINPUT120), .Z(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(new_n1219), .B2(new_n999), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1232), .A2(new_n1260), .ZN(G375));
  NAND2_X1  g1061(.A1(new_n1113), .A2(new_n781), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n845), .A2(new_n534), .B1(new_n791), .B2(new_n471), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(G283), .B2(new_n797), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n811), .A2(new_n473), .B1(new_n806), .B2(new_n857), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n329), .B(new_n1265), .C1(G107), .C2(new_n823), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1264), .A2(new_n962), .A3(new_n1054), .A4(new_n1266), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n842), .A2(new_n844), .B1(new_n202), .B2(new_n800), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1268), .B1(G159), .B2(new_n819), .ZN(new_n1269));
  OAI22_X1  g1069(.A1(new_n812), .A2(new_n342), .B1(new_n806), .B2(new_n1245), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n332), .B(new_n1270), .C1(new_n821), .C2(new_n1153), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n803), .A2(G132), .B1(new_n854), .B2(G58), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1269), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n787), .B1(new_n1267), .B2(new_n1273), .ZN(new_n1274));
  AOI211_X1 g1074(.A(new_n773), .B(new_n1274), .C1(new_n244), .C2(new_n839), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n1182), .A2(new_n999), .B1(new_n1262), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1134), .A2(new_n1020), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1182), .A2(new_n1123), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1276), .B1(new_n1277), .B2(new_n1278), .ZN(G381));
  OR2_X1    g1079(.A1(G393), .A2(G396), .ZN(new_n1280));
  OR3_X1    g1080(.A1(G390), .A2(G384), .A3(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(G378), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1232), .A2(new_n1282), .A3(new_n1260), .ZN(new_n1283));
  OR4_X1    g1083(.A1(G387), .A2(new_n1281), .A3(G381), .A4(new_n1283), .ZN(G407));
  OAI211_X1 g1084(.A(G407), .B(G213), .C1(G343), .C2(new_n1283), .ZN(G409));
  OAI21_X1  g1085(.A(KEYINPUT127), .B1(G387), .B2(new_n1091), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(G393), .B(G396), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(G387), .A2(new_n1091), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(G387), .A2(new_n1091), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1288), .B1(new_n1289), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1289), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1293), .A2(new_n1290), .A3(new_n1286), .A4(new_n1287), .ZN(new_n1294));
  AND2_X1   g1094(.A1(new_n1292), .A2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT61), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT60), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1297), .B1(new_n1182), .B2(new_n1123), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n721), .B1(new_n1298), .B2(new_n1278), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1299), .B1(new_n1278), .B2(new_n1298), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1276), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1301), .A2(new_n838), .A3(new_n867), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1300), .A2(G384), .A3(new_n1276), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n699), .A2(G213), .A3(G2897), .ZN(new_n1304));
  AND3_X1   g1104(.A1(new_n1302), .A2(new_n1303), .A3(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1304), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1282), .B1(new_n1232), .B2(new_n1260), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1219), .A2(new_n1020), .A3(new_n1220), .ZN(new_n1309));
  XNOR2_X1  g1109(.A(new_n1309), .B(KEYINPUT126), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1162), .A2(new_n1164), .A3(new_n1260), .ZN(new_n1311));
  OAI22_X1  g1111(.A1(new_n1310), .A2(new_n1311), .B1(new_n696), .B2(G343), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1307), .B1(new_n1308), .B2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1314));
  NOR3_X1   g1114(.A1(new_n1308), .A2(new_n1314), .A3(new_n1312), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT62), .ZN(new_n1316));
  OAI211_X1 g1116(.A(new_n1296), .B(new_n1313), .C1(new_n1315), .C2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(G375), .A2(G378), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1312), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1314), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1318), .A2(new_n1319), .A3(new_n1320), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1321), .A2(KEYINPUT62), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1295), .B1(new_n1317), .B2(new_n1322), .ZN(new_n1323));
  AND2_X1   g1123(.A1(new_n1313), .A2(new_n1296), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1292), .A2(new_n1294), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT63), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1321), .A2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1315), .A2(KEYINPUT63), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1324), .A2(new_n1325), .A3(new_n1327), .A4(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1323), .A2(new_n1329), .ZN(G405));
  INV_X1    g1130(.A(new_n1283), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1320), .B1(new_n1331), .B2(new_n1308), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1318), .A2(new_n1283), .A3(new_n1314), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  XNOR2_X1  g1134(.A(new_n1334), .B(new_n1325), .ZN(G402));
endmodule


