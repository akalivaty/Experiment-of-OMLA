//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 0 1 0 1 1 1 1 0 1 1 0 0 0 1 1 0 1 0 0 0 0 0 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1213, new_n1214, new_n1215, new_n1217, new_n1218, new_n1219,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  XNOR2_X1  g0013(.A(KEYINPUT66), .B(G68), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G58), .A2(G232), .ZN(new_n221));
  NAND4_X1  g0021(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n213), .B1(new_n217), .B2(new_n222), .ZN(new_n223));
  OR2_X1    g0023(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n213), .A2(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XOR2_X1   g0026(.A(KEYINPUT65), .B(KEYINPUT0), .Z(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n229));
  INV_X1    g0029(.A(new_n201), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n233), .A2(new_n211), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  AND4_X1   g0035(.A1(new_n224), .A2(new_n228), .A3(new_n229), .A4(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  INV_X1    g0037(.A(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n202), .A2(G68), .ZN(new_n249));
  INV_X1    g0049(.A(G68), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G50), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G58), .B(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n248), .B(new_n254), .ZN(G351));
  INV_X1    g0055(.A(G274), .ZN(new_n256));
  AND2_X1   g0056(.A1(G1), .A2(G13), .ZN(new_n257));
  NAND2_X1  g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n257), .A2(new_n258), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n260), .ZN(new_n264));
  INV_X1    g0064(.A(G226), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n262), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT3), .B(G33), .ZN(new_n267));
  INV_X1    g0067(.A(G1698), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(G222), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G77), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n267), .A2(G1698), .ZN(new_n271));
  INV_X1    g0071(.A(G223), .ZN(new_n272));
  OAI221_X1 g0072(.A(new_n269), .B1(new_n270), .B2(new_n267), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT67), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n257), .A2(new_n274), .A3(new_n258), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n274), .B1(new_n257), .B2(new_n258), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n266), .B1(new_n273), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G190), .ZN(new_n280));
  INV_X1    g0080(.A(G200), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n280), .B1(new_n281), .B2(new_n279), .ZN(new_n282));
  INV_X1    g0082(.A(G13), .ZN(new_n283));
  NOR3_X1   g0083(.A1(new_n283), .A2(new_n211), .A3(G1), .ZN(new_n284));
  NAND3_X1  g0084(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n233), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n210), .A2(G20), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n287), .A2(G50), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n284), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT8), .B(G58), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n211), .A2(G33), .ZN(new_n292));
  INV_X1    g0092(.A(G150), .ZN(new_n293));
  INV_X1    g0093(.A(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n211), .A2(new_n294), .ZN(new_n295));
  OAI22_X1  g0095(.A1(new_n291), .A2(new_n292), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n296), .B1(G20), .B2(new_n203), .ZN(new_n297));
  INV_X1    g0097(.A(new_n286), .ZN(new_n298));
  OAI221_X1 g0098(.A(new_n289), .B1(G50), .B2(new_n290), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT9), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(KEYINPUT68), .A2(KEYINPUT10), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n299), .A2(new_n300), .ZN(new_n304));
  NOR3_X1   g0104(.A1(new_n282), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(KEYINPUT68), .A2(KEYINPUT10), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n305), .B(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G179), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n279), .A2(new_n308), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n309), .B(new_n299), .C1(G169), .C2(new_n279), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n263), .A2(KEYINPUT67), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n275), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n294), .A2(KEYINPUT3), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT3), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G33), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n314), .A2(new_n316), .A3(G226), .A4(new_n268), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT69), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n267), .A2(KEYINPUT69), .A3(G226), .A4(new_n268), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n314), .A2(new_n316), .A3(G232), .A4(G1698), .ZN(new_n322));
  NAND2_X1  g0122(.A1(G33), .A2(G97), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n313), .B1(new_n321), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n262), .B1(new_n264), .B2(new_n216), .ZN(new_n327));
  OAI21_X1  g0127(.A(KEYINPUT13), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n327), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT13), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n324), .B1(new_n319), .B2(new_n320), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n329), .B(new_n330), .C1(new_n331), .C2(new_n313), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G169), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n335), .B1(new_n328), .B2(new_n332), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT14), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n334), .A2(G179), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT70), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n339), .B1(new_n336), .B2(new_n337), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NOR3_X1   g0141(.A1(new_n336), .A2(new_n339), .A3(new_n337), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n338), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n214), .A2(new_n211), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n295), .A2(new_n202), .B1(new_n292), .B2(new_n270), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n286), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT11), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(KEYINPUT12), .B1(new_n284), .B2(new_n250), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n283), .A2(G1), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n350), .A2(KEYINPUT12), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n349), .B1(new_n344), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n287), .A2(G68), .A3(new_n288), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n352), .B(new_n353), .C1(new_n347), .C2(new_n346), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n343), .B1(new_n348), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n333), .A2(G200), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n354), .A2(new_n348), .ZN(new_n357));
  INV_X1    g0157(.A(G190), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n356), .B(new_n357), .C1(new_n358), .C2(new_n333), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n291), .ZN(new_n361));
  NOR2_X1   g0161(.A1(G20), .A2(G33), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n361), .A2(new_n362), .B1(G20), .B2(G77), .ZN(new_n363));
  XOR2_X1   g0163(.A(KEYINPUT15), .B(G87), .Z(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n363), .B1(new_n292), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n286), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n287), .A2(G77), .A3(new_n288), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n367), .B(new_n368), .C1(G77), .C2(new_n290), .ZN(new_n369));
  INV_X1    g0169(.A(G244), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n262), .B1(new_n264), .B2(new_n370), .ZN(new_n371));
  OAI22_X1  g0171(.A1(new_n271), .A2(new_n216), .B1(new_n207), .B2(new_n267), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n314), .A2(new_n316), .ZN(new_n373));
  NOR3_X1   g0173(.A1(new_n373), .A2(new_n238), .A3(G1698), .ZN(new_n374));
  OR2_X1    g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n371), .B1(new_n375), .B2(new_n278), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n369), .B1(G190), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n281), .B2(new_n376), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n376), .A2(new_n308), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n379), .B(new_n369), .C1(G169), .C2(new_n376), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NOR3_X1   g0181(.A1(new_n311), .A2(new_n360), .A3(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n262), .B1(new_n264), .B2(new_n238), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n267), .A2(G223), .A3(new_n268), .ZN(new_n384));
  INV_X1    g0184(.A(G87), .ZN(new_n385));
  OAI221_X1 g0185(.A(new_n384), .B1(new_n294), .B2(new_n385), .C1(new_n271), .C2(new_n265), .ZN(new_n386));
  AOI211_X1 g0186(.A(new_n358), .B(new_n383), .C1(new_n386), .C2(new_n278), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n383), .B1(new_n386), .B2(new_n278), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n387), .B1(G200), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n287), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n361), .A2(new_n288), .ZN(new_n392));
  OAI22_X1  g0192(.A1(new_n391), .A2(new_n392), .B1(new_n290), .B2(new_n361), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT16), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT7), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n267), .B2(G20), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n373), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n215), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G159), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT71), .B1(new_n295), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT71), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n362), .A2(new_n402), .A3(G159), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n201), .B1(new_n214), .B2(G58), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n404), .B1(new_n405), .B2(new_n211), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n395), .B1(new_n399), .B2(new_n406), .ZN(new_n407));
  NOR3_X1   g0207(.A1(new_n267), .A2(new_n396), .A3(G20), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT7), .B1(new_n373), .B2(new_n211), .ZN(new_n409));
  OAI21_X1  g0209(.A(G68), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  AND2_X1   g0210(.A1(KEYINPUT66), .A2(G68), .ZN(new_n411));
  NOR2_X1   g0211(.A1(KEYINPUT66), .A2(G68), .ZN(new_n412));
  OAI21_X1  g0212(.A(G58), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n230), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n414), .A2(G20), .B1(new_n401), .B2(new_n403), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n410), .A2(KEYINPUT16), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n407), .A2(new_n416), .A3(new_n286), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT72), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n407), .A2(new_n416), .A3(KEYINPUT72), .A4(new_n286), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n390), .B(new_n394), .C1(new_n419), .C2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT17), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n422), .A2(KEYINPUT74), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n417), .A2(new_n418), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n393), .B1(new_n425), .B2(new_n420), .ZN(new_n426));
  OR2_X1    g0226(.A1(new_n423), .A2(KEYINPUT74), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n423), .A2(KEYINPUT74), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n426), .A2(new_n427), .A3(new_n390), .A4(new_n428), .ZN(new_n429));
  AND3_X1   g0229(.A1(new_n424), .A2(KEYINPUT75), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(KEYINPUT75), .B1(new_n424), .B2(new_n429), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n394), .B1(new_n419), .B2(new_n421), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT18), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n389), .A2(new_n308), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n388), .A2(new_n335), .ZN(new_n436));
  OR2_X1    g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n433), .A2(new_n434), .A3(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n435), .A2(new_n436), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT18), .B1(new_n426), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT73), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT73), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n438), .A2(new_n443), .A3(new_n440), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n432), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n382), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n287), .B1(G1), .B2(new_n294), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n448), .A2(new_n385), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n208), .A2(G87), .ZN(new_n450));
  INV_X1    g0250(.A(new_n323), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT80), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n452), .A2(KEYINPUT19), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT19), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(KEYINPUT80), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n451), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n450), .B1(new_n456), .B2(new_n211), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n454), .A2(KEYINPUT80), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n452), .A2(KEYINPUT19), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n458), .B(new_n459), .C1(new_n292), .C2(new_n206), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n314), .A2(new_n316), .A3(new_n211), .A4(G68), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(KEYINPUT81), .B1(new_n457), .B2(new_n462), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n460), .A2(new_n461), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n323), .B1(new_n458), .B2(new_n459), .ZN(new_n465));
  OAI22_X1  g0265(.A1(new_n465), .A2(G20), .B1(G87), .B2(new_n208), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT81), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n464), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n463), .A2(new_n286), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n365), .A2(new_n284), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT82), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT82), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n469), .A2(new_n473), .A3(new_n470), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n449), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(G45), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(G1), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n478), .A2(new_n263), .A3(G250), .ZN(new_n479));
  NOR2_X1   g0279(.A1(G238), .A2(G1698), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n480), .B1(new_n370), .B2(G1698), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n481), .A2(new_n267), .B1(G33), .B2(G116), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n479), .B1(new_n482), .B2(new_n313), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT78), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n259), .A2(new_n484), .A3(new_n477), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n484), .B1(new_n259), .B2(new_n477), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(KEYINPUT79), .B1(new_n483), .B2(new_n487), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n481), .A2(new_n267), .ZN(new_n489));
  INV_X1    g0289(.A(G116), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n294), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n278), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n263), .A2(G274), .ZN(new_n493));
  OAI21_X1  g0293(.A(KEYINPUT78), .B1(new_n493), .B2(new_n478), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n259), .A2(new_n484), .A3(new_n477), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT79), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n492), .A2(new_n496), .A3(new_n497), .A4(new_n479), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n488), .A2(new_n498), .A3(G190), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT83), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT83), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n488), .A2(new_n498), .A3(new_n501), .A4(G190), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n488), .A2(new_n498), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G200), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n475), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n469), .A2(new_n473), .A3(new_n470), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n473), .B1(new_n469), .B2(new_n470), .ZN(new_n508));
  OAI22_X1  g0308(.A1(new_n507), .A2(new_n508), .B1(new_n365), .B2(new_n448), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n504), .A2(new_n335), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n488), .A2(new_n498), .A3(new_n308), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n506), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n314), .A2(new_n316), .A3(G257), .A4(G1698), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n314), .A2(new_n316), .A3(G250), .A4(new_n268), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G33), .A2(G294), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  XNOR2_X1  g0317(.A(KEYINPUT5), .B(G41), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n518), .A2(new_n477), .B1(new_n257), .B2(new_n258), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n278), .A2(new_n517), .B1(new_n519), .B2(G264), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n259), .A2(new_n477), .A3(new_n518), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n335), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(G179), .B2(new_n522), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT86), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n314), .A2(new_n316), .A3(new_n211), .A4(G87), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(KEYINPUT84), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT84), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n267), .A2(new_n528), .A3(new_n211), .A4(G87), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT22), .ZN(new_n531));
  OAI21_X1  g0331(.A(KEYINPUT23), .B1(new_n211), .B2(G107), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT23), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n533), .A2(new_n207), .A3(G20), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n211), .A2(G33), .A3(G116), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT85), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n532), .A2(new_n534), .A3(new_n535), .A4(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n532), .A2(new_n534), .A3(new_n535), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT85), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n530), .A2(new_n531), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n527), .A2(new_n529), .A3(KEYINPUT22), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n525), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT24), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n298), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n530), .A2(new_n531), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n539), .A2(new_n537), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n541), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT86), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n540), .A2(new_n525), .A3(new_n541), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n548), .A2(KEYINPUT24), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n544), .A2(new_n550), .ZN(new_n551));
  AND2_X1   g0351(.A1(KEYINPUT87), .A2(KEYINPUT25), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n284), .A2(new_n207), .ZN(new_n553));
  NOR2_X1   g0353(.A1(KEYINPUT87), .A2(KEYINPUT25), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(new_n554), .B2(new_n553), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(new_n207), .B2(new_n448), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n524), .B1(new_n551), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n278), .A2(new_n517), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n519), .A2(G264), .ZN(new_n561));
  AND4_X1   g0361(.A1(new_n358), .A2(new_n560), .A3(new_n561), .A4(new_n521), .ZN(new_n562));
  AOI21_X1  g0362(.A(G200), .B1(new_n520), .B2(new_n521), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI211_X1 g0364(.A(new_n557), .B(new_n564), .C1(new_n544), .C2(new_n550), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n559), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n284), .A2(new_n490), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n287), .B(G116), .C1(G1), .C2(new_n294), .ZN(new_n568));
  NAND2_X1  g0368(.A1(G33), .A2(G283), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n569), .B(new_n211), .C1(G33), .C2(new_n206), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n570), .B(new_n286), .C1(new_n211), .C2(G116), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT20), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n571), .A2(new_n572), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n567), .B(new_n568), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n267), .A2(G257), .A3(new_n268), .ZN(new_n576));
  INV_X1    g0376(.A(G303), .ZN(new_n577));
  INV_X1    g0377(.A(G264), .ZN(new_n578));
  OAI221_X1 g0378(.A(new_n576), .B1(new_n577), .B2(new_n267), .C1(new_n271), .C2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n278), .ZN(new_n580));
  INV_X1    g0380(.A(new_n521), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(G270), .B2(new_n519), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n583), .A2(new_n358), .ZN(new_n584));
  AOI211_X1 g0384(.A(new_n575), .B(new_n584), .C1(G200), .C2(new_n583), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n583), .A2(G169), .A3(new_n575), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT21), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n575), .A2(G179), .A3(new_n580), .A4(new_n582), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n583), .A2(KEYINPUT21), .A3(G169), .A4(new_n575), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n585), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n314), .A2(new_n316), .A3(G244), .A4(new_n268), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT4), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n267), .A2(KEYINPUT4), .A3(G244), .A4(new_n268), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n595), .A2(new_n596), .A3(new_n569), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n314), .A2(new_n316), .A3(G250), .A4(G1698), .ZN(new_n598));
  XNOR2_X1  g0398(.A(new_n598), .B(KEYINPUT76), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n313), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT77), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n519), .A2(G257), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n521), .ZN(new_n603));
  NOR3_X1   g0403(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT76), .ZN(new_n605));
  XNOR2_X1  g0405(.A(new_n598), .B(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n595), .A2(new_n596), .A3(new_n569), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n278), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n603), .ZN(new_n609));
  AOI21_X1  g0409(.A(KEYINPUT77), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n335), .B1(new_n604), .B2(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n600), .A2(new_n603), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT6), .ZN(new_n613));
  NOR3_X1   g0413(.A1(new_n613), .A2(new_n206), .A3(G107), .ZN(new_n614));
  XNOR2_X1  g0414(.A(G97), .B(G107), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n614), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  OAI22_X1  g0416(.A1(new_n616), .A2(new_n211), .B1(new_n270), .B2(new_n295), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n207), .B1(new_n397), .B2(new_n398), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n286), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  MUX2_X1   g0419(.A(new_n290), .B(new_n448), .S(G97), .Z(new_n620));
  AOI22_X1  g0420(.A1(new_n612), .A2(new_n308), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n601), .B1(new_n600), .B2(new_n603), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n608), .A2(KEYINPUT77), .A3(new_n609), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n622), .A2(G190), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n281), .B1(new_n608), .B2(new_n609), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n620), .A2(new_n619), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n611), .A2(new_n621), .B1(new_n624), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n566), .A2(new_n592), .A3(new_n628), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n447), .A2(new_n513), .A3(new_n629), .ZN(new_n630));
  XOR2_X1   g0430(.A(new_n630), .B(KEYINPUT88), .Z(G372));
  NAND2_X1  g0431(.A1(new_n424), .A2(new_n429), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT75), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n424), .A2(KEYINPUT75), .A3(new_n429), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n359), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n355), .B1(new_n637), .B2(new_n380), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n307), .B1(new_n639), .B2(new_n441), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n310), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n604), .A2(new_n610), .A3(new_n358), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n625), .A2(new_n626), .ZN(new_n644));
  AOI21_X1  g0444(.A(G169), .B1(new_n622), .B2(new_n623), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n608), .A2(new_n609), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n626), .B1(new_n646), .B2(G179), .ZN(new_n647));
  OAI22_X1  g0447(.A1(new_n643), .A2(new_n644), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n648), .A2(new_n565), .ZN(new_n649));
  INV_X1    g0449(.A(new_n449), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n492), .A2(new_n496), .A3(new_n479), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(G200), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n650), .B(new_n652), .C1(new_n507), .C2(new_n508), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT89), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n472), .A2(new_n474), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n656), .A2(KEYINPUT89), .A3(new_n650), .A4(new_n652), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n655), .A2(new_n657), .A3(new_n503), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n651), .A2(new_n335), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n509), .A2(new_n511), .A3(new_n659), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n557), .B1(new_n544), .B2(new_n550), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n661), .B1(new_n662), .B2(new_n524), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n649), .A2(new_n658), .A3(new_n660), .A4(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n645), .A2(new_n647), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n658), .A2(new_n665), .A3(new_n666), .A4(new_n660), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n506), .A2(new_n512), .A3(new_n666), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(KEYINPUT26), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n664), .A2(new_n667), .A3(new_n660), .A4(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n642), .B1(new_n447), .B2(new_n671), .ZN(G369));
  NAND2_X1  g0472(.A1(new_n350), .A2(new_n211), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G213), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n575), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n591), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n592), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n680), .B1(new_n681), .B2(new_n679), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(G330), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n678), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n566), .B1(new_n662), .B2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n559), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n687), .B1(new_n688), .B2(new_n686), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT90), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n661), .A2(new_n678), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n566), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n559), .A2(new_n686), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n691), .A2(new_n695), .ZN(G399));
  INV_X1    g0496(.A(new_n225), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(G41), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n450), .A2(new_n490), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n698), .A2(new_n699), .A3(new_n210), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n700), .B1(new_n232), .B2(new_n698), .ZN(new_n701));
  XOR2_X1   g0501(.A(new_n701), .B(KEYINPUT28), .Z(new_n702));
  OR3_X1    g0502(.A1(new_n629), .A2(new_n513), .A3(new_n678), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT30), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n580), .A2(G179), .A3(new_n582), .A4(new_n520), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n504), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n622), .A2(new_n623), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n704), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n651), .A2(new_n308), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n709), .A2(new_n522), .A3(new_n583), .A4(new_n646), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n706), .A2(new_n707), .A3(new_n704), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n678), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT31), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n684), .B1(new_n703), .B2(new_n714), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n655), .A2(new_n657), .A3(new_n503), .ZN(new_n716));
  INV_X1    g0516(.A(new_n564), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n662), .A2(new_n717), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n718), .B(new_n628), .C1(new_n559), .C2(new_n591), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n660), .B1(new_n716), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n668), .A2(new_n665), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n658), .A2(KEYINPUT26), .A3(new_n666), .A4(new_n660), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(KEYINPUT91), .B1(new_n723), .B2(new_n678), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT91), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n722), .A2(new_n721), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n725), .B(new_n686), .C1(new_n726), .C2(new_n720), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(KEYINPUT29), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n670), .A2(new_n686), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT29), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n715), .B1(new_n729), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n702), .B1(new_n733), .B2(G1), .ZN(G364));
  INV_X1    g0534(.A(new_n685), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n683), .A2(new_n684), .ZN(new_n736));
  INV_X1    g0536(.A(new_n698), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n283), .A2(G20), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n210), .B1(new_n738), .B2(G45), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n735), .A2(new_n736), .A3(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n225), .A2(G355), .A3(new_n267), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n697), .A2(new_n267), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(G45), .B2(new_n231), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n254), .A2(new_n476), .ZN(new_n745));
  OAI221_X1 g0545(.A(new_n742), .B1(G116), .B2(new_n225), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G13), .A2(G33), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(G20), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n233), .B1(G20), .B2(new_n335), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n740), .B1(new_n746), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT92), .ZN(new_n753));
  INV_X1    g0553(.A(new_n750), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n211), .A2(G179), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G190), .A2(G200), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT95), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n755), .A2(new_n358), .A3(G200), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n758), .A2(G329), .B1(G283), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT96), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n211), .A2(new_n308), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(new_n756), .ZN(new_n764));
  INV_X1    g0564(.A(G311), .ZN(new_n765));
  INV_X1    g0565(.A(G322), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n763), .A2(G190), .A3(new_n281), .ZN(new_n767));
  OAI221_X1 g0567(.A(new_n373), .B1(new_n764), .B2(new_n765), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n763), .A2(G200), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G190), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  XOR2_X1   g0571(.A(KEYINPUT33), .B(G317), .Z(new_n772));
  NAND3_X1  g0572(.A1(new_n755), .A2(G190), .A3(G200), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n771), .A2(new_n772), .B1(new_n773), .B2(new_n577), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n769), .A2(new_n358), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G326), .ZN(new_n777));
  INV_X1    g0577(.A(G294), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n358), .A2(G179), .A3(G200), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n211), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n776), .A2(new_n777), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n768), .B(new_n774), .C1(KEYINPUT94), .C2(new_n781), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n762), .B(new_n782), .C1(KEYINPUT94), .C2(new_n781), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n776), .A2(new_n202), .B1(new_n759), .B2(new_n207), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n771), .A2(new_n250), .B1(new_n206), .B2(new_n780), .ZN(new_n785));
  INV_X1    g0585(.A(G58), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n267), .B1(new_n764), .B2(new_n270), .C1(new_n786), .C2(new_n767), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n784), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  XOR2_X1   g0588(.A(KEYINPUT93), .B(G159), .Z(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n757), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n773), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n792), .A2(KEYINPUT32), .B1(new_n793), .B2(G87), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n788), .B(new_n794), .C1(KEYINPUT32), .C2(new_n792), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n783), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n749), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n753), .B1(new_n754), .B2(new_n796), .C1(new_n682), .C2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n741), .A2(new_n798), .ZN(G396));
  NAND2_X1  g0599(.A1(new_n369), .A2(new_n678), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n378), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(new_n380), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n380), .A2(new_n678), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n748), .ZN(new_n806));
  INV_X1    g0606(.A(new_n740), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n750), .A2(new_n747), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n807), .B1(G77), .B2(new_n809), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n385), .A2(new_n759), .B1(new_n773), .B2(new_n207), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(G283), .B2(new_n770), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n758), .A2(G311), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n373), .B1(new_n764), .B2(new_n490), .ZN(new_n814));
  INV_X1    g0614(.A(new_n767), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n814), .B1(G294), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n780), .ZN(new_n817));
  AOI22_X1  g0617(.A1(G97), .A2(new_n817), .B1(new_n775), .B2(G303), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n812), .A2(new_n813), .A3(new_n816), .A4(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(KEYINPUT97), .B(G143), .ZN(new_n820));
  INV_X1    g0620(.A(new_n764), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n815), .A2(new_n820), .B1(new_n790), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n775), .A2(G137), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n822), .B(new_n823), .C1(new_n293), .C2(new_n771), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT34), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n202), .A2(new_n773), .B1(new_n759), .B2(new_n250), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n373), .B(new_n827), .C1(G58), .C2(new_n817), .ZN(new_n828));
  INV_X1    g0628(.A(G132), .ZN(new_n829));
  INV_X1    g0629(.A(new_n758), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n826), .B(new_n828), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n824), .A2(new_n825), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n819), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n810), .B1(new_n833), .B2(new_n750), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT98), .Z(new_n835));
  NOR2_X1   g0635(.A1(new_n806), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n670), .A2(new_n686), .A3(new_n805), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n838), .A2(KEYINPUT99), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n730), .A2(new_n804), .ZN(new_n840));
  XOR2_X1   g0640(.A(new_n839), .B(new_n840), .Z(new_n841));
  INV_X1    g0641(.A(new_n715), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n807), .B1(new_n841), .B2(new_n842), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n836), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(G384));
  NOR2_X1   g0647(.A1(new_n738), .A2(new_n210), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT104), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT37), .ZN(new_n850));
  INV_X1    g0650(.A(new_n676), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n433), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n850), .B1(new_n852), .B2(KEYINPUT103), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n433), .A2(new_n437), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n854), .A2(new_n852), .A3(new_n422), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n853), .B(new_n855), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n433), .B(new_n851), .C1(new_n632), .C2(new_n441), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT38), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n416), .A2(new_n286), .ZN(new_n861));
  AND2_X1   g0661(.A1(new_n410), .A2(new_n415), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n861), .B1(KEYINPUT16), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n394), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n851), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n432), .B2(new_n445), .ZN(new_n867));
  INV_X1    g0667(.A(new_n422), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n439), .A2(new_n676), .B1(new_n863), .B2(new_n394), .ZN(new_n869));
  OAI21_X1  g0669(.A(KEYINPUT37), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n852), .A2(new_n850), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n854), .A2(new_n422), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT38), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n867), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n860), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(KEYINPUT40), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n357), .A2(new_n686), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n333), .A2(G169), .ZN(new_n881));
  OAI22_X1  g0681(.A1(new_n881), .A2(KEYINPUT14), .B1(new_n308), .B2(new_n333), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n881), .A2(KEYINPUT70), .A3(KEYINPUT14), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n882), .B1(new_n340), .B2(new_n883), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n359), .B(new_n880), .C1(new_n884), .C2(new_n357), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT100), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n359), .B(new_n338), .C1(new_n341), .C2(new_n342), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n886), .B1(new_n887), .B2(new_n879), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n355), .A2(new_n886), .A3(new_n359), .A4(new_n880), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT101), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n703), .A2(new_n714), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT101), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n889), .A2(new_n890), .A3(new_n894), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n892), .A2(new_n893), .A3(new_n805), .A4(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n849), .B1(new_n878), .B2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n896), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n898), .A2(KEYINPUT104), .A3(KEYINPUT40), .A4(new_n877), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n438), .A2(new_n443), .A3(new_n440), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n443), .B1(new_n438), .B2(new_n440), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n865), .B1(new_n636), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n873), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n859), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NOR3_X1   g0705(.A1(new_n903), .A2(KEYINPUT102), .A3(new_n874), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT102), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n867), .B2(new_n875), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n905), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n898), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT40), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n897), .A2(new_n899), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(G330), .ZN(new_n913));
  INV_X1    g0713(.A(new_n447), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n715), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT105), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n912), .A2(new_n914), .A3(new_n893), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT106), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n859), .A2(new_n858), .B1(new_n867), .B2(new_n875), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT39), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT102), .B1(new_n903), .B2(new_n874), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n867), .A2(new_n907), .A3(new_n875), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n867), .A2(new_n873), .ZN(new_n927));
  AOI22_X1  g0727(.A1(new_n925), .A2(new_n926), .B1(new_n927), .B2(new_n859), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n924), .B1(new_n928), .B2(new_n923), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n355), .A2(new_n678), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n441), .A2(new_n676), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n837), .A2(new_n803), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n892), .A2(new_n895), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n932), .B1(new_n935), .B2(new_n928), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n931), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n729), .A2(new_n914), .A3(new_n732), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n938), .A2(new_n642), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n937), .B(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n848), .B1(new_n921), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n921), .B2(new_n940), .ZN(new_n942));
  INV_X1    g0742(.A(new_n616), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n943), .A2(KEYINPUT35), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(KEYINPUT35), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n944), .A2(G116), .A3(new_n234), .A4(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT36), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n232), .A2(G77), .A3(new_n413), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n249), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n949), .A2(G1), .A3(new_n283), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n942), .A2(new_n947), .A3(new_n950), .ZN(G367));
  INV_X1    g0751(.A(new_n743), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n751), .B1(new_n225), .B2(new_n365), .C1(new_n952), .C2(new_n244), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n953), .A2(new_n807), .ZN(new_n954));
  INV_X1    g0754(.A(G283), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n767), .A2(new_n577), .B1(new_n764), .B2(new_n955), .ZN(new_n956));
  AOI211_X1 g0756(.A(new_n267), .B(new_n956), .C1(G317), .C2(new_n791), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n775), .A2(G311), .B1(new_n760), .B2(G97), .ZN(new_n958));
  AOI22_X1  g0758(.A1(G107), .A2(new_n817), .B1(new_n770), .B2(G294), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT46), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n773), .B2(new_n490), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n957), .A2(new_n958), .A3(new_n959), .A4(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n793), .A2(KEYINPUT46), .A3(G116), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT110), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n770), .A2(new_n790), .B1(new_n821), .B2(G50), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT111), .Z(new_n966));
  OAI21_X1  g0766(.A(new_n267), .B1(new_n767), .B2(new_n293), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(G137), .B2(new_n791), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n780), .A2(new_n250), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(G77), .B2(new_n760), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n775), .A2(new_n820), .B1(new_n793), .B2(G58), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n968), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n962), .A2(new_n964), .B1(new_n966), .B2(new_n972), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n973), .B(KEYINPUT47), .Z(new_n974));
  OAI211_X1 g0774(.A(new_n658), .B(new_n660), .C1(new_n475), .C2(new_n686), .ZN(new_n975));
  OR3_X1    g0775(.A1(new_n660), .A2(new_n475), .A3(new_n686), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n954), .B1(new_n754), .B2(new_n974), .C1(new_n977), .C2(new_n797), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n739), .B(KEYINPUT109), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n666), .A2(new_n678), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n686), .B1(new_n619), .B2(new_n620), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n981), .B1(new_n648), .B2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT44), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n983), .B1(KEYINPUT107), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n695), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n984), .A2(KEYINPUT107), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n986), .B(new_n987), .Z(new_n988));
  NAND3_X1  g0788(.A1(new_n693), .A2(new_n694), .A3(new_n983), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT45), .Z(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n691), .B(new_n991), .Z(new_n992));
  OAI211_X1 g0792(.A(KEYINPUT108), .B(new_n693), .C1(new_n689), .C2(new_n692), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(KEYINPUT108), .B2(new_n693), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(new_n735), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n992), .A2(new_n733), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n733), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n698), .B(KEYINPUT41), .Z(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n980), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n691), .A2(new_n983), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n977), .A2(KEYINPUT43), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n688), .B1(new_n624), .B2(new_n627), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n686), .B1(new_n1003), .B2(new_n666), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n983), .A2(new_n566), .A3(new_n692), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(KEYINPUT42), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1005), .A2(KEYINPUT42), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1002), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n977), .A2(KEYINPUT43), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1001), .B(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n978), .B1(new_n1000), .B2(new_n1012), .ZN(G387));
  OR2_X1    g0813(.A1(new_n689), .A2(new_n797), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n225), .A2(new_n699), .A3(new_n267), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(G107), .B2(new_n225), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n241), .A2(new_n476), .ZN(new_n1017));
  AOI211_X1 g0817(.A(G45), .B(new_n699), .C1(G68), .C2(G77), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n291), .A2(G50), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT50), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n952), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1016), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n751), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n807), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n817), .A2(G283), .B1(new_n793), .B2(G294), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n815), .A2(G317), .B1(new_n821), .B2(G303), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n776), .B2(new_n766), .C1(new_n765), .C2(new_n771), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT48), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1025), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT114), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT115), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n1033), .A2(KEYINPUT49), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1033), .A2(KEYINPUT49), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n373), .B1(new_n757), .B2(new_n777), .C1(new_n490), .C2(new_n759), .ZN(new_n1036));
  NOR3_X1   g0836(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(KEYINPUT112), .B(G150), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n773), .A2(new_n270), .B1(new_n757), .B2(new_n1038), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT113), .Z(new_n1040));
  NOR2_X1   g0840(.A1(new_n365), .A2(new_n780), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n291), .B2(new_n771), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n267), .B1(new_n764), .B2(new_n250), .C1(new_n202), .C2(new_n767), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n776), .A2(new_n400), .B1(new_n759), .B2(new_n206), .ZN(new_n1045));
  NOR4_X1   g0845(.A1(new_n1040), .A2(new_n1043), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1037), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1024), .B1(new_n1047), .B2(new_n750), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n1014), .A2(new_n1048), .B1(new_n995), .B2(new_n980), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n733), .A2(new_n995), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(new_n698), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n733), .A2(new_n995), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1049), .B1(new_n1051), .B2(new_n1052), .ZN(G393));
  INV_X1    g0853(.A(new_n992), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n1050), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1055), .A2(new_n698), .A3(new_n996), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n751), .B1(new_n206), .B2(new_n225), .C1(new_n952), .C2(new_n248), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n807), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(G150), .A2(new_n775), .B1(new_n815), .B2(G159), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT51), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n780), .A2(new_n270), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(G50), .B2(new_n770), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n821), .A2(new_n361), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n373), .B1(new_n791), .B2(new_n820), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G87), .A2(new_n760), .B1(new_n793), .B2(new_n214), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1060), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1068), .A2(KEYINPUT116), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G317), .A2(new_n775), .B1(new_n815), .B2(G311), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT52), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n373), .B1(new_n757), .B2(new_n766), .C1(new_n778), .C2(new_n764), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n771), .A2(new_n577), .B1(new_n759), .B2(new_n207), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n780), .A2(new_n490), .B1(new_n773), .B2(new_n955), .ZN(new_n1074));
  OR4_X1    g0874(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1068), .A2(KEYINPUT116), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1069), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1058), .B1(new_n1077), .B2(new_n750), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n983), .B2(new_n797), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1056), .B(new_n1079), .C1(new_n1054), .C2(new_n979), .ZN(G390));
  NAND4_X1  g0880(.A1(new_n715), .A2(new_n805), .A3(new_n892), .A4(new_n895), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n930), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n933), .B2(new_n934), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1084), .B(new_n924), .C1(new_n923), .C2(new_n928), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT117), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n724), .A2(new_n727), .A3(new_n803), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n934), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1087), .A2(new_n1088), .A3(new_n802), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n922), .A2(new_n930), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  AND3_X1   g0891(.A1(new_n1085), .A2(new_n1086), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1086), .B1(new_n1085), .B2(new_n1091), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1082), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n1085), .A2(new_n1091), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1081), .B1(new_n1095), .B2(new_n1086), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n934), .B1(new_n842), .B2(new_n804), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n933), .B1(new_n1098), .B2(new_n1081), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1087), .A2(new_n802), .ZN(new_n1100));
  AND2_X1   g0900(.A1(new_n1098), .A2(new_n1081), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1099), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n938), .A2(new_n642), .A3(new_n915), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n737), .B1(new_n1097), .B2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1094), .A2(new_n1096), .A3(new_n1108), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n807), .B1(new_n361), .B2(new_n809), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1061), .B1(G283), .B2(new_n775), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n207), .B2(new_n771), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n830), .A2(new_n778), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n373), .B1(new_n764), .B2(new_n206), .C1(new_n490), .C2(new_n767), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n250), .A2(new_n759), .B1(new_n773), .B2(new_n385), .ZN(new_n1116));
  OR4_X1    g0916(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .A4(new_n1116), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(G128), .A2(new_n775), .B1(new_n815), .B2(G132), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1118), .B(KEYINPUT119), .ZN(new_n1119));
  OR3_X1    g0919(.A1(new_n773), .A2(new_n1038), .A3(KEYINPUT53), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n758), .A2(G125), .ZN(new_n1121));
  OAI21_X1  g0921(.A(KEYINPUT53), .B1(new_n773), .B2(new_n1038), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n267), .B1(new_n759), .B2(new_n202), .ZN(new_n1124));
  OR2_X1    g0924(.A1(new_n1124), .A2(KEYINPUT118), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(KEYINPUT118), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n770), .A2(G137), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(KEYINPUT54), .B(G143), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n817), .A2(G159), .B1(new_n821), .B2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .A4(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1117), .B1(new_n1123), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1111), .B1(new_n1132), .B2(new_n750), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n929), .B2(new_n748), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1134), .B1(new_n1097), .B2(new_n979), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1110), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(G378));
  NAND3_X1  g0937(.A1(new_n1109), .A2(KEYINPUT120), .A3(new_n1105), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n299), .A2(new_n851), .ZN(new_n1139));
  XOR2_X1   g0939(.A(new_n311), .B(new_n1139), .Z(new_n1140));
  XNOR2_X1  g0940(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1140), .B(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(new_n912), .B2(G330), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n912), .A2(G330), .A3(new_n1143), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1145), .A2(new_n937), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n937), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n912), .A2(G330), .A3(new_n1143), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1148), .B1(new_n1149), .B2(new_n1144), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1138), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(KEYINPUT120), .B1(new_n1109), .B2(new_n1105), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n737), .B1(new_n1154), .B2(KEYINPUT57), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT57), .ZN(new_n1156));
  OAI211_X1 g0956(.A(KEYINPUT121), .B(new_n1156), .C1(new_n1152), .C2(new_n1153), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1156), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT121), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1155), .A2(new_n1157), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1142), .A2(new_n747), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n809), .A2(G50), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n775), .A2(G125), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(new_n771), .B2(new_n829), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n815), .A2(G128), .B1(new_n821), .B2(G137), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n773), .B2(new_n1128), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1165), .B(new_n1167), .C1(G150), .C2(new_n817), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  OR2_X1    g0969(.A1(new_n1169), .A2(KEYINPUT59), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(KEYINPUT59), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n790), .A2(new_n760), .ZN(new_n1172));
  AOI211_X1 g0972(.A(G33), .B(G41), .C1(new_n791), .C2(G124), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .A4(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n267), .A2(G41), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1175), .B1(new_n767), .B2(new_n207), .C1(new_n365), .C2(new_n764), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n969), .B(new_n1176), .C1(G77), .C2(new_n793), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n955), .B2(new_n830), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n759), .A2(new_n786), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n206), .A2(new_n771), .B1(new_n776), .B2(new_n490), .ZN(new_n1180));
  NOR3_X1   g0980(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  OR2_X1    g0981(.A1(new_n1181), .A2(KEYINPUT58), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(KEYINPUT58), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1175), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1184), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1174), .A2(new_n1182), .A3(new_n1183), .A4(new_n1185), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n740), .B(new_n1163), .C1(new_n1186), .C2(new_n750), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n1151), .A2(new_n980), .B1(new_n1162), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1161), .A2(new_n1188), .ZN(G375));
  NAND2_X1  g0989(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1106), .A2(new_n999), .A3(new_n1190), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n1191), .B(KEYINPUT122), .Z(new_n1192));
  NAND2_X1  g0992(.A1(new_n934), .A2(new_n747), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n807), .B1(G68), .B2(new_n809), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n776), .A2(new_n829), .B1(new_n773), .B2(new_n400), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(new_n770), .B2(new_n1129), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n758), .A2(G128), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n267), .B1(new_n764), .B2(new_n293), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(G137), .B2(new_n815), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1179), .B1(G50), .B2(new_n817), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1196), .A2(new_n1197), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n776), .A2(new_n778), .B1(new_n773), .B2(new_n206), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G116), .B2(new_n770), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n758), .A2(G303), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n815), .A2(G283), .B1(new_n821), .B2(G107), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1203), .A2(new_n1042), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n373), .B1(new_n759), .B2(new_n270), .ZN(new_n1207));
  XOR2_X1   g1007(.A(new_n1207), .B(KEYINPUT123), .Z(new_n1208));
  OAI21_X1  g1008(.A(new_n1201), .B1(new_n1206), .B2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1194), .B1(new_n1209), .B2(new_n750), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1103), .A2(new_n980), .B1(new_n1193), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1192), .A2(new_n1211), .ZN(G381));
  NOR2_X1   g1012(.A1(G375), .A2(G378), .ZN(new_n1213));
  OR2_X1    g1013(.A1(G393), .A2(G396), .ZN(new_n1214));
  NOR4_X1   g1014(.A1(G387), .A2(G390), .A3(G384), .A4(new_n1214), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1213), .A2(new_n1211), .A3(new_n1192), .A4(new_n1215), .ZN(G407));
  NAND2_X1  g1016(.A1(new_n677), .A2(G213), .ZN(new_n1217));
  XOR2_X1   g1017(.A(new_n1217), .B(KEYINPUT124), .Z(new_n1218));
  NAND2_X1  g1018(.A1(new_n1213), .A2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(G407), .A2(G213), .A3(new_n1219), .ZN(G409));
  INV_X1    g1020(.A(KEYINPUT61), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1161), .A2(G378), .A3(new_n1188), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(new_n1152), .A2(new_n998), .A3(new_n1153), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1188), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1136), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1218), .B1(new_n1222), .B2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT60), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n1106), .B2(new_n1190), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1190), .A2(new_n1227), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(new_n698), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1211), .B1(new_n1228), .B2(new_n1230), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1231), .A2(new_n846), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n846), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1234), .A2(G2897), .A3(new_n1218), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT125), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(KEYINPUT125), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1217), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1240), .A2(G2897), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1235), .B1(new_n1239), .B2(new_n1241), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1221), .B1(new_n1226), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(KEYINPUT126), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1222), .A2(new_n1225), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1218), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1239), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1245), .A2(KEYINPUT62), .A3(new_n1246), .A4(new_n1247), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1240), .B(new_n1239), .C1(new_n1222), .C2(new_n1225), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1248), .B1(new_n1249), .B2(KEYINPUT62), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT126), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1251), .B(new_n1221), .C1(new_n1226), .C2(new_n1242), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1244), .A2(new_n1250), .A3(new_n1252), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(G387), .B(G390), .ZN(new_n1254));
  XOR2_X1   g1054(.A(G393), .B(G396), .Z(new_n1255));
  XNOR2_X1  g1055(.A(new_n1254), .B(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1253), .A2(new_n1256), .ZN(new_n1257));
  OR2_X1    g1057(.A1(new_n1249), .A2(KEYINPUT63), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1226), .A2(KEYINPUT63), .A3(new_n1247), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1240), .B1(new_n1222), .B2(new_n1225), .ZN(new_n1260));
  OR2_X1    g1060(.A1(new_n1260), .A2(new_n1242), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1256), .A2(KEYINPUT61), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1258), .A2(new_n1259), .A3(new_n1261), .A4(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1257), .A2(new_n1263), .ZN(G405));
  NAND2_X1  g1064(.A1(G375), .A2(new_n1136), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1265), .A2(new_n1222), .A3(new_n1234), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1222), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1247), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1266), .B(new_n1268), .C1(KEYINPUT127), .C2(new_n1256), .ZN(new_n1269));
  AND2_X1   g1069(.A1(new_n1256), .A2(KEYINPUT127), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(new_n1269), .B(new_n1270), .ZN(G402));
endmodule


