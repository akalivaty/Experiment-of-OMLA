//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 1 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0 0 1 1 0 1 0 0 1 0 1 0 0 1 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041;
  INV_X1    g000(.A(KEYINPUT86), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G116), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT66), .B(G116), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(new_n188), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT2), .B(G113), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n192), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n194), .B(new_n189), .C1(new_n188), .C2(new_n190), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT4), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n198));
  INV_X1    g012(.A(G107), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  AND2_X1   g014(.A1(KEYINPUT80), .A2(G104), .ZN(new_n201));
  NOR2_X1   g015(.A1(KEYINPUT80), .A2(G104), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n200), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n198), .A2(new_n199), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n198), .A2(new_n199), .A3(G104), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n203), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(KEYINPUT81), .A2(G101), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G101), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n203), .A2(new_n205), .A3(new_n211), .A4(new_n206), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n197), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  AOI21_X1  g027(.A(KEYINPUT4), .B1(new_n207), .B2(new_n209), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n196), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n199), .B1(new_n201), .B2(new_n202), .ZN(new_n216));
  NAND2_X1  g030(.A1(G104), .A2(G107), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(G101), .A3(new_n217), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n212), .A2(new_n218), .ZN(new_n219));
  OR2_X1    g033(.A1(new_n189), .A2(KEYINPUT5), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT5), .ZN(new_n221));
  OAI211_X1 g035(.A(G113), .B(new_n220), .C1(new_n191), .C2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n219), .A2(new_n195), .A3(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(G110), .B(G122), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n215), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n224), .B(KEYINPUT8), .ZN(new_n226));
  AND3_X1   g040(.A1(new_n219), .A2(new_n195), .A3(new_n222), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n222), .A2(new_n195), .B1(new_n212), .B2(new_n218), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G146), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G143), .ZN(new_n231));
  INV_X1    g045(.A(G143), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G146), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT64), .B(G128), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT1), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n236), .B1(G143), .B2(new_n230), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n234), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n231), .A2(new_n233), .A3(new_n236), .A4(G128), .ZN(new_n239));
  AOI21_X1  g053(.A(G125), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT0), .ZN(new_n242));
  INV_X1    g056(.A(G128), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(KEYINPUT0), .A2(G128), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n234), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n231), .B(new_n233), .C1(new_n242), .C2(new_n243), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G125), .ZN(new_n249));
  INV_X1    g063(.A(G224), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n250), .A2(G953), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n241), .A2(new_n249), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G125), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n254), .B1(new_n246), .B2(new_n247), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n251), .B1(new_n240), .B2(new_n255), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n253), .B(new_n256), .C1(KEYINPUT7), .C2(new_n251), .ZN(new_n257));
  OR4_X1    g071(.A1(KEYINPUT7), .A2(new_n240), .A3(new_n255), .A4(new_n251), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n225), .A2(new_n229), .A3(new_n257), .A4(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G902), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT85), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n224), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n193), .A2(new_n195), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT80), .B(G104), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n204), .B1(new_n266), .B2(new_n200), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n208), .B1(new_n267), .B2(new_n206), .ZN(new_n268));
  INV_X1    g082(.A(new_n212), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT4), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n214), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n265), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n264), .B1(new_n272), .B2(new_n227), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n273), .A2(KEYINPUT6), .A3(new_n225), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n253), .A2(new_n256), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n276), .B(new_n264), .C1(new_n272), .C2(new_n227), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n274), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n259), .A2(KEYINPUT85), .A3(new_n260), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n263), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(G210), .B1(G237), .B2(G902), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n187), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n278), .A2(new_n279), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT85), .B1(new_n259), .B2(new_n260), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n282), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n263), .A2(new_n281), .A3(new_n278), .A4(new_n279), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n283), .B1(new_n288), .B2(new_n187), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT93), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT89), .ZN(new_n291));
  INV_X1    g105(.A(G116), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT66), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT66), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G116), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n291), .B1(new_n296), .B2(G122), .ZN(new_n297));
  INV_X1    g111(.A(G122), .ZN(new_n298));
  AOI211_X1 g112(.A(KEYINPUT89), .B(new_n298), .C1(new_n293), .C2(new_n295), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT14), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT91), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n292), .A2(G122), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n300), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT14), .ZN(new_n305));
  OAI21_X1  g119(.A(KEYINPUT89), .B1(new_n190), .B2(new_n298), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n294), .A2(G116), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n292), .A2(KEYINPUT66), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n291), .B(G122), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n305), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(KEYINPUT91), .B1(new_n310), .B2(new_n302), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n306), .A2(new_n305), .A3(new_n309), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n304), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G107), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n306), .A2(new_n309), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(new_n199), .A3(new_n303), .ZN(new_n316));
  AND2_X1   g130(.A1(KEYINPUT64), .A2(G128), .ZN(new_n317));
  NOR2_X1   g131(.A1(KEYINPUT64), .A2(G128), .ZN(new_n318));
  OAI21_X1  g132(.A(G143), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n243), .A2(G143), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G134), .ZN(new_n323));
  INV_X1    g137(.A(G134), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n319), .A2(new_n324), .A3(new_n321), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n316), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n314), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT90), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n319), .A2(KEYINPUT13), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n330), .B1(new_n331), .B2(new_n321), .ZN(new_n332));
  AOI211_X1 g146(.A(KEYINPUT90), .B(new_n320), .C1(new_n319), .C2(KEYINPUT13), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n320), .A2(KEYINPUT13), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n324), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n199), .B1(new_n315), .B2(new_n303), .ZN(new_n337));
  AOI211_X1 g151(.A(G107), .B(new_n302), .C1(new_n306), .C2(new_n309), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n325), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  OR2_X1    g153(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  XOR2_X1   g154(.A(KEYINPUT9), .B(G234), .Z(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G217), .ZN(new_n343));
  NOR3_X1   g157(.A1(new_n342), .A2(new_n343), .A3(G953), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n329), .A2(new_n340), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n344), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n327), .B1(new_n313), .B2(G107), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n336), .A2(new_n339), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(G902), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(G478), .ZN(new_n351));
  NOR2_X1   g165(.A1(KEYINPUT92), .A2(KEYINPUT15), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(KEYINPUT92), .A2(KEYINPUT15), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n351), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n290), .B1(new_n350), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n344), .B1(new_n329), .B2(new_n340), .ZN(new_n358));
  NOR3_X1   g172(.A1(new_n347), .A2(new_n348), .A3(new_n346), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n260), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n360), .A2(KEYINPUT93), .A3(new_n355), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n260), .B(new_n356), .C1(new_n358), .C2(new_n359), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT94), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT94), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n350), .A2(new_n365), .A3(new_n356), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G953), .ZN(new_n368));
  NAND2_X1  g182(.A1(G234), .A2(G237), .ZN(new_n369));
  INV_X1    g183(.A(G952), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n370), .A2(KEYINPUT95), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n370), .A2(KEYINPUT95), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n368), .B(new_n369), .C1(new_n371), .C2(new_n372), .ZN(new_n373));
  XOR2_X1   g187(.A(KEYINPUT21), .B(G898), .Z(new_n374));
  NAND3_X1  g188(.A1(new_n369), .A2(G902), .A3(G953), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NOR2_X1   g190(.A1(G475), .A2(G902), .ZN(new_n377));
  XNOR2_X1  g191(.A(G125), .B(G140), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(KEYINPUT16), .ZN(new_n379));
  OR3_X1    g193(.A1(new_n254), .A2(KEYINPUT16), .A3(G140), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n379), .A2(G146), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(G146), .B1(new_n379), .B2(new_n380), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(G237), .A2(G953), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(G143), .A3(G214), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(G143), .B1(new_n384), .B2(G214), .ZN(new_n387));
  OAI211_X1 g201(.A(KEYINPUT17), .B(G131), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G237), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(new_n368), .A3(G214), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n232), .ZN(new_n391));
  INV_X1    g205(.A(G131), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n392), .A3(new_n385), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT87), .ZN(new_n394));
  OAI21_X1  g208(.A(G131), .B1(new_n386), .B2(new_n387), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT87), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n391), .A2(new_n396), .A3(new_n392), .A4(new_n385), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n394), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n383), .B(new_n388), .C1(new_n398), .C2(KEYINPUT17), .ZN(new_n399));
  XNOR2_X1  g213(.A(G113), .B(G122), .ZN(new_n400));
  XOR2_X1   g214(.A(new_n400), .B(G104), .Z(new_n401));
  XNOR2_X1  g215(.A(new_n378), .B(new_n230), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT18), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n391), .B(new_n385), .C1(new_n403), .C2(new_n392), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n402), .B(new_n404), .C1(new_n403), .C2(new_n395), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n399), .A2(new_n401), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n379), .A2(G146), .A3(new_n380), .ZN(new_n407));
  XOR2_X1   g221(.A(new_n378), .B(KEYINPUT19), .Z(new_n408));
  OAI211_X1 g222(.A(new_n398), .B(new_n407), .C1(G146), .C2(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n401), .B1(new_n409), .B2(new_n405), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n377), .B1(new_n406), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT20), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n409), .A2(new_n405), .ZN(new_n414));
  INV_X1    g228(.A(new_n401), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n399), .A2(new_n401), .A3(new_n405), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(KEYINPUT20), .A3(new_n377), .ZN(new_n419));
  AOI21_X1  g233(.A(KEYINPUT88), .B1(new_n416), .B2(new_n417), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n413), .A2(new_n419), .B1(new_n412), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n401), .B1(new_n399), .B2(new_n405), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n260), .B1(new_n406), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G475), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT88), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n418), .A2(new_n425), .A3(new_n412), .ZN(new_n426));
  INV_X1    g240(.A(new_n377), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n424), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n421), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n362), .A2(new_n367), .A3(new_n376), .A4(new_n429), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n289), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(G221), .B1(new_n342), .B2(G902), .ZN(new_n432));
  OAI21_X1  g246(.A(G214), .B1(G237), .B2(G902), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n248), .B1(new_n213), .B2(new_n214), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n234), .B1(new_n237), .B2(new_n243), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n239), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n219), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT10), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n238), .A2(new_n239), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n219), .A2(KEYINPUT10), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT11), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n443), .B1(new_n324), .B2(G137), .ZN(new_n444));
  INV_X1    g258(.A(G137), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n445), .A2(KEYINPUT11), .A3(G134), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n324), .A2(G137), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n444), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(G131), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n444), .A2(new_n446), .A3(new_n392), .A4(new_n447), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n451), .B(KEYINPUT82), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n435), .A2(new_n440), .A3(new_n442), .A4(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n368), .A2(G227), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n454), .B(KEYINPUT79), .ZN(new_n455));
  XNOR2_X1  g269(.A(G110), .B(G140), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n455), .B(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n435), .A2(new_n440), .A3(new_n442), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n459), .B1(new_n451), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(KEYINPUT83), .B1(new_n219), .B2(new_n441), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n212), .A2(new_n218), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n231), .A2(new_n233), .A3(G128), .ZN(new_n464));
  OAI21_X1  g278(.A(KEYINPUT1), .B1(new_n232), .B2(G146), .ZN(new_n465));
  OR2_X1    g279(.A1(KEYINPUT64), .A2(G128), .ZN(new_n466));
  NAND2_X1  g280(.A1(KEYINPUT64), .A2(G128), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  AOI22_X1  g282(.A1(new_n236), .A2(new_n464), .B1(new_n468), .B2(new_n234), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT83), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n463), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n462), .A2(new_n438), .A3(new_n471), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n472), .A2(KEYINPUT12), .A3(new_n451), .ZN(new_n473));
  AOI21_X1  g287(.A(KEYINPUT12), .B1(new_n472), .B2(new_n451), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n453), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT84), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI211_X1 g291(.A(KEYINPUT84), .B(new_n453), .C1(new_n473), .C2(new_n474), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n461), .B1(new_n479), .B2(new_n457), .ZN(new_n480));
  OAI21_X1  g294(.A(G469), .B1(new_n480), .B2(G902), .ZN(new_n481));
  INV_X1    g295(.A(G469), .ZN(new_n482));
  INV_X1    g296(.A(new_n473), .ZN(new_n483));
  INV_X1    g297(.A(new_n474), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n459), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n460), .A2(new_n451), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n458), .B1(new_n486), .B2(new_n453), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n482), .B(new_n260), .C1(new_n485), .C2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n434), .B1(new_n481), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n235), .A2(KEYINPUT23), .A3(G119), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n188), .A2(G128), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT23), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT74), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT74), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(KEYINPUT23), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n491), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(KEYINPUT75), .B1(new_n188), .B2(G128), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT75), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(new_n243), .A3(G119), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n490), .B1(new_n496), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT76), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n490), .B(KEYINPUT76), .C1(new_n496), .C2(new_n500), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n503), .A2(G110), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n188), .B1(new_n466), .B2(new_n467), .ZN(new_n506));
  INV_X1    g320(.A(new_n491), .ZN(new_n507));
  XNOR2_X1  g321(.A(KEYINPUT24), .B(G110), .ZN(new_n508));
  NOR3_X1   g322(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n382), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n509), .B1(new_n510), .B2(new_n407), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n505), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n508), .B1(new_n506), .B2(new_n507), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n513), .B1(new_n501), .B2(G110), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n378), .A2(new_n230), .ZN(new_n515));
  AND2_X1   g329(.A1(new_n407), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n368), .A2(G221), .A3(G234), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT77), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n518), .B(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(KEYINPUT22), .B(G137), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n518), .B(KEYINPUT77), .ZN(new_n523));
  INV_X1    g337(.A(new_n521), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n512), .A2(new_n517), .A3(new_n527), .ZN(new_n528));
  AOI22_X1  g342(.A1(new_n505), .A2(new_n511), .B1(new_n514), .B2(new_n516), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT78), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n522), .A2(new_n525), .A3(KEYINPUT78), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n528), .B(new_n260), .C1(new_n529), .C2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT25), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n512), .A2(new_n517), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n533), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n539), .A2(KEYINPUT25), .A3(new_n260), .A4(new_n528), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n343), .B1(G234), .B2(new_n260), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n542), .A2(G902), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n539), .A2(new_n528), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT28), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n451), .A2(new_n248), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n324), .A2(G137), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n445), .A2(G134), .ZN(new_n550));
  OAI21_X1  g364(.A(G131), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n450), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n441), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT70), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n548), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n265), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n554), .B1(new_n548), .B2(new_n553), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n547), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n548), .A2(new_n553), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n559), .A2(new_n196), .ZN(new_n560));
  AOI22_X1  g374(.A1(new_n548), .A2(new_n553), .B1(new_n193), .B2(new_n195), .ZN(new_n561));
  OAI21_X1  g375(.A(KEYINPUT28), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n384), .A2(G210), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT68), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT68), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n384), .A2(new_n565), .A3(G210), .ZN(new_n566));
  XNOR2_X1  g380(.A(KEYINPUT26), .B(G101), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n564), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  XOR2_X1   g382(.A(KEYINPUT26), .B(G101), .Z(new_n569));
  INV_X1    g383(.A(G210), .ZN(new_n570));
  NOR4_X1   g384(.A1(new_n570), .A2(KEYINPUT68), .A3(G237), .A4(G953), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n565), .B1(new_n384), .B2(G210), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n569), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n568), .A2(new_n573), .A3(new_n575), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT69), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(KEYINPUT69), .B1(new_n577), .B2(new_n578), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n558), .A2(new_n562), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT30), .ZN(new_n585));
  OR2_X1    g399(.A1(new_n585), .A2(KEYINPUT65), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(KEYINPUT65), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n450), .A2(new_n551), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n469), .A2(new_n588), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n449), .A2(new_n450), .B1(new_n246), .B2(new_n247), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n586), .B(new_n587), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n548), .A2(new_n553), .A3(KEYINPUT65), .A4(new_n585), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n265), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n579), .B1(new_n593), .B2(new_n560), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT29), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n584), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n558), .A2(KEYINPUT72), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n559), .A2(new_n196), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n265), .A2(new_n548), .A3(new_n553), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n598), .A2(KEYINPUT71), .A3(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT71), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n561), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n600), .A2(KEYINPUT28), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT72), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n604), .B(new_n547), .C1(new_n556), .C2(new_n557), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n579), .A2(new_n595), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n597), .A2(new_n603), .A3(new_n605), .A4(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n596), .A2(new_n607), .A3(new_n260), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(G472), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(KEYINPUT73), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT73), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n608), .A2(new_n611), .A3(G472), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n558), .A2(new_n562), .ZN(new_n614));
  INV_X1    g428(.A(new_n583), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n591), .A2(new_n592), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n560), .B1(new_n617), .B2(new_n196), .ZN(new_n618));
  INV_X1    g432(.A(new_n579), .ZN(new_n619));
  AOI21_X1  g433(.A(KEYINPUT31), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT31), .ZN(new_n621));
  NOR4_X1   g435(.A1(new_n593), .A2(new_n621), .A3(new_n560), .A4(new_n579), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n616), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(G472), .A2(G902), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n623), .A2(KEYINPUT32), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(KEYINPUT32), .B1(new_n623), .B2(new_n624), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n546), .B1(new_n613), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n431), .A2(new_n489), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G101), .ZN(G3));
  INV_X1    g444(.A(new_n429), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT97), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT33), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n633), .B1(new_n358), .B2(new_n359), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n345), .A2(KEYINPUT33), .A3(new_n349), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n634), .A2(new_n260), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(G478), .ZN(new_n637));
  AOI211_X1 g451(.A(G478), .B(G902), .C1(new_n345), .C2(new_n349), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n632), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  AOI211_X1 g454(.A(KEYINPUT97), .B(new_n638), .C1(new_n636), .C2(G478), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n631), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT98), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  OAI211_X1 g458(.A(KEYINPUT98), .B(new_n631), .C1(new_n640), .C2(new_n641), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n288), .A2(new_n433), .ZN(new_n647));
  INV_X1    g461(.A(new_n376), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n479), .A2(new_n457), .ZN(new_n650));
  INV_X1    g464(.A(new_n461), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n650), .A2(G469), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(G469), .A2(G902), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n652), .A2(new_n488), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n432), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n583), .B1(new_n558), .B2(new_n562), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n617), .A2(new_n196), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n657), .A2(new_n599), .A3(new_n619), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n621), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n618), .A2(KEYINPUT31), .A3(new_n619), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n656), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g475(.A(G472), .B1(new_n661), .B2(G902), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT96), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n623), .A2(new_n624), .ZN(new_n665));
  INV_X1    g479(.A(G472), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n666), .B1(new_n623), .B2(new_n260), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(KEYINPUT96), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n664), .A2(new_n665), .A3(new_n668), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n655), .A2(new_n546), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n646), .A2(new_n649), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT34), .B(G104), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G6));
  AND2_X1   g487(.A1(new_n362), .A2(new_n367), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n424), .A2(new_n413), .A3(new_n419), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n670), .A2(new_n649), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT35), .B(G107), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G9));
  AND3_X1   g493(.A1(new_n664), .A2(new_n665), .A3(new_n668), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT36), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n531), .A2(new_n681), .A3(new_n532), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n682), .A2(new_n529), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n682), .A2(new_n529), .ZN(new_n684));
  INV_X1    g498(.A(new_n544), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n686), .B1(new_n541), .B2(new_n542), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n431), .A2(new_n489), .A3(new_n680), .A4(new_n688), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT37), .B(G110), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G12));
  INV_X1    g505(.A(KEYINPUT32), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n665), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n623), .A2(KEYINPUT32), .A3(new_n624), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n608), .A2(new_n611), .A3(G472), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n611), .B1(new_n608), .B2(G472), .ZN(new_n696));
  OAI211_X1 g510(.A(new_n693), .B(new_n694), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n433), .ZN(new_n698));
  AOI211_X1 g512(.A(new_n698), .B(new_n687), .C1(new_n286), .C2(new_n287), .ZN(new_n699));
  AND4_X1   g513(.A1(new_n697), .A2(new_n699), .A3(new_n654), .A4(new_n432), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n373), .B(KEYINPUT101), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT99), .B(G900), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n703), .A2(new_n375), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  OR2_X1    g519(.A1(new_n705), .A2(KEYINPUT100), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(KEYINPUT100), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n702), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  AOI211_X1 g523(.A(new_n675), .B(new_n709), .C1(new_n362), .C2(new_n367), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n700), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G128), .ZN(G30));
  INV_X1    g526(.A(KEYINPUT38), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n289), .B(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NOR4_X1   g529(.A1(new_n715), .A2(new_n698), .A3(new_n674), .A4(new_n429), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n615), .A2(new_n602), .A3(new_n600), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(G472), .A3(new_n658), .ZN(new_n718));
  NAND2_X1  g532(.A1(G472), .A2(G902), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(KEYINPUT102), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT102), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n718), .A2(new_n722), .A3(new_n719), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n693), .A2(new_n721), .A3(new_n694), .A4(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n688), .ZN(new_n726));
  XOR2_X1   g540(.A(new_n708), .B(KEYINPUT39), .Z(new_n727));
  OR3_X1    g541(.A1(new_n655), .A2(KEYINPUT103), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g542(.A(KEYINPUT103), .B1(new_n655), .B2(new_n727), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n728), .A2(KEYINPUT40), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT40), .B1(new_n728), .B2(new_n729), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n716), .B(new_n726), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G143), .ZN(G45));
  OAI211_X1 g547(.A(new_n631), .B(new_n708), .C1(new_n640), .C2(new_n641), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n700), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G146), .ZN(G48));
  INV_X1    g551(.A(KEYINPUT104), .ZN(new_n738));
  INV_X1    g552(.A(new_n546), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n260), .B1(new_n485), .B2(new_n487), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(G469), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n741), .A2(new_n432), .A3(new_n488), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n697), .A2(new_n739), .A3(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n646), .A2(new_n738), .A3(new_n649), .A4(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n644), .A2(new_n649), .A3(new_n645), .A4(new_n744), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(KEYINPUT104), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(KEYINPUT41), .B(G113), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(G15));
  NOR2_X1   g564(.A1(new_n647), .A2(new_n742), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n676), .A2(new_n697), .A3(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n546), .A2(new_n648), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(new_n292), .ZN(G18));
  AND2_X1   g570(.A1(new_n699), .A2(new_n697), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n430), .A2(new_n742), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G119), .ZN(G21));
  INV_X1    g574(.A(new_n624), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n659), .A2(new_n660), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n597), .A2(new_n603), .A3(new_n605), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n615), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n761), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n667), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n743), .A2(new_n753), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n362), .A2(new_n367), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n768), .A2(new_n433), .A3(new_n631), .A4(new_n288), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(KEYINPUT105), .B(G122), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n770), .B(new_n771), .ZN(G24));
  NAND3_X1  g586(.A1(new_n743), .A2(new_n433), .A3(new_n288), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n766), .A2(new_n688), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n734), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(new_n254), .ZN(G27));
  AND3_X1   g590(.A1(new_n489), .A2(new_n628), .A3(new_n289), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n734), .A2(KEYINPUT42), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT106), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n780), .B(new_n692), .C1(new_n661), .C2(new_n761), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n694), .B(new_n781), .C1(new_n695), .C2(new_n696), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n626), .A2(new_n780), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n739), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n434), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n654), .A2(new_n289), .A3(new_n785), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n734), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT42), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n779), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(new_n392), .ZN(G33));
  NAND4_X1  g604(.A1(new_n489), .A2(new_n628), .A3(new_n289), .A4(new_n710), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT107), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G134), .ZN(G36));
  NAND2_X1  g607(.A1(new_n480), .A2(KEYINPUT45), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT45), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n458), .B1(new_n477), .B2(new_n478), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n795), .B1(new_n796), .B2(new_n461), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n794), .A2(G469), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n798), .A2(KEYINPUT46), .A3(new_n653), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n488), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT46), .B1(new_n798), .B2(new_n653), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n432), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n802), .A2(new_n727), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(KEYINPUT108), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n429), .B1(new_n640), .B2(new_n641), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT109), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT43), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n805), .A2(new_n806), .A3(KEYINPUT43), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n669), .A3(new_n688), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT44), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n289), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(new_n698), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(KEYINPUT110), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n811), .A2(KEYINPUT44), .A3(new_n669), .A4(new_n688), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n814), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n804), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(new_n445), .ZN(G39));
  XNOR2_X1  g635(.A(new_n802), .B(KEYINPUT47), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n816), .A2(new_n613), .A3(new_n627), .A4(new_n546), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n822), .A2(new_n734), .A3(new_n823), .ZN(new_n824));
  XOR2_X1   g638(.A(new_n824), .B(G140), .Z(G42));
  NOR3_X1   g639(.A1(new_n815), .A2(new_n698), .A3(new_n742), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n724), .A2(new_n373), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n826), .A2(new_n739), .A3(new_n827), .ZN(new_n828));
  NOR4_X1   g642(.A1(new_n828), .A2(new_n631), .A3(new_n640), .A4(new_n641), .ZN(new_n829));
  INV_X1    g643(.A(new_n766), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n830), .A2(new_n546), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n809), .A2(new_n701), .A3(new_n810), .A4(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(new_n433), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n833), .A2(new_n715), .A3(new_n743), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT50), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n833), .A2(KEYINPUT50), .A3(new_n715), .A4(new_n743), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n829), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n832), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT47), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n802), .B(new_n840), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n741), .A2(new_n488), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n843), .A2(new_n432), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n817), .B(new_n839), .C1(new_n841), .C2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n811), .A2(new_n701), .A3(new_n826), .ZN(new_n846));
  OR2_X1    g660(.A1(new_n846), .A2(new_n774), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n838), .A2(KEYINPUT51), .A3(new_n845), .A4(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n368), .B1(new_n371), .B2(new_n372), .ZN(new_n849));
  OR3_X1    g663(.A1(new_n846), .A2(KEYINPUT48), .A3(new_n784), .ZN(new_n850));
  OAI21_X1  g664(.A(KEYINPUT48), .B1(new_n846), .B2(new_n784), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT52), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n699), .A2(new_n654), .A3(new_n697), .A4(new_n432), .ZN(new_n855));
  INV_X1    g669(.A(new_n710), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n855), .B1(new_n856), .B2(new_n734), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n857), .A2(new_n775), .ZN(new_n858));
  INV_X1    g672(.A(new_n655), .ZN(new_n859));
  INV_X1    g673(.A(new_n769), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n859), .A2(new_n726), .A3(new_n860), .A4(new_n708), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n854), .B1(new_n858), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n700), .B1(new_n735), .B2(new_n710), .ZN(new_n863));
  OR3_X1    g677(.A1(new_n734), .A2(new_n773), .A3(new_n774), .ZN(new_n864));
  AND4_X1   g678(.A1(new_n854), .A2(new_n863), .A3(new_n864), .A4(new_n861), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n862), .A2(new_n865), .A3(KEYINPUT113), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT113), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n863), .A2(new_n864), .A3(new_n861), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(KEYINPUT52), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n858), .A2(new_n854), .A3(new_n861), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n867), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n866), .A2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n770), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n759), .B1(new_n754), .B2(new_n752), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n746), .A2(KEYINPUT104), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n746), .A2(KEYINPUT104), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n873), .B(new_n875), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n689), .A2(new_n629), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT86), .B1(new_n286), .B2(new_n287), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n376), .B1(new_n880), .B2(new_n283), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n768), .A2(new_n429), .ZN(new_n882));
  AOI211_X1 g696(.A(new_n698), .B(new_n881), .C1(new_n642), .C2(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n879), .B1(new_n670), .B2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(new_n782), .ZN(new_n885));
  INV_X1    g699(.A(new_n783), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n546), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n786), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n735), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  AOI22_X1  g703(.A1(new_n889), .A2(KEYINPUT42), .B1(new_n777), .B2(new_n778), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n697), .A2(new_n674), .ZN(new_n891));
  OAI22_X1  g705(.A1(new_n642), .A2(new_n830), .B1(new_n891), .B2(new_n675), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n892), .A2(new_n688), .A3(new_n708), .A4(new_n888), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n884), .A2(new_n890), .A3(new_n792), .A4(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n878), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT53), .B1(new_n872), .B2(new_n895), .ZN(new_n896));
  AOI211_X1 g710(.A(new_n770), .B(new_n874), .C1(new_n745), .C2(new_n747), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n881), .B1(new_n642), .B2(new_n882), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n670), .A2(new_n898), .A3(new_n433), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n893), .A2(new_n899), .A3(new_n629), .A4(new_n689), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT107), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n791), .B(new_n901), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n900), .A2(new_n789), .A3(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n862), .A2(new_n865), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n897), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT53), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT54), .B1(new_n896), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n905), .A2(new_n906), .ZN(new_n909));
  OAI21_X1  g723(.A(KEYINPUT113), .B1(new_n862), .B2(new_n865), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n869), .A2(new_n870), .A3(new_n867), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n895), .A2(KEYINPUT53), .A3(new_n910), .A4(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT54), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n909), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n908), .A2(KEYINPUT114), .A3(new_n914), .ZN(new_n915));
  OR2_X1    g729(.A1(new_n914), .A2(KEYINPUT114), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n853), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n839), .A2(new_n751), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n646), .A2(new_n739), .A3(new_n827), .A4(new_n826), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n822), .B1(new_n432), .B2(new_n843), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n920), .A2(KEYINPUT115), .A3(new_n817), .A4(new_n839), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT115), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n845), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n838), .A2(new_n921), .A3(new_n923), .A4(new_n847), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT51), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n924), .A2(KEYINPUT116), .A3(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(KEYINPUT116), .B1(new_n924), .B2(new_n925), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n917), .A2(new_n918), .A3(new_n919), .A4(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n370), .A2(new_n368), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n843), .A2(KEYINPUT49), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT112), .Z(new_n934));
  AOI211_X1 g748(.A(new_n805), .B(new_n934), .C1(KEYINPUT49), .C2(new_n843), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n546), .A2(new_n434), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT111), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n935), .A2(new_n725), .A3(new_n715), .A4(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n932), .A2(new_n938), .ZN(G75));
  INV_X1    g753(.A(KEYINPUT56), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n909), .A2(new_n912), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(G902), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n940), .B1(new_n942), .B2(new_n570), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n274), .A2(new_n277), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(new_n275), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT55), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n943), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n368), .A2(G952), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n940), .B(new_n946), .C1(new_n942), .C2(new_n570), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n948), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT117), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(G51));
  NOR2_X1   g768(.A1(new_n485), .A2(new_n487), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n914), .A2(KEYINPUT119), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n941), .A2(KEYINPUT54), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT119), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n909), .A2(new_n912), .A3(new_n958), .A4(new_n913), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n956), .A2(new_n957), .A3(new_n959), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n653), .B(KEYINPUT118), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT57), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n955), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n798), .B(KEYINPUT120), .Z(new_n964));
  NOR2_X1   g778(.A1(new_n942), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n950), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(KEYINPUT121), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT121), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n968), .B(new_n950), .C1(new_n963), .C2(new_n965), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n967), .A2(new_n969), .ZN(G54));
  NAND4_X1  g784(.A1(new_n941), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(new_n418), .Z(new_n972));
  NOR2_X1   g786(.A1(new_n972), .A2(new_n949), .ZN(G60));
  NAND2_X1  g787(.A1(G478), .A2(G902), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT59), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n915), .A2(new_n916), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n634), .A2(new_n635), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n949), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n960), .A2(new_n634), .A3(new_n635), .A4(new_n975), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n978), .A2(new_n979), .ZN(G63));
  XNOR2_X1  g794(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n981));
  NAND2_X1  g795(.A1(G217), .A2(G902), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT60), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n983), .B1(new_n909), .B2(new_n912), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n683), .A2(new_n684), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(new_n950), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n984), .B1(new_n539), .B2(new_n528), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n981), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OR2_X1    g803(.A1(new_n989), .A2(KEYINPUT123), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n987), .A2(new_n988), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(KEYINPUT61), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n989), .A2(KEYINPUT123), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n990), .A2(new_n992), .A3(new_n993), .ZN(G66));
  AOI21_X1  g808(.A(new_n368), .B1(new_n374), .B2(G224), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n897), .A2(new_n884), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n995), .B1(new_n996), .B2(new_n368), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(KEYINPUT124), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n944), .B1(G898), .B2(new_n368), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n998), .B(new_n999), .Z(G69));
  XOR2_X1   g814(.A(new_n617), .B(KEYINPUT125), .Z(new_n1001));
  XNOR2_X1  g815(.A(new_n1001), .B(new_n408), .ZN(new_n1002));
  INV_X1    g816(.A(G227), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n368), .B1(new_n1004), .B2(G900), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n642), .A2(new_n882), .ZN(new_n1006));
  OAI211_X1 g820(.A(new_n628), .B(new_n816), .C1(new_n1006), .C2(KEYINPUT126), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n728), .A2(new_n729), .ZN(new_n1008));
  AOI211_X1 g822(.A(new_n1007), .B(new_n1008), .C1(KEYINPUT126), .C2(new_n1006), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n820), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n732), .A2(new_n858), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT62), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n732), .A2(KEYINPUT62), .A3(new_n858), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n824), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g829(.A(G953), .B1(new_n1010), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1005), .B1(new_n1016), .B2(new_n1002), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n887), .A2(new_n860), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n819), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(new_n804), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n792), .A2(new_n858), .ZN(new_n1022));
  INV_X1    g836(.A(new_n1022), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n1021), .A2(new_n890), .A3(new_n1023), .ZN(new_n1024));
  NOR3_X1   g838(.A1(new_n1024), .A2(G953), .A3(new_n824), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1025), .B1(G227), .B2(G953), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1017), .B1(new_n1026), .B2(new_n1002), .ZN(G72));
  NAND2_X1  g841(.A1(new_n658), .A2(new_n594), .ZN(new_n1028));
  INV_X1    g842(.A(new_n1028), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n1010), .A2(new_n1015), .A3(new_n619), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n824), .A2(new_n619), .ZN(new_n1031));
  NAND4_X1  g845(.A1(new_n1021), .A2(new_n890), .A3(new_n1023), .A4(new_n1031), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n996), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g847(.A(new_n719), .B(KEYINPUT63), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1029), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g849(.A(new_n1034), .ZN(new_n1036));
  OAI211_X1 g850(.A(new_n1036), .B(new_n1028), .C1(new_n896), .C2(new_n907), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n1035), .A2(new_n950), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1038), .A2(KEYINPUT127), .ZN(new_n1039));
  INV_X1    g853(.A(KEYINPUT127), .ZN(new_n1040));
  NAND4_X1  g854(.A1(new_n1035), .A2(new_n1040), .A3(new_n950), .A4(new_n1037), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1039), .A2(new_n1041), .ZN(G57));
endmodule


