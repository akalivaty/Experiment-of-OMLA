//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 1 1 0 1 0 0 0 1 1 1 0 1 1 0 1 0 1 0 0 0 0 1 1 1 0 1 1 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 1 1 1 1 0 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(G137), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT11), .A3(G134), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n190), .A3(new_n192), .ZN(new_n193));
  OR2_X1    g007(.A1(new_n193), .A2(G131), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT66), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n195), .B1(new_n188), .B2(G137), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n191), .A2(KEYINPUT66), .A3(G134), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n190), .A3(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G131), .ZN(new_n199));
  AND3_X1   g013(.A1(new_n194), .A2(KEYINPUT71), .A3(new_n199), .ZN(new_n200));
  AOI21_X1  g014(.A(KEYINPUT71), .B1(new_n194), .B2(new_n199), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(G143), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT1), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(G128), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n204), .A2(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n202), .A2(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT67), .B(G128), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n207), .B1(G143), .B2(new_n204), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n208), .A2(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(KEYINPUT72), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT72), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n217), .B1(new_n208), .B2(new_n214), .ZN(new_n218));
  OAI22_X1  g032(.A1(new_n200), .A2(new_n201), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(G116), .B(G119), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT2), .B(G113), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n220), .B(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT0), .ZN(new_n225));
  INV_X1    g039(.A(G128), .ZN(new_n226));
  NOR3_X1   g040(.A1(new_n211), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(KEYINPUT0), .A2(G128), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n229), .B1(new_n209), .B2(new_n210), .ZN(new_n230));
  AND3_X1   g044(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n231));
  AOI21_X1  g045(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AND3_X1   g047(.A1(new_n230), .A2(KEYINPUT65), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(KEYINPUT65), .B1(new_n230), .B2(new_n233), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n228), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT65), .ZN(new_n239));
  INV_X1    g053(.A(new_n229), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n240), .B1(new_n203), .B2(new_n205), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT64), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n242), .B1(new_n225), .B2(new_n226), .ZN(new_n243));
  NAND3_X1  g057(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n239), .B1(new_n241), .B2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n230), .A2(new_n233), .A3(KEYINPUT65), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(KEYINPUT69), .A3(new_n228), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n238), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G131), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n193), .B(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(KEYINPUT70), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT70), .ZN(new_n255));
  AOI211_X1 g069(.A(new_n255), .B(new_n252), .C1(new_n238), .C2(new_n249), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n224), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT26), .B(G101), .ZN(new_n258));
  NOR2_X1   g072(.A1(G237), .A2(G953), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G210), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n258), .B(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT73), .B(KEYINPUT27), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n261), .B(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT68), .ZN(new_n264));
  INV_X1    g078(.A(new_n215), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n194), .A2(new_n199), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n215), .A2(KEYINPUT68), .A3(new_n194), .A4(new_n199), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n267), .B(new_n268), .C1(new_n252), .C2(new_n236), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n269), .A2(KEYINPUT30), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n219), .B1(new_n254), .B2(new_n256), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n270), .B1(new_n271), .B2(KEYINPUT30), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n257), .B(new_n263), .C1(new_n272), .C2(new_n222), .ZN(new_n273));
  INV_X1    g087(.A(new_n263), .ZN(new_n274));
  XOR2_X1   g088(.A(KEYINPUT75), .B(KEYINPUT28), .Z(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n222), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n269), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n276), .B1(new_n257), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n252), .B1(new_n238), .B2(new_n249), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n223), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n281), .A2(KEYINPUT28), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n274), .B1(new_n279), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n273), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT29), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT76), .ZN(new_n287));
  INV_X1    g101(.A(new_n219), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT69), .B1(new_n248), .B2(new_n228), .ZN(new_n289));
  AOI211_X1 g103(.A(new_n237), .B(new_n227), .C1(new_n246), .C2(new_n247), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n253), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n255), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n280), .A2(KEYINPUT70), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n288), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n257), .B1(new_n294), .B2(new_n222), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n282), .B1(new_n295), .B2(KEYINPUT28), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n263), .A2(new_n285), .ZN(new_n297));
  AOI21_X1  g111(.A(G902), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT76), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n284), .A2(new_n299), .A3(new_n285), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n287), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G472), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n223), .B1(new_n292), .B2(new_n293), .ZN(new_n303));
  INV_X1    g117(.A(new_n278), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n275), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n282), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n274), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n303), .A2(new_n263), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n308), .B1(new_n272), .B2(new_n222), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n307), .B1(KEYINPUT31), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT74), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n257), .A2(new_n274), .ZN(new_n312));
  INV_X1    g126(.A(new_n270), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT30), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n313), .B1(new_n294), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n312), .B1(new_n315), .B2(new_n277), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT31), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n311), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n317), .B(new_n308), .C1(new_n272), .C2(new_n222), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n319), .A2(KEYINPUT74), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n310), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  NOR2_X1   g135(.A1(G472), .A2(G902), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(KEYINPUT32), .A3(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT32), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n263), .B1(new_n279), .B2(new_n282), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n325), .B1(new_n316), .B2(new_n317), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n315), .A2(new_n277), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n327), .A2(new_n311), .A3(new_n317), .A4(new_n308), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n319), .A2(KEYINPUT74), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n326), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n322), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n324), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n302), .A2(new_n323), .A3(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(G214), .B1(G237), .B2(G902), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G952), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n336), .A2(G953), .ZN(new_n337));
  NAND2_X1  g151(.A1(G234), .A2(G237), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(G902), .A3(G953), .ZN(new_n341));
  XOR2_X1   g155(.A(new_n341), .B(KEYINPUT98), .Z(new_n342));
  XNOR2_X1  g156(.A(KEYINPUT21), .B(G898), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n340), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  XOR2_X1   g158(.A(G110), .B(G122), .Z(new_n345));
  XOR2_X1   g159(.A(new_n345), .B(KEYINPUT8), .Z(new_n346));
  INV_X1    g160(.A(G101), .ZN(new_n347));
  INV_X1    g161(.A(G104), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT82), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT82), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G104), .ZN(new_n351));
  INV_X1    g165(.A(G107), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n349), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n348), .A2(G107), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n347), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT85), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n355), .B(new_n356), .ZN(new_n357));
  XNOR2_X1  g171(.A(KEYINPUT82), .B(G104), .ZN(new_n358));
  OAI21_X1  g172(.A(KEYINPUT83), .B1(new_n358), .B2(new_n352), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n349), .A2(new_n351), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT83), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(new_n361), .A3(G107), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n353), .A2(KEYINPUT3), .ZN(new_n364));
  OR3_X1    g178(.A1(new_n348), .A2(KEYINPUT3), .A3(G107), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n363), .A2(new_n347), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n220), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n367), .A2(new_n221), .ZN(new_n368));
  INV_X1    g182(.A(G116), .ZN(new_n369));
  NOR3_X1   g183(.A1(new_n369), .A2(KEYINPUT5), .A3(G119), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n370), .B1(new_n220), .B2(KEYINPUT5), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n368), .B1(G113), .B2(new_n371), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n357), .A2(new_n366), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n372), .B1(new_n357), .B2(new_n366), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n346), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n375), .B(KEYINPUT93), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n361), .B1(new_n360), .B2(G107), .ZN(new_n377));
  AOI211_X1 g191(.A(KEYINPUT83), .B(new_n352), .C1(new_n349), .C2(new_n351), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n364), .B(new_n365), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT4), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(G101), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n381), .A2(new_n277), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n379), .A2(G101), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(KEYINPUT4), .A3(new_n366), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n373), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n345), .ZN(new_n386));
  XNOR2_X1  g200(.A(KEYINPUT92), .B(G224), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n388), .A2(G953), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(KEYINPUT7), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n236), .A2(G125), .ZN(new_n392));
  INV_X1    g206(.A(G125), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n265), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  AOI22_X1  g209(.A1(new_n385), .A2(new_n386), .B1(new_n391), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT91), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n392), .B(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(new_n394), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n376), .B(new_n396), .C1(new_n391), .C2(new_n399), .ZN(new_n400));
  AND2_X1   g214(.A1(new_n382), .A2(new_n384), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n345), .B1(new_n401), .B2(new_n373), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n385), .A2(new_n386), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n403), .A3(KEYINPUT6), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n399), .A2(new_n389), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n398), .A2(new_n390), .A3(new_n394), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OR3_X1    g221(.A1(new_n385), .A2(KEYINPUT6), .A3(new_n386), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n404), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(G902), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n400), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(G210), .B1(G237), .B2(G902), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n400), .A2(new_n409), .A3(new_n410), .A4(new_n412), .ZN(new_n415));
  AOI211_X1 g229(.A(new_n335), .B(new_n344), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n212), .A2(G143), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n226), .A2(G143), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n417), .A2(new_n188), .A3(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(G116), .B(G122), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n421), .B(new_n352), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n418), .B1(new_n417), .B2(KEYINPUT13), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT13), .ZN(new_n424));
  OAI21_X1  g238(.A(KEYINPUT97), .B1(new_n419), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(G134), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  AOI211_X1 g240(.A(KEYINPUT97), .B(new_n418), .C1(new_n417), .C2(KEYINPUT13), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n420), .B(new_n422), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  OR2_X1    g242(.A1(new_n369), .A2(G122), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n352), .B1(new_n429), .B2(KEYINPUT14), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n430), .B(new_n421), .ZN(new_n431));
  INV_X1    g245(.A(new_n420), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n188), .B1(new_n417), .B2(new_n419), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n431), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  XOR2_X1   g248(.A(KEYINPUT9), .B(G234), .Z(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(KEYINPUT81), .ZN(new_n436));
  INV_X1    g250(.A(G217), .ZN(new_n437));
  NOR3_X1   g251(.A1(new_n436), .A2(new_n437), .A3(G953), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n428), .A2(new_n434), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n438), .B1(new_n428), .B2(new_n434), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n410), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G478), .ZN(new_n443));
  OR2_X1    g257(.A1(new_n443), .A2(KEYINPUT15), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n442), .B(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT95), .ZN(new_n446));
  INV_X1    g260(.A(G140), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(G125), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n393), .A2(G140), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(new_n449), .A3(KEYINPUT16), .ZN(new_n450));
  OR3_X1    g264(.A1(new_n393), .A2(KEYINPUT16), .A3(G140), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n450), .A2(G146), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(G146), .B1(new_n450), .B2(new_n451), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n446), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n450), .A2(new_n451), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n204), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n450), .A2(new_n451), .A3(G146), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(KEYINPUT95), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(G237), .ZN(new_n459));
  INV_X1    g273(.A(G953), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n460), .A3(G214), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n202), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n259), .A2(G143), .A3(G214), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n251), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT17), .ZN(new_n465));
  INV_X1    g279(.A(new_n463), .ZN(new_n466));
  AOI21_X1  g280(.A(G143), .B1(new_n259), .B2(G214), .ZN(new_n467));
  OAI21_X1  g281(.A(G131), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT17), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n462), .A2(new_n251), .A3(new_n463), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n454), .A2(new_n458), .A3(new_n465), .A4(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(G113), .B(G122), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(new_n348), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n464), .A2(KEYINPUT18), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n448), .A2(new_n449), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n476), .B(G146), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n462), .A2(new_n463), .ZN(new_n478));
  AND2_X1   g292(.A1(KEYINPUT18), .A2(G131), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n475), .B(new_n477), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n472), .A2(new_n474), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n474), .B1(new_n472), .B2(new_n480), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n410), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT96), .B(G475), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(G475), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n476), .A2(KEYINPUT19), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT19), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n448), .A2(new_n449), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n487), .A2(new_n204), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT94), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n468), .A2(new_n470), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n487), .A2(KEYINPUT94), .A3(new_n204), .A4(new_n489), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n492), .A2(new_n493), .A3(new_n457), .A4(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n474), .B1(new_n495), .B2(new_n480), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n486), .B(new_n410), .C1(new_n481), .C2(new_n496), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n497), .A2(KEYINPUT20), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT20), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n495), .A2(new_n480), .ZN(new_n500));
  INV_X1    g314(.A(new_n474), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n472), .A2(new_n474), .A3(new_n480), .ZN(new_n503));
  AOI21_X1  g317(.A(G475), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n499), .B1(new_n504), .B2(new_n410), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n485), .B1(new_n498), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n416), .A2(new_n445), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n212), .A2(G119), .ZN(new_n509));
  OR2_X1    g323(.A1(new_n509), .A2(KEYINPUT77), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(KEYINPUT77), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n510), .B(new_n511), .C1(G119), .C2(new_n226), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT24), .B(G110), .ZN(new_n513));
  OAI21_X1  g327(.A(KEYINPUT23), .B1(new_n226), .B2(G119), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT78), .ZN(new_n515));
  OR2_X1    g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n514), .A2(new_n515), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n226), .A2(G119), .ZN(new_n519));
  INV_X1    g333(.A(new_n509), .ZN(new_n520));
  AOI22_X1  g334(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(KEYINPUT23), .ZN(new_n521));
  INV_X1    g335(.A(G110), .ZN(new_n522));
  AOI22_X1  g336(.A1(new_n512), .A2(new_n513), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n457), .B1(G146), .B2(new_n476), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI22_X1  g339(.A1(new_n512), .A2(new_n513), .B1(new_n452), .B2(new_n453), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n521), .A2(new_n522), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n460), .A2(G221), .A3(G234), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n530), .B(KEYINPUT22), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n531), .B(G137), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n532), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n534), .B1(new_n525), .B2(new_n528), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n533), .A2(new_n410), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT79), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(KEYINPUT25), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n437), .B1(G234), .B2(new_n410), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n533), .A2(new_n535), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(KEYINPUT80), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n539), .A2(G902), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  OR2_X1    g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(G469), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n381), .B1(new_n289), .B2(new_n290), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n383), .A2(KEYINPUT4), .A3(new_n366), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT84), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT10), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n265), .A2(new_n217), .ZN(new_n553));
  INV_X1    g367(.A(new_n218), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n357), .A2(new_n366), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n211), .B1(new_n213), .B2(new_n226), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n208), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n357), .A2(new_n558), .A3(new_n366), .ZN(new_n559));
  AOI22_X1  g373(.A1(new_n555), .A2(new_n556), .B1(new_n559), .B2(new_n552), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT84), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n250), .A2(new_n384), .A3(new_n561), .A4(new_n381), .ZN(new_n562));
  XOR2_X1   g376(.A(new_n252), .B(KEYINPUT86), .Z(new_n563));
  NAND4_X1  g377(.A1(new_n551), .A2(new_n560), .A3(new_n562), .A4(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(G110), .B(G140), .ZN(new_n565));
  INV_X1    g379(.A(G227), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n566), .A2(G953), .ZN(new_n567));
  XOR2_X1   g381(.A(new_n565), .B(new_n567), .Z(new_n568));
  AND3_X1   g382(.A1(new_n564), .A2(KEYINPUT90), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n559), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n215), .B1(new_n357), .B2(new_n366), .ZN(new_n571));
  OAI211_X1 g385(.A(KEYINPUT12), .B(new_n253), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT87), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n559), .B1(new_n556), .B2(new_n215), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n575), .A2(KEYINPUT87), .A3(KEYINPUT12), .A4(new_n253), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n253), .B1(new_n570), .B2(new_n571), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT12), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n574), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(KEYINPUT90), .B1(new_n564), .B2(new_n568), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n569), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n551), .A2(new_n560), .A3(new_n562), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(KEYINPUT89), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT89), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n551), .A2(new_n586), .A3(new_n560), .A4(new_n562), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(new_n253), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n568), .B1(new_n588), .B2(new_n564), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n548), .B(new_n410), .C1(new_n583), .C2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n580), .A2(new_n564), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT88), .ZN(new_n592));
  INV_X1    g406(.A(new_n568), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT88), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n580), .A2(new_n594), .A3(new_n564), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n588), .A2(new_n564), .A3(new_n568), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(G469), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(G469), .A2(G902), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n590), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(G221), .B1(new_n436), .B2(G902), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n333), .A2(new_n508), .A3(new_n547), .A4(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT99), .B(G101), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G3));
  NAND2_X1  g420(.A1(new_n329), .A2(new_n328), .ZN(new_n607));
  AOI21_X1  g421(.A(G902), .B1(new_n607), .B2(new_n310), .ZN(new_n608));
  INV_X1    g422(.A(G472), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n331), .B1(new_n607), .B2(new_n310), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n601), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n546), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n612), .A2(new_n600), .A3(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n416), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT33), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n617), .B1(new_n440), .B2(new_n441), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n428), .A2(new_n434), .ZN(new_n619));
  INV_X1    g433(.A(new_n438), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n621), .A2(KEYINPUT33), .A3(new_n439), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n443), .A2(G902), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n618), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n442), .A2(new_n443), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n506), .A2(new_n626), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n615), .A2(new_n616), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(KEYINPUT34), .B(G104), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G6));
  AOI21_X1  g444(.A(new_n335), .B1(new_n414), .B2(new_n415), .ZN(new_n631));
  INV_X1    g445(.A(new_n344), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n445), .A2(new_n506), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT100), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n416), .A2(KEYINPUT100), .A3(new_n633), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n615), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT101), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT35), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G107), .ZN(G9));
  NOR2_X1   g455(.A1(new_n534), .A2(KEYINPUT36), .ZN(new_n642));
  XOR2_X1   g456(.A(new_n529), .B(new_n642), .Z(new_n643));
  AOI22_X1  g457(.A1(new_n538), .A2(new_n539), .B1(new_n543), .B2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n508), .A2(new_n612), .A3(new_n603), .A4(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT37), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(new_n522), .ZN(G12));
  INV_X1    g462(.A(G900), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n342), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(new_n339), .B(KEYINPUT102), .Z(new_n651));
  NOR2_X1   g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n633), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n602), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n333), .A2(new_n655), .A3(new_n631), .A4(new_n645), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G128), .ZN(G30));
  NAND2_X1  g471(.A1(new_n414), .A2(new_n415), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT38), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n507), .A2(new_n335), .A3(new_n445), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(new_n652), .B(KEYINPUT39), .Z(new_n662));
  NAND2_X1  g476(.A1(new_n603), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n661), .B1(new_n663), .B2(KEYINPUT40), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n303), .B1(new_n315), .B2(new_n277), .ZN(new_n665));
  OR2_X1    g479(.A1(new_n665), .A2(new_n263), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n410), .B1(new_n295), .B2(new_n274), .ZN(new_n668));
  OAI21_X1  g482(.A(G472), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n332), .A2(new_n323), .A3(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(new_n645), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n664), .B(new_n671), .C1(KEYINPUT40), .C2(new_n663), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G143), .ZN(G45));
  NAND4_X1  g487(.A1(new_n333), .A2(new_n603), .A3(new_n631), .A4(new_n645), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT103), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n497), .A2(KEYINPUT20), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n504), .A2(new_n499), .A3(new_n410), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AOI22_X1  g492(.A1(new_n678), .A2(new_n485), .B1(new_n624), .B2(new_n625), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n675), .B1(new_n679), .B2(new_n653), .ZN(new_n680));
  AND4_X1   g494(.A1(new_n675), .A2(new_n506), .A3(new_n626), .A4(new_n653), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n674), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(new_n204), .ZN(G48));
  NOR2_X1   g499(.A1(new_n616), .A2(new_n627), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n410), .B1(new_n583), .B2(new_n589), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(G469), .ZN(new_n688));
  AND3_X1   g502(.A1(new_n688), .A2(new_n601), .A3(new_n590), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n333), .A2(new_n686), .A3(new_n547), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(KEYINPUT41), .B(G113), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G15));
  NAND2_X1  g506(.A1(new_n636), .A2(new_n637), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n693), .A2(new_n333), .A3(new_n547), .A4(new_n689), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G116), .ZN(G18));
  NAND4_X1  g509(.A1(new_n333), .A2(new_n508), .A3(new_n645), .A4(new_n689), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G119), .ZN(G21));
  NOR2_X1   g511(.A1(new_n296), .A2(new_n274), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n698), .B1(new_n328), .B2(new_n329), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n309), .A2(KEYINPUT31), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n331), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT104), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n702), .B1(new_n608), .B2(new_n609), .ZN(new_n703));
  OAI211_X1 g517(.A(KEYINPUT104), .B(G472), .C1(new_n330), .C2(G902), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n701), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT105), .ZN(new_n706));
  AND3_X1   g520(.A1(new_n705), .A2(new_n706), .A3(new_n547), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n706), .B1(new_n705), .B2(new_n547), .ZN(new_n708));
  OR2_X1    g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n507), .A2(new_n445), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n709), .A2(new_n416), .A3(new_n710), .A4(new_n689), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G122), .ZN(G24));
  AND4_X1   g526(.A1(new_n601), .A2(new_n631), .A3(new_n688), .A4(new_n590), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT106), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n714), .B1(new_n680), .B2(new_n681), .ZN(new_n715));
  OAI21_X1  g529(.A(KEYINPUT103), .B1(new_n627), .B2(new_n652), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n679), .A2(new_n675), .A3(new_n653), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(KEYINPUT106), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n705), .A2(new_n645), .A3(new_n713), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G125), .ZN(G27));
  NOR4_X1   g535(.A1(new_n330), .A2(KEYINPUT107), .A3(new_n324), .A4(new_n331), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n723), .B1(new_n611), .B2(KEYINPUT32), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n611), .ZN(new_n726));
  AOI22_X1  g540(.A1(new_n301), .A2(G472), .B1(new_n726), .B2(new_n324), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n546), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n414), .A2(new_n334), .A3(new_n415), .ZN(new_n729));
  AND4_X1   g543(.A1(new_n601), .A2(new_n719), .A3(new_n600), .A4(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n728), .A2(KEYINPUT108), .A3(KEYINPUT42), .A4(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n323), .A2(KEYINPUT107), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n611), .A2(new_n723), .A3(KEYINPUT32), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n302), .A2(new_n732), .A3(new_n332), .A4(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n734), .A2(KEYINPUT42), .A3(new_n547), .A4(new_n730), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT108), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n600), .A2(new_n601), .A3(new_n729), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n333), .A2(new_n547), .A3(new_n719), .A4(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT42), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n731), .A2(new_n737), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G131), .ZN(G33));
  INV_X1    g557(.A(new_n654), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n333), .A2(new_n547), .A3(new_n744), .A4(new_n738), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G134), .ZN(G36));
  NAND2_X1  g560(.A1(new_n596), .A2(new_n597), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(KEYINPUT45), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(G469), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(KEYINPUT46), .A3(new_n599), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT46), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n753), .B(G469), .C1(new_n748), .C2(G902), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n749), .A2(KEYINPUT109), .A3(KEYINPUT46), .A4(new_n599), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n752), .A2(new_n590), .A3(new_n754), .A4(new_n755), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n756), .A2(new_n601), .A3(new_n662), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n729), .B(KEYINPUT111), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n759));
  AOI21_X1  g573(.A(KEYINPUT43), .B1(new_n507), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n507), .A2(new_n626), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n760), .B(new_n761), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n645), .B(new_n762), .C1(new_n610), .C2(new_n611), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT44), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n758), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n757), .B(new_n765), .C1(new_n764), .C2(new_n763), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G137), .ZN(G39));
  INV_X1    g581(.A(KEYINPUT47), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n756), .A2(new_n768), .A3(new_n601), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n768), .B1(new_n756), .B2(new_n601), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n333), .A2(new_n547), .A3(new_n683), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(new_n729), .A3(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G140), .ZN(G42));
  AND2_X1   g588(.A1(new_n688), .A2(new_n590), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT49), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n614), .A2(new_n334), .ZN(new_n778));
  AOI211_X1 g592(.A(new_n659), .B(new_n777), .C1(KEYINPUT112), .C2(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n778), .A2(KEYINPUT112), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(new_n761), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n775), .A2(new_n776), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n779), .A2(new_n781), .A3(new_n670), .A4(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT53), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n705), .A2(new_n645), .A3(new_n719), .A4(new_n738), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT114), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AOI211_X1 g602(.A(new_n644), .B(new_n701), .C1(new_n703), .C2(new_n704), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n789), .A2(KEYINPUT114), .A3(new_n719), .A4(new_n738), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n507), .A2(new_n445), .A3(new_n653), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n333), .A2(new_n645), .A3(new_n738), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n745), .A2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n633), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n796), .A2(KEYINPUT113), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(KEYINPUT113), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n797), .A2(new_n627), .A3(new_n798), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n799), .A2(new_n416), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n800), .A2(new_n612), .A3(new_n600), .A4(new_n614), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n604), .A2(new_n646), .A3(new_n801), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n791), .A2(new_n795), .A3(new_n802), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n694), .A2(new_n690), .A3(new_n696), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n803), .A2(new_n711), .A3(new_n742), .A4(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n684), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n656), .A2(new_n720), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n658), .A2(new_n660), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n602), .A2(new_n652), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n671), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n806), .A2(new_n807), .A3(new_n808), .A4(new_n811), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n656), .B(new_n720), .C1(new_n674), .C2(new_n683), .ZN(new_n813));
  INV_X1    g627(.A(new_n811), .ZN(new_n814));
  OAI21_X1  g628(.A(KEYINPUT52), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n785), .B1(new_n805), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n604), .A2(new_n646), .A3(new_n801), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n818), .A2(new_n794), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n742), .A2(new_n819), .A3(new_n791), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n710), .B(new_n689), .C1(new_n707), .C2(new_n708), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n804), .B1(new_n821), .B2(new_n616), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n812), .A2(new_n815), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(KEYINPUT53), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n817), .A2(new_n825), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n826), .A2(KEYINPUT54), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n826), .A2(KEYINPUT54), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n784), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n826), .A2(KEYINPUT54), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n826), .A2(KEYINPUT54), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n830), .A2(KEYINPUT115), .A3(new_n831), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT51), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n762), .A2(new_n651), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n709), .A2(new_n689), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT50), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n659), .A2(new_n334), .ZN(new_n838));
  OR3_X1    g652(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n837), .B1(new_n836), .B2(new_n838), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n775), .A2(new_n613), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n844), .B1(new_n769), .B2(new_n770), .ZN(new_n845));
  INV_X1    g659(.A(new_n758), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n845), .A2(new_n709), .A3(new_n846), .A4(new_n835), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n839), .A2(KEYINPUT116), .A3(new_n840), .ZN(new_n848));
  AND4_X1   g662(.A1(new_n834), .A2(new_n843), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n689), .ZN(new_n850));
  INV_X1    g664(.A(new_n729), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n852), .A2(new_n547), .A3(new_n340), .A4(new_n670), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n853), .A2(KEYINPUT117), .ZN(new_n854));
  INV_X1    g668(.A(new_n626), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n853), .A2(KEYINPUT117), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n854), .A2(new_n507), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n852), .A2(new_n835), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n789), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n847), .A2(new_n841), .A3(new_n861), .ZN(new_n862));
  AOI22_X1  g676(.A1(new_n849), .A2(new_n861), .B1(KEYINPUT51), .B2(new_n862), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n854), .A2(new_n679), .A3(new_n856), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n859), .A2(new_n728), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT48), .ZN(new_n866));
  INV_X1    g680(.A(new_n631), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n866), .B(new_n337), .C1(new_n867), .C2(new_n836), .ZN(new_n868));
  NOR4_X1   g682(.A1(new_n833), .A2(new_n863), .A3(new_n864), .A4(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(G952), .A2(G953), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n783), .B1(new_n869), .B2(new_n870), .ZN(G75));
  NAND2_X1  g685(.A1(new_n336), .A2(G953), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n872), .B(KEYINPUT119), .Z(new_n873));
  AOI21_X1  g687(.A(new_n410), .B1(new_n817), .B2(new_n825), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT56), .B1(new_n874), .B2(G210), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n404), .A2(new_n408), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(new_n407), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(KEYINPUT55), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n873), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n874), .B(KEYINPUT118), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(new_n413), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT56), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n879), .B1(new_n881), .B2(new_n883), .ZN(G51));
  INV_X1    g698(.A(new_n749), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n880), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(KEYINPUT120), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n599), .B(KEYINPUT57), .Z(new_n888));
  OAI21_X1  g702(.A(new_n888), .B1(new_n827), .B2(new_n828), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n889), .B1(new_n589), .B2(new_n583), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT120), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n880), .A2(new_n891), .A3(new_n885), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n887), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n893), .A2(new_n873), .ZN(G54));
  INV_X1    g708(.A(new_n873), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n880), .A2(KEYINPUT58), .A3(G475), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n502), .A2(new_n503), .ZN(new_n897));
  OR2_X1    g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n896), .A2(new_n897), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n895), .B1(new_n898), .B2(new_n899), .ZN(G60));
  AND2_X1   g714(.A1(new_n618), .A2(new_n622), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT121), .Z(new_n902));
  NAND2_X1  g716(.A1(G478), .A2(G902), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT59), .Z(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n902), .B1(new_n833), .B2(new_n905), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n905), .B(new_n902), .C1(new_n827), .C2(new_n828), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT122), .B1(new_n907), .B2(new_n873), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n873), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT122), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n906), .A2(new_n908), .A3(new_n911), .ZN(G63));
  NAND2_X1  g726(.A1(G217), .A2(G902), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT60), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT53), .B1(new_n823), .B2(new_n824), .ZN(new_n916));
  NOR4_X1   g730(.A1(new_n816), .A2(new_n820), .A3(new_n785), .A4(new_n822), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT123), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n826), .A2(KEYINPUT123), .A3(new_n915), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n920), .A2(new_n542), .A3(new_n921), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n643), .B(KEYINPUT124), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(KEYINPUT123), .B1(new_n826), .B2(new_n915), .ZN(new_n925));
  AOI211_X1 g739(.A(new_n919), .B(new_n914), .C1(new_n817), .C2(new_n825), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n920), .A2(new_n921), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n930), .A2(KEYINPUT125), .A3(new_n924), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n895), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(KEYINPUT126), .B1(new_n929), .B2(new_n931), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n922), .B(new_n932), .C1(new_n933), .C2(KEYINPUT61), .ZN(new_n934));
  AOI21_X1  g748(.A(KEYINPUT125), .B1(new_n930), .B2(new_n924), .ZN(new_n935));
  AOI211_X1 g749(.A(new_n928), .B(new_n923), .C1(new_n920), .C2(new_n921), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n873), .B(new_n922), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT126), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n939), .B1(new_n935), .B2(new_n936), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n937), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n934), .A2(new_n941), .ZN(G66));
  OAI21_X1  g756(.A(G953), .B1(new_n388), .B2(new_n343), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n711), .A2(new_n804), .A3(new_n802), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n943), .B1(new_n945), .B2(G953), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n876), .B1(G898), .B2(new_n460), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT127), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n946), .B(new_n948), .ZN(G69));
  NAND2_X1  g763(.A1(new_n487), .A2(new_n489), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n272), .B(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n813), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n742), .A2(new_n745), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n757), .A2(new_n728), .A3(new_n809), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n766), .A2(new_n773), .A3(new_n954), .A4(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n952), .B1(new_n956), .B2(new_n460), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(G227), .B2(new_n460), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n953), .A2(new_n672), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT62), .Z(new_n960));
  NOR2_X1   g774(.A1(new_n663), .A2(new_n851), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n961), .A2(new_n547), .A3(new_n333), .A4(new_n799), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n960), .A2(new_n766), .A3(new_n773), .A4(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n963), .A2(new_n460), .A3(new_n952), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n649), .B1(new_n952), .B2(new_n566), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n958), .B(new_n964), .C1(new_n460), .C2(new_n965), .ZN(G72));
  NAND2_X1  g780(.A1(G472), .A2(G902), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT63), .Z(new_n968));
  OAI21_X1  g782(.A(new_n968), .B1(new_n956), .B2(new_n944), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n969), .A2(new_n263), .A3(new_n665), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n826), .A2(new_n273), .A3(new_n666), .A4(new_n968), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n970), .A2(new_n873), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n968), .B1(new_n963), .B2(new_n944), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n972), .B1(new_n667), .B2(new_n973), .ZN(G57));
endmodule


