//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 1 0 1 0 1 1 0 1 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0 0 1 1 0 0 0 0 1 1 1 0 0 1 0 1 1 1 1 0 0 0 1 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n786, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014;
  INV_X1    g000(.A(KEYINPUT75), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT32), .ZN(new_n188));
  NOR3_X1   g002(.A1(new_n188), .A2(G472), .A3(G902), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT0), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT66), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(G143), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT65), .B(G146), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n195), .B1(new_n196), .B2(G143), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(KEYINPUT65), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G146), .ZN(new_n200));
  AND4_X1   g014(.A1(KEYINPUT66), .A2(new_n198), .A3(new_n200), .A4(G143), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n192), .B1(new_n197), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT11), .ZN(new_n203));
  INV_X1    g017(.A(G134), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(G137), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(G137), .ZN(new_n206));
  INV_X1    g020(.A(G137), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(KEYINPUT11), .A3(G134), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n205), .A2(new_n206), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G131), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT67), .B(G131), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n211), .A2(new_n205), .A3(new_n206), .A4(new_n208), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G143), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(G146), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n216), .B1(new_n196), .B2(G143), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT64), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n218), .B1(KEYINPUT0), .B2(G128), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n190), .A2(new_n191), .A3(KEYINPUT64), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n192), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n202), .A2(new_n213), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT69), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT69), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n226), .A2(new_n228), .A3(G128), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n230), .B1(new_n197), .B2(new_n201), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT70), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n198), .A2(new_n200), .A3(G143), .ZN(new_n233));
  INV_X1    g047(.A(new_n195), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n196), .A2(KEYINPUT66), .A3(G143), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT70), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n237), .A2(new_n238), .A3(new_n230), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n226), .A2(new_n228), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n233), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G128), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(KEYINPUT71), .A3(new_n217), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT71), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n191), .B1(new_n233), .B2(new_n240), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n198), .A2(new_n200), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n215), .B1(new_n246), .B2(new_n214), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n244), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n232), .A2(new_n239), .B1(new_n243), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n207), .A2(G134), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n250), .A2(new_n206), .A3(new_n251), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n252), .B(G131), .C1(new_n251), .C2(new_n250), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(new_n212), .ZN(new_n254));
  OAI211_X1 g068(.A(KEYINPUT30), .B(new_n224), .C1(new_n249), .C2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G119), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G116), .ZN(new_n257));
  INV_X1    g071(.A(G116), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G119), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT2), .B(G113), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n260), .B(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n255), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n265));
  AOI211_X1 g079(.A(KEYINPUT70), .B(new_n229), .C1(new_n235), .C2(new_n236), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n238), .B1(new_n237), .B2(new_n230), .ZN(new_n267));
  AOI21_X1  g081(.A(KEYINPUT71), .B1(new_n242), .B2(new_n217), .ZN(new_n268));
  NOR3_X1   g082(.A1(new_n245), .A2(new_n247), .A3(new_n244), .ZN(new_n269));
  OAI22_X1  g083(.A1(new_n266), .A2(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n254), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n223), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n265), .B1(new_n272), .B2(KEYINPUT30), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n224), .B1(new_n249), .B2(new_n254), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT30), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n274), .A2(KEYINPUT72), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n264), .B1(new_n273), .B2(new_n276), .ZN(new_n277));
  AOI211_X1 g091(.A(new_n223), .B(new_n263), .C1(new_n270), .C2(new_n271), .ZN(new_n278));
  NOR2_X1   g092(.A1(G237), .A2(G953), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G210), .ZN(new_n280));
  XOR2_X1   g094(.A(new_n280), .B(KEYINPUT27), .Z(new_n281));
  XNOR2_X1  g095(.A(KEYINPUT26), .B(G101), .ZN(new_n282));
  XOR2_X1   g096(.A(new_n281), .B(new_n282), .Z(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n278), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(KEYINPUT73), .B1(new_n277), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n262), .B1(new_n272), .B2(KEYINPUT30), .ZN(new_n288));
  NOR3_X1   g102(.A1(new_n272), .A2(new_n265), .A3(KEYINPUT30), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT72), .B1(new_n274), .B2(new_n275), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT73), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n291), .A2(new_n292), .A3(new_n285), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n287), .A2(new_n293), .A3(KEYINPUT31), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT28), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n274), .A2(new_n263), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n224), .B(new_n262), .C1(new_n249), .C2(new_n254), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT74), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n297), .A2(new_n299), .A3(new_n295), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n299), .B1(new_n297), .B2(new_n295), .ZN(new_n302));
  NOR3_X1   g116(.A1(new_n298), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n291), .A2(new_n285), .ZN(new_n304));
  OAI22_X1  g118(.A1(new_n283), .A2(new_n303), .B1(new_n304), .B2(KEYINPUT31), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n189), .B1(new_n294), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n284), .B1(new_n277), .B2(new_n278), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT29), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n270), .A2(new_n271), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n262), .B1(new_n309), .B2(new_n224), .ZN(new_n310));
  OAI21_X1  g124(.A(KEYINPUT28), .B1(new_n310), .B2(new_n278), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n297), .A2(new_n295), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT74), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n311), .A2(new_n283), .A3(new_n300), .A4(new_n313), .ZN(new_n314));
  AND3_X1   g128(.A1(new_n307), .A2(new_n308), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G902), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n316), .B1(new_n314), .B2(new_n308), .ZN(new_n317));
  OAI21_X1  g131(.A(G472), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n306), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n277), .A2(new_n286), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT31), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n311), .A2(new_n300), .A3(new_n313), .ZN(new_n322));
  AOI22_X1  g136(.A1(new_n320), .A2(new_n321), .B1(new_n322), .B2(new_n284), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n287), .A2(new_n293), .A3(KEYINPUT31), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(G472), .A2(G902), .ZN(new_n326));
  AOI21_X1  g140(.A(KEYINPUT32), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n187), .B1(new_n319), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n325), .A2(new_n326), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n188), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n298), .A2(new_n302), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n331), .A2(KEYINPUT29), .A3(new_n283), .A4(new_n300), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n314), .A2(new_n308), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n283), .B1(new_n291), .B2(new_n297), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n316), .B(new_n332), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n325), .A2(new_n189), .B1(new_n335), .B2(G472), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n330), .A2(new_n336), .A3(KEYINPUT75), .ZN(new_n337));
  INV_X1    g151(.A(G125), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT78), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G125), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT16), .ZN(new_n343));
  INV_X1    g157(.A(G140), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(G125), .A2(G140), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n346), .B1(new_n342), .B2(G140), .ZN(new_n347));
  OAI211_X1 g161(.A(G146), .B(new_n345), .C1(new_n347), .C2(new_n343), .ZN(new_n348));
  AND2_X1   g162(.A1(G125), .A2(G140), .ZN(new_n349));
  OR2_X1    g163(.A1(new_n349), .A2(new_n346), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n196), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT77), .B1(new_n256), .B2(G128), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT23), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n256), .A2(G128), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n191), .A2(G119), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT23), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n355), .A2(KEYINPUT77), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n353), .A2(new_n354), .A3(new_n357), .ZN(new_n358));
  OR2_X1    g172(.A1(new_n358), .A2(G110), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT79), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n355), .A2(new_n354), .ZN(new_n361));
  XNOR2_X1  g175(.A(KEYINPUT24), .B(G110), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n359), .A2(new_n360), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n360), .B1(new_n359), .B2(new_n363), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n348), .B(new_n351), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n345), .B1(new_n347), .B2(new_n343), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n194), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n348), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n358), .A2(G110), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n369), .B(new_n370), .C1(new_n361), .C2(new_n362), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  XNOR2_X1  g186(.A(KEYINPUT22), .B(G137), .ZN(new_n373));
  INV_X1    g187(.A(G221), .ZN(new_n374));
  INV_X1    g188(.A(G234), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n374), .A2(new_n375), .A3(G953), .ZN(new_n376));
  XOR2_X1   g190(.A(new_n373), .B(new_n376), .Z(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n372), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n377), .B1(new_n366), .B2(new_n371), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(KEYINPUT76), .B(G217), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n382), .B1(G234), .B2(new_n316), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n383), .A2(G902), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(KEYINPUT25), .B1(new_n381), .B2(new_n316), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT25), .ZN(new_n387));
  NOR4_X1   g201(.A1(new_n379), .A2(new_n380), .A3(new_n387), .A4(G902), .ZN(new_n388));
  OR2_X1    g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n385), .B1(new_n389), .B2(new_n383), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n328), .A2(new_n337), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT80), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n328), .A2(new_n337), .A3(KEYINPUT80), .A4(new_n390), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G107), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n396), .A2(G104), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(G104), .ZN(new_n398));
  OR2_X1    g212(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n397), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(G101), .ZN(new_n401));
  AND2_X1   g215(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n402));
  NOR2_X1   g216(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n403));
  OAI211_X1 g217(.A(G104), .B(new_n396), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n400), .A2(new_n401), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT82), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT82), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n400), .A2(new_n407), .A3(new_n404), .A4(new_n401), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  OR2_X1    g223(.A1(new_n398), .A2(KEYINPUT83), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n398), .A2(KEYINPUT83), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT84), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n412), .B1(new_n396), .B2(G104), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n397), .A2(KEYINPUT84), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n410), .A2(new_n411), .A3(new_n413), .A4(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G101), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n409), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT85), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI22_X1  g233(.A1(new_n406), .A2(new_n408), .B1(G101), .B2(new_n415), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT85), .ZN(new_n421));
  INV_X1    g235(.A(G113), .ZN(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT89), .B(KEYINPUT5), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n422), .B1(new_n260), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT90), .ZN(new_n425));
  XOR2_X1   g239(.A(KEYINPUT89), .B(KEYINPUT5), .Z(new_n426));
  INV_X1    g240(.A(new_n257), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NOR3_X1   g242(.A1(new_n423), .A2(KEYINPUT90), .A3(new_n257), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n424), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n260), .ZN(new_n431));
  OR2_X1    g245(.A1(new_n431), .A2(new_n261), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n419), .A2(new_n421), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n400), .A2(new_n404), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G101), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT4), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n406), .A2(new_n408), .B1(G101), .B2(new_n435), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n438), .B1(new_n439), .B2(new_n437), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n263), .ZN(new_n441));
  XNOR2_X1  g255(.A(G110), .B(G122), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n434), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  AOI221_X4 g257(.A(new_n418), .B1(new_n415), .B2(G101), .C1(new_n406), .C2(new_n408), .ZN(new_n444));
  AOI21_X1  g258(.A(KEYINPUT85), .B1(new_n409), .B2(new_n416), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n446), .A2(new_n433), .B1(new_n263), .B2(new_n440), .ZN(new_n447));
  XOR2_X1   g261(.A(new_n442), .B(KEYINPUT91), .Z(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  OAI211_X1 g263(.A(KEYINPUT6), .B(new_n443), .C1(new_n447), .C2(new_n449), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n202), .A2(new_n222), .A3(new_n342), .ZN(new_n451));
  XNOR2_X1  g265(.A(KEYINPUT78), .B(G125), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n451), .B1(new_n270), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(G224), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n454), .A2(G953), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n453), .B(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT92), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n434), .A2(new_n441), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT6), .ZN(new_n459));
  AND4_X1   g273(.A1(new_n457), .A2(new_n458), .A3(new_n459), .A4(new_n448), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n449), .B1(new_n434), .B2(new_n441), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n457), .B1(new_n461), .B2(new_n459), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n450), .B(new_n456), .C1(new_n460), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n417), .A2(new_n433), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n422), .B1(new_n260), .B2(KEYINPUT5), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n465), .B1(new_n428), .B2(new_n429), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n432), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n420), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n442), .B(KEYINPUT8), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n464), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n451), .ZN(new_n471));
  INV_X1    g285(.A(new_n455), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(KEYINPUT7), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n471), .B(new_n473), .C1(new_n249), .C2(new_n342), .ZN(new_n474));
  OR2_X1    g288(.A1(new_n472), .A2(KEYINPUT93), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n472), .A2(KEYINPUT93), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n475), .A2(KEYINPUT7), .A3(new_n476), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n470), .B(new_n474), .C1(new_n453), .C2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT94), .ZN(new_n479));
  AOI22_X1  g293(.A1(new_n478), .A2(new_n479), .B1(new_n447), .B2(new_n442), .ZN(new_n480));
  OR2_X1    g294(.A1(new_n453), .A2(new_n477), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n481), .A2(KEYINPUT94), .A3(new_n474), .A4(new_n470), .ZN(new_n482));
  AOI21_X1  g296(.A(G902), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n463), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(G210), .B1(G237), .B2(G902), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n463), .A2(new_n483), .A3(new_n485), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(G214), .B1(G237), .B2(G902), .ZN(new_n490));
  XOR2_X1   g304(.A(new_n490), .B(KEYINPUT87), .Z(new_n491));
  XOR2_X1   g305(.A(new_n491), .B(KEYINPUT88), .Z(new_n492));
  INV_X1    g306(.A(G952), .ZN(new_n493));
  AOI211_X1 g307(.A(G953), .B(new_n493), .C1(G234), .C2(G237), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(KEYINPUT21), .B(G898), .ZN(new_n496));
  XOR2_X1   g310(.A(new_n496), .B(KEYINPUT100), .Z(new_n497));
  INV_X1    g311(.A(G237), .ZN(new_n498));
  OAI211_X1 g312(.A(G902), .B(G953), .C1(new_n375), .C2(new_n498), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n499), .B(KEYINPUT99), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n495), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  AND2_X1   g315(.A1(new_n492), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n489), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(G469), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n267), .A2(new_n266), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n191), .B1(new_n216), .B2(KEYINPUT1), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n237), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n420), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT10), .ZN(new_n509));
  AND2_X1   g323(.A1(new_n202), .A2(new_n222), .ZN(new_n510));
  AOI22_X1  g324(.A1(new_n508), .A2(new_n509), .B1(new_n440), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n213), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n419), .A2(KEYINPUT10), .A3(new_n270), .A4(new_n421), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(G110), .B(G140), .ZN(new_n515));
  INV_X1    g329(.A(G953), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(G227), .ZN(new_n517));
  XOR2_X1   g331(.A(new_n515), .B(new_n517), .Z(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n249), .A2(new_n417), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n508), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n520), .B1(new_n522), .B2(new_n213), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT86), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n524), .A2(KEYINPUT12), .ZN(new_n525));
  AOI211_X1 g339(.A(new_n512), .B(new_n525), .C1(new_n508), .C2(new_n521), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n514), .B(new_n519), .C1(new_n523), .C2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n508), .A2(new_n509), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n440), .A2(new_n510), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(new_n513), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n213), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n519), .B1(new_n532), .B2(new_n514), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n504), .B(new_n316), .C1(new_n528), .C2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n514), .B1(new_n523), .B2(new_n526), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n518), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n532), .A2(new_n514), .A3(new_n519), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(G469), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(G469), .A2(G902), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n534), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT9), .B(G234), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n374), .B1(new_n542), .B2(new_n316), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(G475), .A2(G902), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n546), .B(KEYINPUT98), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n547), .A2(KEYINPUT20), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT96), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT19), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n350), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n346), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n553), .B1(new_n452), .B2(new_n344), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n552), .B(new_n196), .C1(new_n554), .C2(new_n551), .ZN(new_n555));
  INV_X1    g369(.A(new_n211), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n279), .A2(G143), .A3(G214), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(G143), .B1(new_n279), .B2(G214), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n556), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n498), .A2(new_n516), .A3(G214), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n214), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n562), .A2(new_n211), .A3(new_n557), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n348), .A2(new_n555), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT18), .ZN(new_n566));
  INV_X1    g380(.A(G131), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n568), .B1(new_n558), .B2(new_n559), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n562), .B(new_n557), .C1(new_n566), .C2(new_n567), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OAI211_X1 g385(.A(G146), .B(new_n553), .C1(new_n452), .C2(new_n344), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT95), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n572), .A2(new_n573), .B1(new_n196), .B2(new_n350), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n347), .A2(KEYINPUT95), .A3(G146), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n571), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n550), .B1(new_n565), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n574), .A2(new_n575), .ZN(new_n578));
  INV_X1    g392(.A(new_n571), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n348), .A2(new_n555), .A3(new_n564), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n580), .A2(KEYINPUT96), .A3(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(G113), .B(G122), .ZN(new_n583));
  INV_X1    g397(.A(G104), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n583), .B(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n577), .A2(new_n582), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT17), .ZN(new_n588));
  OR2_X1    g402(.A1(new_n560), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n560), .A2(new_n588), .A3(new_n563), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n368), .A2(new_n589), .A3(new_n348), .A4(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n591), .A2(new_n580), .A3(new_n585), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n549), .B1(new_n587), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n587), .A2(new_n592), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT97), .ZN(new_n595));
  INV_X1    g409(.A(new_n547), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT97), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n587), .A2(new_n597), .A3(new_n592), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n595), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n593), .B1(new_n599), .B2(KEYINPUT20), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n591), .A2(new_n580), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n586), .ZN(new_n602));
  AOI21_X1  g416(.A(G902), .B1(new_n602), .B2(new_n592), .ZN(new_n603));
  INV_X1    g417(.A(G475), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(G122), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(G116), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n258), .A2(G122), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(new_n396), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n214), .A2(G128), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT13), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n191), .A2(G143), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n612), .A2(new_n613), .ZN(new_n617));
  OAI21_X1  g431(.A(G134), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n612), .A2(new_n615), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n204), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n611), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n619), .B(new_n204), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n610), .A2(new_n396), .ZN(new_n623));
  OR2_X1    g437(.A1(new_n609), .A2(KEYINPUT14), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n609), .A2(KEYINPUT14), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n624), .A2(new_n625), .A3(new_n608), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(G107), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n622), .A2(new_n623), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n621), .A2(new_n628), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n382), .A2(new_n541), .A3(G953), .ZN(new_n630));
  XOR2_X1   g444(.A(new_n629), .B(new_n630), .Z(new_n631));
  INV_X1    g445(.A(G478), .ZN(new_n632));
  OR2_X1    g446(.A1(new_n632), .A2(KEYINPUT15), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n631), .A2(new_n316), .A3(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n633), .B1(new_n631), .B2(new_n316), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n606), .A2(new_n637), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n503), .A2(new_n545), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n395), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G101), .ZN(G3));
  INV_X1    g455(.A(G472), .ZN(new_n642));
  AOI21_X1  g456(.A(G902), .B1(new_n323), .B2(new_n324), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n329), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n390), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n644), .A2(new_n545), .A3(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT101), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n487), .A2(new_n647), .A3(new_n488), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n463), .A2(new_n483), .A3(KEYINPUT101), .A4(new_n485), .ZN(new_n649));
  INV_X1    g463(.A(new_n491), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(new_n631), .B(KEYINPUT33), .Z(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(G478), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n631), .A2(new_n632), .A3(new_n316), .ZN(new_n654));
  NAND2_X1  g468(.A1(G478), .A2(G902), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n606), .A2(new_n658), .ZN(new_n659));
  AND4_X1   g473(.A1(new_n501), .A2(new_n648), .A3(new_n651), .A4(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n646), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(KEYINPUT102), .ZN(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT34), .B(G104), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G6));
  NAND4_X1  g478(.A1(new_n595), .A2(KEYINPUT103), .A3(new_n598), .A4(new_n548), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n665), .B1(new_n604), .B2(new_n603), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n599), .A2(KEYINPUT20), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT103), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n595), .A2(new_n598), .A3(new_n548), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n637), .ZN(new_n672));
  AND3_X1   g486(.A1(new_n667), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  AND4_X1   g487(.A1(new_n501), .A2(new_n648), .A3(new_n651), .A4(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n646), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT105), .B(G107), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(KEYINPUT104), .B(KEYINPUT35), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G9));
  INV_X1    g493(.A(new_n644), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n383), .B1(new_n386), .B2(new_n388), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n372), .B(KEYINPUT106), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n682), .B1(KEYINPUT36), .B2(new_n378), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n372), .B(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n378), .A2(KEYINPUT36), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n683), .A2(new_n384), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n681), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n639), .A2(new_n680), .A3(new_n689), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT37), .B(G110), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G12));
  NOR2_X1   g506(.A1(new_n500), .A2(G900), .ZN(new_n693));
  OR2_X1    g507(.A1(new_n693), .A2(KEYINPUT107), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(KEYINPUT107), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n694), .A2(new_n495), .A3(new_n695), .ZN(new_n696));
  AND4_X1   g510(.A1(new_n672), .A2(new_n667), .A3(new_n671), .A4(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n697), .A2(new_n648), .A3(new_n651), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n545), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n328), .A2(new_n337), .A3(new_n701), .A4(new_n689), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n191), .ZN(G30));
  XNOR2_X1  g518(.A(new_n696), .B(KEYINPUT39), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n545), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(KEYINPUT40), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n284), .B1(new_n310), .B2(new_n278), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n287), .A2(new_n293), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g524(.A(G472), .B1(new_n710), .B2(G902), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n330), .A2(new_n306), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT109), .B(KEYINPUT38), .ZN(new_n713));
  XOR2_X1   g527(.A(new_n489), .B(new_n713), .Z(new_n714));
  NOR4_X1   g528(.A1(new_n689), .A2(new_n606), .A3(new_n491), .A4(new_n637), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n708), .A2(new_n712), .A3(new_n714), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G143), .ZN(G45));
  INV_X1    g531(.A(new_n702), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n648), .A2(new_n651), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n656), .B1(new_n652), .B2(G478), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n720), .B(new_n696), .C1(new_n600), .C2(new_n605), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n718), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G146), .ZN(G48));
  NOR2_X1   g540(.A1(new_n531), .A2(new_n213), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n512), .B1(new_n511), .B2(new_n513), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n518), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n527), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n504), .B1(new_n730), .B2(new_n316), .ZN(new_n731));
  AOI211_X1 g545(.A(G469), .B(G902), .C1(new_n729), .C2(new_n527), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n733), .A2(new_n390), .A3(new_n544), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n660), .A2(new_n328), .A3(new_n337), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(KEYINPUT41), .B(G113), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G15));
  NAND4_X1  g551(.A1(new_n674), .A2(new_n328), .A3(new_n337), .A4(new_n734), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G116), .ZN(G18));
  AND2_X1   g553(.A1(new_n328), .A2(new_n337), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT110), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n733), .A2(new_n544), .A3(new_n606), .A4(new_n637), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n648), .A2(new_n651), .A3(new_n501), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n740), .A2(new_n741), .A3(new_n689), .A4(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n328), .A2(new_n337), .A3(new_n689), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n742), .A2(new_n743), .ZN(new_n747));
  OAI21_X1  g561(.A(KEYINPUT110), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  XOR2_X1   g563(.A(KEYINPUT111), .B(G119), .Z(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(G21));
  NOR2_X1   g565(.A1(new_n606), .A2(new_n637), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n733), .A2(new_n544), .A3(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n743), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n643), .A2(new_n642), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n322), .A2(new_n284), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n324), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(KEYINPUT112), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n320), .A2(new_n321), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT112), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n324), .A2(new_n756), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n758), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n755), .B1(new_n762), .B2(new_n326), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n754), .A2(new_n390), .A3(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G122), .ZN(G24));
  NAND2_X1  g579(.A1(new_n762), .A2(new_n326), .ZN(new_n766));
  INV_X1    g580(.A(new_n755), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(new_n767), .A3(new_n689), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n731), .A2(new_n732), .A3(new_n543), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n719), .A2(new_n722), .A3(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(new_n338), .ZN(G27));
  INV_X1    g586(.A(KEYINPUT42), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n539), .B(KEYINPUT113), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n538), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n544), .B1(new_n775), .B2(new_n732), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n487), .A2(new_n488), .A3(new_n650), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n328), .A2(new_n337), .A3(new_n390), .A4(new_n778), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n773), .B1(new_n779), .B2(new_n721), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n776), .A2(new_n777), .A3(new_n721), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n330), .A2(new_n336), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n781), .A2(KEYINPUT42), .A3(new_n782), .A4(new_n390), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G131), .ZN(G33));
  INV_X1    g599(.A(new_n697), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n779), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(new_n204), .ZN(G36));
  NAND2_X1  g602(.A1(new_n536), .A2(new_n537), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT45), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n504), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n791), .B1(new_n790), .B2(new_n789), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n774), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT46), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n732), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n792), .A2(KEYINPUT46), .A3(new_n774), .ZN(new_n796));
  AOI211_X1 g610(.A(new_n543), .B(new_n706), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  XOR2_X1   g611(.A(new_n777), .B(KEYINPUT114), .Z(new_n798));
  NAND2_X1  g612(.A1(new_n606), .A2(new_n720), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT43), .ZN(new_n800));
  INV_X1    g614(.A(new_n689), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n800), .A2(new_n680), .A3(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT44), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR4_X1   g618(.A1(new_n800), .A2(new_n680), .A3(KEYINPUT44), .A4(new_n801), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n797), .B(new_n798), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G137), .ZN(G39));
  AOI21_X1  g621(.A(new_n543), .B1(new_n795), .B2(new_n796), .ZN(new_n808));
  XOR2_X1   g622(.A(KEYINPUT115), .B(KEYINPUT47), .Z(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n777), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n645), .A3(new_n722), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n740), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT115), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n814), .A2(KEYINPUT47), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n810), .B(new_n813), .C1(new_n808), .C2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G140), .ZN(G42));
  XOR2_X1   g631(.A(new_n733), .B(KEYINPUT49), .Z(new_n818));
  NAND3_X1  g632(.A1(new_n390), .A2(new_n492), .A3(new_n544), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n819), .A2(new_n799), .ZN(new_n820));
  OR4_X1    g634(.A1(new_n712), .A2(new_n818), .A3(new_n714), .A4(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n800), .A2(new_n495), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n822), .A2(new_n769), .A3(new_n811), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n782), .A2(new_n390), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XOR2_X1   g639(.A(new_n825), .B(KEYINPUT48), .Z(new_n826));
  INV_X1    g640(.A(new_n769), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n390), .A2(new_n494), .ZN(new_n828));
  NOR4_X1   g642(.A1(new_n712), .A2(new_n827), .A3(new_n777), .A4(new_n828), .ZN(new_n829));
  AOI211_X1 g643(.A(new_n493), .B(G953), .C1(new_n829), .C2(new_n659), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n719), .A2(new_n769), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n822), .A2(new_n390), .A3(new_n763), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n826), .B(new_n830), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n829), .A2(new_n606), .A3(new_n658), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n834), .B1(new_n768), .B2(new_n823), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n810), .B1(new_n808), .B2(new_n815), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n733), .A2(new_n543), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n832), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n798), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n835), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n714), .A2(new_n650), .A3(new_n827), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n839), .B(new_n843), .C1(KEYINPUT118), .C2(KEYINPUT50), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n839), .A2(new_n843), .ZN(new_n845));
  XOR2_X1   g659(.A(KEYINPUT118), .B(KEYINPUT50), .Z(new_n846));
  OAI21_X1  g660(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(KEYINPUT51), .B1(new_n842), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n833), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n840), .B1(new_n838), .B2(KEYINPUT120), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n850), .B1(KEYINPUT120), .B2(new_n838), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT51), .B1(new_n835), .B2(KEYINPUT119), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n852), .B1(KEYINPUT119), .B2(new_n835), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n851), .A2(new_n847), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n849), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n698), .B(KEYINPUT108), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n771), .B1(new_n718), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n719), .A2(new_n752), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n801), .A2(new_n696), .ZN(new_n859));
  INV_X1    g673(.A(new_n776), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n306), .A2(new_n711), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n859), .B(new_n860), .C1(new_n327), .C2(new_n861), .ZN(new_n862));
  OAI22_X1  g676(.A1(new_n702), .A2(new_n723), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT52), .B1(new_n857), .B2(new_n864), .ZN(new_n865));
  OAI22_X1  g679(.A1(new_n700), .A2(new_n702), .B1(new_n768), .B2(new_n770), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT52), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n866), .A2(new_n863), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n637), .A2(new_n696), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n870), .B1(new_n681), .B2(new_n688), .ZN(new_n871));
  INV_X1    g685(.A(new_n598), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n597), .B1(new_n587), .B2(new_n592), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT103), .B1(new_n874), .B2(new_n548), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n666), .B1(new_n875), .B2(new_n668), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n871), .A2(new_n876), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n545), .A2(new_n877), .A3(new_n777), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n878), .A2(new_n328), .A3(new_n337), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n763), .A2(new_n781), .A3(new_n689), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n879), .B(new_n880), .C1(new_n779), .C2(new_n786), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n881), .B1(new_n780), .B2(new_n783), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n600), .A2(new_n605), .A3(new_n637), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n463), .A2(new_n483), .A3(new_n485), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n485), .B1(new_n463), .B2(new_n483), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n883), .B(new_n502), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(KEYINPUT116), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT116), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n489), .A2(new_n888), .A3(new_n502), .A4(new_n883), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n489), .A2(new_n659), .A3(new_n502), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n887), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n646), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n764), .A2(new_n738), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n735), .A2(new_n690), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n882), .A2(new_n640), .A3(new_n749), .A4(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT53), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n869), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n895), .A2(new_n640), .A3(new_n749), .ZN(new_n899));
  INV_X1    g713(.A(new_n787), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n879), .A2(new_n880), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n784), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n857), .A2(new_n864), .A3(KEYINPUT52), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n867), .B1(new_n866), .B2(new_n863), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT53), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT54), .B1(new_n898), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT117), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n897), .B1(new_n869), .B2(new_n896), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT54), .ZN(new_n911));
  INV_X1    g725(.A(new_n899), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n912), .A2(new_n906), .A3(KEYINPUT53), .A4(new_n882), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n910), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n908), .A2(new_n909), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n911), .B1(new_n910), .B2(new_n913), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(KEYINPUT117), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n855), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(G952), .A2(G953), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT121), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n821), .B1(new_n918), .B2(new_n920), .ZN(G75));
  AOI21_X1  g735(.A(new_n316), .B1(new_n910), .B2(new_n913), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(G210), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n450), .B1(new_n460), .B2(new_n462), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(new_n456), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT55), .ZN(new_n926));
  XNOR2_X1  g740(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n923), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n516), .A2(G952), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT56), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n926), .B1(new_n923), .B2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n931), .A2(new_n933), .ZN(G51));
  XNOR2_X1  g748(.A(new_n774), .B(KEYINPUT123), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT57), .Z(new_n936));
  AND3_X1   g750(.A1(new_n910), .A2(new_n911), .A3(new_n913), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n936), .B1(new_n937), .B2(new_n916), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n730), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n792), .B(KEYINPUT124), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n922), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n929), .B1(new_n939), .B2(new_n941), .ZN(G54));
  AND2_X1   g756(.A1(KEYINPUT58), .A2(G475), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n922), .A2(new_n874), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n874), .B1(new_n922), .B2(new_n943), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n944), .A2(new_n945), .A3(new_n929), .ZN(G60));
  XOR2_X1   g760(.A(new_n655), .B(KEYINPUT59), .Z(new_n947));
  NOR2_X1   g761(.A1(new_n652), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n948), .B1(new_n937), .B2(new_n916), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n930), .ZN(new_n950));
  INV_X1    g764(.A(new_n947), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n915), .A2(new_n917), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n950), .B1(new_n652), .B2(new_n952), .ZN(G63));
  NAND2_X1  g767(.A1(new_n910), .A2(new_n913), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n683), .A2(new_n687), .ZN(new_n955));
  NAND2_X1  g769(.A1(G217), .A2(G902), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT60), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n954), .A2(new_n955), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n957), .B1(new_n910), .B2(new_n913), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n959), .B(new_n930), .C1(new_n381), .C2(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(KEYINPUT61), .B1(new_n959), .B2(KEYINPUT125), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OR2_X1    g777(.A1(new_n960), .A2(new_n381), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n929), .B1(new_n960), .B2(new_n955), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT125), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n966), .B1(new_n960), .B2(new_n955), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n964), .B(new_n965), .C1(new_n967), .C2(KEYINPUT61), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n963), .A2(new_n968), .ZN(G66));
  INV_X1    g783(.A(new_n497), .ZN(new_n970));
  OAI21_X1  g784(.A(G953), .B1(new_n970), .B2(new_n454), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n971), .B1(new_n912), .B2(G953), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n924), .B1(G898), .B2(new_n516), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n972), .B(new_n973), .ZN(G69));
  AOI21_X1  g788(.A(new_n866), .B1(new_n718), .B2(new_n724), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n716), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(KEYINPUT62), .ZN(new_n977));
  OR2_X1    g791(.A1(new_n659), .A2(new_n883), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n395), .A2(new_n707), .A3(new_n811), .A4(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT126), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n979), .B(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT62), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n975), .A2(new_n982), .A3(new_n716), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n816), .A2(new_n806), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n977), .A2(new_n981), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n516), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n255), .B1(new_n289), .B2(new_n290), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n552), .B1(new_n554), .B2(new_n551), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n858), .A2(new_n824), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n787), .B1(new_n797), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n816), .A2(new_n806), .A3(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(new_n784), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n857), .A2(new_n725), .ZN(new_n995));
  NOR3_X1   g809(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(new_n516), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n990), .B1(G900), .B2(G953), .ZN(new_n998));
  AOI22_X1  g812(.A1(new_n986), .A2(new_n990), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n516), .B1(G227), .B2(G900), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n997), .A2(new_n998), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n1000), .B1(new_n1001), .B2(KEYINPUT127), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n999), .B(new_n1002), .ZN(G72));
  NAND2_X1  g817(.A1(G472), .A2(G902), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1004), .B(KEYINPUT63), .Z(new_n1005));
  INV_X1    g819(.A(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1006), .B1(new_n996), .B2(new_n912), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n277), .A2(new_n278), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1008), .A2(new_n284), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n930), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n287), .A2(new_n307), .A3(new_n293), .ZN(new_n1011));
  AND3_X1   g825(.A1(new_n954), .A2(new_n1005), .A3(new_n1011), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1005), .B1(new_n985), .B2(new_n899), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n1008), .A2(new_n284), .ZN(new_n1014));
  AOI211_X1 g828(.A(new_n1010), .B(new_n1012), .C1(new_n1013), .C2(new_n1014), .ZN(G57));
endmodule


