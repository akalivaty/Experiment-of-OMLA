//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 1 0 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1 1 0 1 1 0 1 0 0 0 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1232, new_n1233, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1303, new_n1304;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  AND2_X1   g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G20), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n202), .A2(G50), .ZN(new_n213));
  INV_X1    g0013(.A(G50), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G97), .ZN(new_n216));
  INV_X1    g0016(.A(G257), .ZN(new_n217));
  OAI22_X1  g0017(.A1(new_n214), .A2(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n218), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  AND2_X1   g0021(.A1(KEYINPUT64), .A2(G68), .ZN(new_n222));
  NOR2_X1   g0022(.A1(KEYINPUT64), .A2(G68), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n219), .B(new_n220), .C1(new_n221), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT65), .Z(new_n227));
  OAI21_X1  g0027(.A(new_n207), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n210), .B1(new_n212), .B2(new_n213), .C1(new_n228), .C2(KEYINPUT1), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT67), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G226), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n234), .B(new_n235), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n239), .B(KEYINPUT68), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n236), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(G1), .A2(G13), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(KEYINPUT69), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT69), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n249), .A2(new_n253), .A3(new_n250), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G20), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n256), .B1(new_n201), .B2(new_n214), .ZN(new_n257));
  XOR2_X1   g0057(.A(new_n257), .B(KEYINPUT70), .Z(new_n258));
  XOR2_X1   g0058(.A(KEYINPUT8), .B(G58), .Z(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(G20), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n259), .A2(new_n261), .B1(G150), .B2(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n255), .B1(new_n258), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G13), .ZN(new_n265));
  NOR3_X1   g0065(.A1(new_n265), .A2(new_n256), .A3(G1), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n264), .B1(new_n214), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n266), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n255), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G1), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G20), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n270), .A2(G50), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g0074(.A(new_n274), .B(KEYINPUT9), .ZN(new_n275));
  INV_X1    g0075(.A(G41), .ZN(new_n276));
  INV_X1    g0076(.A(G45), .ZN(new_n277));
  AOI21_X1  g0077(.A(G1), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(G1), .A3(G13), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n278), .A2(new_n280), .A3(G274), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n271), .B1(G41), .B2(G45), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n281), .B1(new_n215), .B2(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT3), .B(G33), .ZN(new_n285));
  NOR2_X1   g0085(.A1(G222), .A2(G1698), .ZN(new_n286));
  INV_X1    g0086(.A(G1698), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(G223), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n285), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT3), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G77), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n280), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n284), .B1(new_n289), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G200), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n298), .B1(G190), .B2(new_n296), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n275), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT10), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT10), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n275), .A2(new_n302), .A3(new_n299), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n296), .A2(G169), .ZN(new_n305));
  INV_X1    g0105(.A(new_n274), .ZN(new_n306));
  INV_X1    g0106(.A(G179), .ZN(new_n307));
  AOI211_X1 g0107(.A(new_n305), .B(new_n306), .C1(new_n307), .C2(new_n296), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G232), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G1698), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n285), .B(new_n311), .C1(G226), .C2(G1698), .ZN(new_n312));
  NAND2_X1  g0112(.A1(G33), .A2(G97), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n280), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n281), .B1(new_n221), .B2(new_n283), .ZN(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT13), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NOR3_X1   g0117(.A1(new_n314), .A2(KEYINPUT13), .A3(new_n315), .ZN(new_n318));
  OAI21_X1  g0118(.A(G169), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT14), .ZN(new_n320));
  INV_X1    g0120(.A(new_n314), .ZN(new_n321));
  INV_X1    g0121(.A(new_n315), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT13), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT72), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n318), .A2(KEYINPUT72), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n326), .A2(new_n327), .A3(G179), .A4(new_n316), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT14), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n329), .B(G169), .C1(new_n317), .C2(new_n318), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n320), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n255), .ZN(new_n332));
  INV_X1    g0132(.A(new_n224), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n333), .A2(new_n256), .ZN(new_n334));
  INV_X1    g0134(.A(new_n262), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n256), .A2(G33), .ZN(new_n336));
  OAI22_X1  g0136(.A1(new_n335), .A2(new_n214), .B1(new_n336), .B2(new_n294), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n332), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT11), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT11), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n332), .B(new_n340), .C1(new_n334), .C2(new_n337), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(G68), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n343), .B1(new_n271), .B2(G20), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n255), .A2(new_n268), .A3(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT73), .ZN(new_n346));
  XNOR2_X1  g0146(.A(new_n345), .B(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(KEYINPUT12), .B1(new_n266), .B2(new_n343), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n265), .A2(G1), .ZN(new_n349));
  AND2_X1   g0149(.A1(new_n349), .A2(KEYINPUT12), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n348), .B1(new_n334), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n342), .A2(new_n347), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n331), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n297), .B1(new_n324), .B2(new_n316), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT74), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n326), .A2(new_n327), .A3(G190), .A4(new_n316), .ZN(new_n357));
  AND3_X1   g0157(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n356), .B1(new_n355), .B2(new_n357), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n353), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n259), .A2(new_n262), .B1(G20), .B2(G77), .ZN(new_n362));
  XNOR2_X1  g0162(.A(KEYINPUT15), .B(G87), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n362), .B1(new_n336), .B2(new_n363), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n364), .A2(new_n332), .B1(new_n294), .B2(new_n266), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n270), .A2(G77), .A3(new_n272), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n280), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n285), .A2(new_n287), .ZN(new_n369));
  INV_X1    g0169(.A(G107), .ZN(new_n370));
  OAI22_X1  g0170(.A1(new_n369), .A2(new_n310), .B1(new_n370), .B2(new_n285), .ZN(new_n371));
  NOR3_X1   g0171(.A1(new_n293), .A2(new_n221), .A3(new_n287), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n368), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n281), .ZN(new_n374));
  INV_X1    g0174(.A(new_n283), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n374), .B1(G244), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n367), .B1(G200), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n377), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n378), .A2(KEYINPUT71), .B1(G190), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(KEYINPUT71), .B2(new_n378), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n307), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n382), .B(new_n367), .C1(G169), .C2(new_n379), .ZN(new_n383));
  AND2_X1   g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n304), .A2(new_n309), .A3(new_n361), .A4(new_n384), .ZN(new_n385));
  AND2_X1   g0185(.A1(new_n259), .A2(new_n272), .ZN(new_n386));
  INV_X1    g0186(.A(new_n259), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n270), .A2(new_n386), .B1(new_n266), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(G20), .B1(new_n290), .B2(new_n292), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT75), .B1(new_n389), .B2(KEYINPUT7), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT75), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT7), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n391), .B(new_n392), .C1(new_n285), .C2(G20), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n293), .A2(KEYINPUT7), .A3(new_n256), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n390), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(G68), .ZN(new_n396));
  INV_X1    g0196(.A(G159), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n335), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(G58), .B1(new_n222), .B2(new_n223), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT76), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI211_X1 g0201(.A(KEYINPUT76), .B(G58), .C1(new_n222), .C2(new_n223), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n401), .A2(new_n202), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n398), .B1(new_n403), .B2(G20), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n396), .A2(KEYINPUT16), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n332), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n256), .A2(KEYINPUT7), .ZN(new_n407));
  AOI21_X1  g0207(.A(KEYINPUT77), .B1(new_n260), .B2(KEYINPUT3), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n260), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n407), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n389), .A2(KEYINPUT7), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n333), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(KEYINPUT16), .B1(new_n404), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n388), .B1(new_n406), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(G169), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT78), .ZN(new_n418));
  OR2_X1    g0218(.A1(G223), .A2(G1698), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n215), .A2(G1698), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n290), .A2(new_n419), .A3(new_n292), .A4(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(G33), .A2(G87), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n368), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n280), .A2(G232), .A3(new_n282), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n281), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n418), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n280), .B1(new_n421), .B2(new_n422), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n281), .A2(new_n425), .ZN(new_n429));
  NOR3_X1   g0229(.A1(new_n428), .A2(new_n429), .A3(KEYINPUT78), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n417), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n428), .A2(new_n429), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n307), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n416), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT18), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n403), .A2(G20), .ZN(new_n439));
  INV_X1    g0239(.A(new_n398), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n414), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT16), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n443), .A2(new_n332), .A3(new_n405), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n434), .B1(new_n444), .B2(new_n388), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT18), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n438), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n297), .B1(new_n427), .B2(new_n430), .ZN(new_n448));
  INV_X1    g0248(.A(G190), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n432), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n451), .B(new_n388), .C1(new_n406), .C2(new_n415), .ZN(new_n452));
  NOR2_X1   g0252(.A1(KEYINPUT79), .A2(KEYINPUT17), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g0254(.A(KEYINPUT79), .B(KEYINPUT17), .Z(new_n455));
  NAND4_X1  g0255(.A1(new_n444), .A2(new_n388), .A3(new_n451), .A4(new_n455), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n447), .A2(new_n457), .ZN(new_n458));
  OR2_X1    g0258(.A1(new_n385), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT4), .ZN(new_n460));
  INV_X1    g0260(.A(G244), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n460), .B1(new_n369), .B2(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n285), .A2(KEYINPUT4), .A3(G244), .A4(new_n287), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n285), .A2(G250), .A3(G1698), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G283), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n462), .A2(new_n463), .A3(new_n464), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n368), .ZN(new_n467));
  XNOR2_X1  g0267(.A(KEYINPUT5), .B(G41), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n277), .A2(G1), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n280), .A2(G274), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n368), .B1(new_n469), .B2(new_n468), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G257), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n467), .A2(new_n449), .A3(new_n473), .A4(new_n475), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n467), .A2(new_n473), .A3(new_n475), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n476), .B1(new_n477), .B2(G200), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n268), .A2(G97), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n271), .A2(G33), .ZN(new_n480));
  XNOR2_X1  g0280(.A(new_n480), .B(KEYINPUT82), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n269), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n479), .B1(new_n483), .B2(G97), .ZN(new_n484));
  OAI21_X1  g0284(.A(G107), .B1(new_n412), .B2(new_n413), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT80), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI211_X1 g0287(.A(KEYINPUT80), .B(G107), .C1(new_n412), .C2(new_n413), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n370), .A2(KEYINPUT6), .A3(G97), .ZN(new_n489));
  XOR2_X1   g0289(.A(G97), .B(G107), .Z(new_n490));
  OAI21_X1  g0290(.A(new_n489), .B1(new_n490), .B2(KEYINPUT6), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n491), .A2(G20), .B1(G77), .B2(new_n262), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n487), .A2(new_n488), .A3(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT81), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n493), .A2(new_n494), .A3(new_n332), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n494), .B1(new_n493), .B2(new_n332), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n478), .B(new_n484), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n484), .ZN(new_n499));
  INV_X1    g0299(.A(new_n497), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n499), .B1(new_n500), .B2(new_n495), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n477), .A2(new_n307), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n467), .A2(new_n473), .A3(new_n475), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n417), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n498), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n474), .A2(G264), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n285), .A2(G250), .A3(new_n287), .ZN(new_n508));
  NAND2_X1  g0308(.A1(G33), .A2(G294), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT85), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n285), .A2(new_n511), .A3(G257), .A4(G1698), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n290), .A2(new_n292), .A3(G257), .A4(G1698), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT85), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n510), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n473), .B(new_n507), .C1(new_n515), .C2(new_n280), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(G200), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n514), .A2(new_n512), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n368), .B1(new_n518), .B2(new_n510), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n519), .A2(G190), .A3(new_n473), .A4(new_n507), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n483), .A2(G107), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n266), .A2(new_n370), .ZN(new_n522));
  XOR2_X1   g0322(.A(new_n522), .B(KEYINPUT25), .Z(new_n523));
  AND2_X1   g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g0324(.A(KEYINPUT83), .B(G116), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n525), .A2(new_n260), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT23), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n527), .B1(new_n256), .B2(G107), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n370), .A2(KEYINPUT23), .A3(G20), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n526), .A2(new_n256), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT24), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n290), .A2(new_n292), .A3(new_n256), .A4(G87), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(KEYINPUT22), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT22), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n285), .A2(new_n534), .A3(new_n256), .A4(G87), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n530), .A2(new_n531), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n531), .B1(new_n530), .B2(new_n536), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n332), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n517), .A2(new_n520), .A3(new_n524), .A4(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT86), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n530), .A2(new_n536), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(KEYINPUT24), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n255), .B1(new_n545), .B2(new_n537), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n521), .A2(new_n523), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n548), .A2(KEYINPUT86), .A3(new_n517), .A4(new_n520), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n543), .A2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT19), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n256), .B1(new_n313), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(G87), .B2(new_n205), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n290), .A2(new_n292), .A3(new_n256), .A4(G68), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n551), .B1(new_n336), .B2(new_n216), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n332), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n255), .A2(new_n481), .A3(G87), .A4(new_n268), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n363), .A2(new_n266), .ZN(new_n559));
  AND3_X1   g0359(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n280), .B(G250), .C1(G1), .C2(new_n277), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n280), .A2(G274), .A3(new_n469), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n285), .A2(G238), .A3(new_n287), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n285), .A2(G244), .A3(G1698), .ZN(new_n565));
  INV_X1    g0365(.A(G116), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT83), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT83), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(G116), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G33), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n564), .A2(new_n565), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n563), .B1(new_n572), .B2(new_n368), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(G190), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n560), .B(new_n574), .C1(new_n297), .C2(new_n573), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n572), .A2(new_n368), .ZN(new_n576));
  INV_X1    g0376(.A(new_n563), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n417), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n573), .A2(new_n307), .ZN(new_n580));
  INV_X1    g0380(.A(new_n363), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n255), .A2(new_n481), .A3(new_n268), .A4(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n557), .A2(new_n559), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n579), .A2(new_n580), .A3(new_n583), .ZN(new_n584));
  AND3_X1   g0384(.A1(new_n575), .A2(new_n584), .A3(KEYINPUT84), .ZN(new_n585));
  AOI21_X1  g0385(.A(KEYINPUT84), .B1(new_n575), .B2(new_n584), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT21), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n255), .A2(new_n481), .A3(G116), .A4(new_n268), .ZN(new_n589));
  INV_X1    g0389(.A(new_n349), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n525), .A2(G20), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n465), .B(new_n256), .C1(G33), .C2(new_n216), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n592), .A2(new_n251), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n593), .A2(KEYINPUT20), .A3(new_n591), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT20), .B1(new_n593), .B2(new_n591), .ZN(new_n595));
  OAI221_X1 g0395(.A(new_n589), .B1(new_n590), .B2(new_n591), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n472), .B1(G270), .B2(new_n474), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n285), .A2(G264), .A3(G1698), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n293), .A2(G303), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n599), .B(new_n600), .C1(new_n369), .C2(new_n217), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n368), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(G169), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n588), .B1(new_n597), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(G200), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n598), .A2(new_n602), .A3(G190), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n597), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n598), .A2(new_n602), .A3(G179), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n596), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n596), .A2(KEYINPUT21), .A3(G169), .A4(new_n603), .ZN(new_n612));
  AND4_X1   g0412(.A1(new_n605), .A2(new_n608), .A3(new_n611), .A4(new_n612), .ZN(new_n613));
  OR2_X1    g0413(.A1(new_n516), .A2(G179), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n524), .A2(new_n540), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n516), .A2(new_n417), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n550), .A2(new_n587), .A3(new_n613), .A4(new_n617), .ZN(new_n618));
  NOR3_X1   g0418(.A1(new_n459), .A2(new_n506), .A3(new_n618), .ZN(G372));
  INV_X1    g0419(.A(new_n459), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n501), .A2(new_n505), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n587), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(KEYINPUT26), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n579), .A2(KEYINPUT87), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n579), .A2(KEYINPUT87), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n580), .B(new_n583), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n575), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n621), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n623), .B1(KEYINPUT26), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n605), .A2(new_n611), .A3(new_n612), .ZN(new_n631));
  INV_X1    g0431(.A(new_n617), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n628), .B(new_n550), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n626), .B1(new_n633), .B2(new_n506), .ZN(new_n634));
  OR2_X1    g0434(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n620), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n454), .A2(new_n456), .ZN(new_n637));
  INV_X1    g0437(.A(new_n383), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n638), .B1(new_n358), .B2(new_n359), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n637), .B1(new_n639), .B2(new_n353), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n438), .A2(KEYINPUT88), .A3(new_n446), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT88), .ZN(new_n642));
  AOI211_X1 g0442(.A(new_n437), .B(new_n434), .C1(new_n444), .C2(new_n388), .ZN(new_n643));
  AOI21_X1  g0443(.A(KEYINPUT18), .B1(new_n416), .B2(new_n435), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n304), .B1(new_n640), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n636), .A2(new_n309), .A3(new_n647), .ZN(G369));
  OR2_X1    g0448(.A1(new_n613), .A2(KEYINPUT89), .ZN(new_n649));
  OR3_X1    g0449(.A1(new_n590), .A2(KEYINPUT27), .A3(G20), .ZN(new_n650));
  OAI21_X1  g0450(.A(KEYINPUT27), .B1(new_n590), .B2(G20), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(G213), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(G343), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n597), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n613), .A2(KEYINPUT89), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n649), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n631), .A2(new_n656), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT90), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(G330), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n632), .A2(new_n655), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n543), .A2(new_n549), .B1(new_n615), .B2(new_n654), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n665), .B1(new_n666), .B2(new_n632), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n631), .A2(new_n655), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n671), .B1(new_n632), .B2(new_n655), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n669), .A2(new_n672), .ZN(G399));
  INV_X1    g0473(.A(new_n208), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(G41), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n205), .A2(G87), .A3(G116), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G1), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n213), .B2(new_n676), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n679), .B(KEYINPUT28), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT29), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n635), .A2(new_n681), .A3(new_n655), .ZN(new_n682));
  INV_X1    g0482(.A(new_n506), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n587), .A2(new_n613), .A3(new_n617), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n683), .A2(new_n684), .A3(new_n550), .A4(new_n655), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n467), .A2(new_n475), .A3(new_n573), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n519), .A2(new_n507), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n686), .A2(new_n687), .A3(new_n609), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(KEYINPUT30), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT30), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n610), .A2(new_n507), .A3(new_n519), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n690), .B1(new_n691), .B2(new_n686), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n573), .A2(G179), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n503), .A2(new_n516), .A3(new_n693), .A4(new_n603), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n689), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n695), .A2(KEYINPUT31), .A3(new_n654), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(KEYINPUT31), .B1(new_n695), .B2(new_n654), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n685), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(G330), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n629), .A2(KEYINPUT26), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(KEYINPUT26), .B2(new_n622), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n655), .B1(new_n703), .B2(new_n634), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(KEYINPUT29), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n682), .A2(new_n701), .A3(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n680), .B1(new_n707), .B2(G1), .ZN(G364));
  NOR2_X1   g0508(.A1(new_n265), .A2(G20), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n271), .B1(new_n709), .B2(G45), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n675), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n712), .B1(new_n663), .B2(G330), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(G330), .B2(new_n663), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n250), .B1(G20), .B2(new_n417), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n256), .A2(new_n307), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  OR3_X1    g0518(.A1(new_n718), .A2(KEYINPUT93), .A3(new_n297), .ZN(new_n719));
  OAI21_X1  g0519(.A(KEYINPUT93), .B1(new_n718), .B2(new_n297), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n719), .A2(G190), .A3(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n297), .A2(G190), .ZN(new_n723));
  OAI21_X1  g0523(.A(G20), .B1(new_n723), .B2(G179), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT95), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  AOI22_X1  g0529(.A1(new_n722), .A2(G326), .B1(new_n729), .B2(G294), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n719), .A2(new_n449), .A3(new_n720), .ZN(new_n731));
  XOR2_X1   g0531(.A(KEYINPUT33), .B(G317), .Z(new_n732));
  OAI21_X1  g0532(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(G190), .A2(G200), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n717), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(G311), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n256), .A2(G179), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n734), .ZN(new_n738));
  INV_X1    g0538(.A(G329), .ZN(new_n739));
  OAI22_X1  g0539(.A1(new_n735), .A2(new_n736), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n737), .A2(G190), .A3(G200), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n740), .B1(G303), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n718), .A2(new_n723), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n285), .B1(new_n744), .B2(G322), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n737), .A2(new_n449), .A3(G200), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(KEYINPUT94), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(G283), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n743), .B(new_n745), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n729), .A2(G97), .ZN(new_n751));
  OAI221_X1 g0551(.A(new_n751), .B1(new_n214), .B2(new_n721), .C1(new_n343), .C2(new_n731), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n747), .A2(G107), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n738), .A2(new_n397), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n754), .B(KEYINPUT32), .ZN(new_n755));
  INV_X1    g0555(.A(new_n735), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n293), .B1(new_n756), .B2(G77), .ZN(new_n757));
  AOI22_X1  g0557(.A1(G58), .A2(new_n744), .B1(new_n742), .B2(G87), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n753), .A2(new_n755), .A3(new_n757), .A4(new_n758), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n733), .A2(new_n750), .B1(new_n752), .B2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT96), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n716), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n762), .B1(new_n761), .B2(new_n760), .ZN(new_n763));
  INV_X1    g0563(.A(new_n712), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n674), .A2(new_n293), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT91), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n766), .A2(G355), .B1(new_n566), .B2(new_n674), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n247), .A2(G45), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT92), .Z(new_n769));
  NOR2_X1   g0569(.A1(new_n674), .A2(new_n285), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n770), .B1(G45), .B2(new_n213), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n767), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G13), .A2(G33), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G20), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n715), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n764), .B1(new_n772), .B2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n775), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n763), .B(new_n777), .C1(new_n663), .C2(new_n778), .ZN(new_n779));
  AND2_X1   g0579(.A1(new_n714), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(G396));
  NAND2_X1  g0581(.A1(new_n635), .A2(new_n655), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n367), .A2(new_n654), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n381), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n383), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n383), .A2(new_n654), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n782), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n786), .B1(new_n784), .B2(new_n383), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n655), .B(new_n790), .C1(new_n630), .C2(new_n634), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n712), .B1(new_n792), .B2(new_n701), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(new_n701), .B2(new_n792), .ZN(new_n794));
  AOI22_X1  g0594(.A1(G143), .A2(new_n744), .B1(new_n756), .B2(G159), .ZN(new_n795));
  INV_X1    g0595(.A(G150), .ZN(new_n796));
  INV_X1    g0596(.A(G137), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n795), .B1(new_n731), .B2(new_n796), .C1(new_n797), .C2(new_n721), .ZN(new_n798));
  XOR2_X1   g0598(.A(new_n798), .B(KEYINPUT34), .Z(new_n799));
  NAND2_X1  g0599(.A1(new_n747), .A2(G68), .ZN(new_n800));
  INV_X1    g0600(.A(G132), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n285), .B1(new_n738), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(G50), .B2(new_n742), .ZN(new_n803));
  INV_X1    g0603(.A(G58), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n800), .B(new_n803), .C1(new_n804), .C2(new_n728), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n747), .A2(G87), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n285), .B1(new_n744), .B2(G294), .ZN(new_n807));
  INV_X1    g0607(.A(new_n738), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(G311), .ZN(new_n809));
  AOI22_X1  g0609(.A1(G107), .A2(new_n742), .B1(new_n756), .B2(new_n570), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n806), .A2(new_n807), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G303), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n751), .B1(new_n749), .B2(new_n731), .C1(new_n812), .C2(new_n721), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n799), .A2(new_n805), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(new_n715), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n715), .A2(new_n773), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n764), .B1(new_n294), .B2(new_n816), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n815), .B(new_n817), .C1(new_n790), .C2(new_n774), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n794), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(G384));
  NOR2_X1   g0620(.A1(new_n212), .A2(new_n566), .ZN(new_n821));
  XOR2_X1   g0621(.A(new_n491), .B(KEYINPUT97), .Z(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT35), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n821), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(new_n824), .B2(new_n823), .ZN(new_n826));
  XNOR2_X1  g0626(.A(KEYINPUT98), .B(KEYINPUT36), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n826), .B(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n213), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n401), .A2(new_n829), .A3(G77), .A4(new_n402), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n214), .A2(G68), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n271), .B(G13), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n828), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n353), .A2(new_n654), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT101), .ZN(new_n836));
  AOI21_X1  g0636(.A(KEYINPUT16), .B1(new_n396), .B2(new_n404), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n388), .B1(new_n406), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n652), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n643), .A2(new_n644), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n841), .B1(new_n842), .B2(new_n637), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n416), .A2(new_n839), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n436), .A2(new_n844), .A3(new_n452), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT37), .ZN(new_n846));
  INV_X1    g0646(.A(new_n452), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n847), .A2(new_n846), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n838), .B1(new_n435), .B2(new_n839), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n845), .A2(new_n846), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n843), .A2(new_n850), .A3(KEYINPUT38), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT39), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT100), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n844), .A2(new_n642), .A3(new_n452), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(KEYINPUT37), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n845), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n652), .B1(new_n444), .B2(new_n388), .ZN(new_n858));
  NOR3_X1   g0658(.A1(new_n847), .A2(new_n445), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n859), .A2(KEYINPUT37), .A3(new_n855), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n641), .A2(new_n645), .A3(new_n457), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n861), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n854), .B1(new_n863), .B2(KEYINPUT38), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n857), .A2(new_n860), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n862), .A2(new_n858), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT38), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n867), .A2(KEYINPUT100), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n853), .B1(new_n864), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n840), .B1(new_n447), .B2(new_n457), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n849), .A2(KEYINPUT37), .A3(new_n452), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n859), .B2(KEYINPUT37), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n868), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n851), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT99), .B1(new_n875), .B2(KEYINPUT39), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT99), .ZN(new_n877));
  AOI211_X1 g0677(.A(new_n877), .B(new_n852), .C1(new_n874), .C2(new_n851), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n836), .B1(new_n870), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n851), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT38), .B1(new_n843), .B2(new_n850), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT39), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n877), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n875), .A2(KEYINPUT99), .A3(KEYINPUT39), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n853), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT100), .B1(new_n867), .B2(new_n868), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n854), .B(KEYINPUT38), .C1(new_n865), .C2(new_n866), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n886), .A2(new_n890), .A3(KEYINPUT101), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n835), .B1(new_n880), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n791), .A2(new_n787), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n352), .A2(new_n654), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n360), .A2(new_n895), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n353), .B(new_n894), .C1(new_n358), .C2(new_n359), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n900), .A2(new_n875), .B1(new_n646), .B2(new_n652), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n892), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n459), .B1(new_n682), .B2(new_n705), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n647), .A2(new_n309), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n903), .B(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n851), .B1(new_n888), .B2(new_n889), .ZN(new_n908));
  NOR3_X1   g0708(.A1(new_n618), .A2(new_n506), .A3(new_n654), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n695), .A2(new_n654), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT31), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n696), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n898), .B(new_n790), .C1(new_n909), .C2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(KEYINPUT40), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n914), .A2(KEYINPUT103), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT103), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n700), .A2(new_n919), .A3(new_n790), .A4(new_n898), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n918), .A2(new_n920), .A3(new_n875), .ZN(new_n921));
  XNOR2_X1  g0721(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n908), .A2(new_n917), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n923), .A2(new_n620), .A3(new_n700), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(G330), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n923), .B1(new_n620), .B2(new_n700), .ZN(new_n926));
  OR2_X1    g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n907), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n271), .B2(new_n709), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n907), .A2(new_n927), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n833), .B1(new_n929), .B2(new_n930), .ZN(G367));
  NAND2_X1  g0731(.A1(new_n239), .A2(new_n770), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n932), .B(new_n776), .C1(new_n208), .C2(new_n363), .ZN(new_n933));
  AOI22_X1  g0733(.A1(G58), .A2(new_n742), .B1(new_n756), .B2(G50), .ZN(new_n934));
  INV_X1    g0734(.A(new_n744), .ZN(new_n935));
  OAI221_X1 g0735(.A(new_n934), .B1(new_n294), .B2(new_n746), .C1(new_n796), .C2(new_n935), .ZN(new_n936));
  AOI211_X1 g0736(.A(new_n293), .B(new_n936), .C1(G137), .C2(new_n808), .ZN(new_n937));
  INV_X1    g0737(.A(new_n731), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(G159), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n729), .A2(G68), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n722), .A2(G143), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n937), .A2(new_n939), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n742), .A2(KEYINPUT46), .A3(G116), .ZN(new_n943));
  INV_X1    g0743(.A(G317), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n943), .B1(new_n944), .B2(new_n738), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n935), .A2(new_n812), .B1(new_n216), .B2(new_n746), .ZN(new_n946));
  AOI21_X1  g0746(.A(KEYINPUT46), .B1(new_n742), .B2(new_n570), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n293), .B1(new_n735), .B2(new_n749), .ZN(new_n948));
  NOR4_X1   g0748(.A1(new_n945), .A2(new_n946), .A3(new_n947), .A4(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(G294), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n949), .B1(new_n950), .B2(new_n731), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n721), .A2(new_n736), .B1(new_n728), .B2(new_n370), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n942), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n953), .B(KEYINPUT47), .Z(new_n954));
  OAI211_X1 g0754(.A(new_n712), .B(new_n933), .C1(new_n954), .C2(new_n716), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT109), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n655), .A2(new_n560), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n628), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n626), .B2(new_n957), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n956), .B1(new_n778), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n501), .A2(new_n655), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n484), .B1(new_n496), .B2(new_n497), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n962), .A2(new_n502), .A3(new_n504), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n506), .A2(new_n961), .B1(new_n963), .B2(new_n655), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n671), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT42), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n964), .B(KEYINPUT104), .Z(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n632), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n963), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n966), .B1(new_n969), .B2(new_n655), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT105), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(KEYINPUT43), .B2(new_n959), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n959), .B(KEYINPUT43), .Z(new_n973));
  OAI21_X1  g0773(.A(new_n972), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n967), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n669), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n974), .B(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n672), .A2(new_n964), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT45), .Z(new_n980));
  NOR2_X1   g0780(.A1(new_n672), .A2(new_n964), .ZN(new_n981));
  OR2_X1    g0781(.A1(KEYINPUT106), .A2(KEYINPUT44), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(KEYINPUT106), .A2(KEYINPUT44), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n981), .B2(new_n982), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n980), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n668), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n667), .B(new_n670), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n664), .B(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n989), .A2(new_n706), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n669), .B(new_n980), .C1(new_n983), .C2(new_n985), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n987), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(KEYINPUT107), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT107), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n987), .A2(new_n994), .A3(new_n990), .A4(new_n991), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n706), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n675), .B(KEYINPUT41), .Z(new_n997));
  OAI21_X1  g0797(.A(new_n710), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT108), .ZN(new_n999));
  AND3_X1   g0799(.A1(new_n978), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n999), .B1(new_n978), .B2(new_n998), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n960), .B1(new_n1000), .B2(new_n1001), .ZN(G387));
  NOR2_X1   g0802(.A1(new_n741), .A2(new_n294), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(G150), .B2(new_n808), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n214), .B2(new_n935), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n293), .B(new_n1005), .C1(G68), .C2(new_n756), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n747), .A2(G97), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n729), .A2(new_n581), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G159), .A2(new_n722), .B1(new_n938), .B2(new_n259), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(G317), .A2(new_n744), .B1(new_n756), .B2(G303), .ZN(new_n1011));
  INV_X1    g0811(.A(G322), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1011), .B1(new_n731), .B2(new_n736), .C1(new_n1012), .C2(new_n721), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT48), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n729), .A2(G283), .B1(G294), .B2(new_n742), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT110), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(KEYINPUT49), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n285), .B1(new_n808), .B2(G326), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1020), .B(new_n1021), .C1(new_n525), .C2(new_n746), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1019), .A2(KEYINPUT49), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1010), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n715), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n236), .A2(new_n277), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n677), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n1026), .A2(new_n770), .B1(new_n1027), .B2(new_n766), .ZN(new_n1028));
  NOR3_X1   g0828(.A1(new_n387), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n677), .B(new_n277), .C1(new_n343), .C2(new_n294), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT50), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(new_n259), .B2(new_n214), .ZN(new_n1032));
  NOR3_X1   g0832(.A1(new_n1029), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n1028), .A2(new_n1033), .B1(G107), .B2(new_n208), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n764), .B1(new_n1034), .B2(new_n776), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1025), .A2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n667), .B2(new_n775), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n664), .B(new_n988), .Z(new_n1038));
  AOI21_X1  g0838(.A(new_n1037), .B1(new_n1038), .B2(new_n711), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1038), .A2(new_n707), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n675), .B1(new_n989), .B2(new_n706), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1039), .B1(new_n1040), .B2(new_n1041), .ZN(G393));
  AOI21_X1  g0842(.A(new_n676), .B1(new_n993), .B2(new_n995), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT111), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(new_n987), .B2(new_n991), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n1044), .B2(new_n991), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1043), .B1(new_n990), .B2(new_n1046), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n721), .A2(new_n796), .B1(new_n397), .B2(new_n935), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT51), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n729), .A2(G77), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n293), .B1(new_n756), .B2(new_n259), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n742), .A2(new_n333), .B1(new_n808), .B2(G143), .ZN(new_n1052));
  AND4_X1   g0852(.A1(new_n806), .A2(new_n1050), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1049), .B(new_n1053), .C1(new_n214), .C2(new_n731), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT113), .Z(new_n1055));
  AOI21_X1  g0855(.A(new_n285), .B1(new_n808), .B2(G322), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n753), .B(new_n1056), .C1(new_n749), .C2(new_n741), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT114), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n721), .A2(new_n944), .B1(new_n736), .B2(new_n935), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT52), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n728), .A2(new_n525), .B1(new_n950), .B2(new_n735), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(G303), .B2(new_n938), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1058), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT115), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n715), .B1(new_n1055), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n776), .B1(new_n216), .B2(new_n208), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n244), .B2(new_n770), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT112), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1065), .A2(new_n712), .A3(new_n1068), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT116), .Z(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n775), .B2(new_n975), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n1046), .B2(new_n711), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1047), .A2(new_n1072), .ZN(G390));
  NAND2_X1  g0873(.A1(new_n899), .A2(new_n835), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n880), .A2(new_n891), .A3(new_n1074), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n700), .A2(G330), .A3(new_n790), .A4(new_n898), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n898), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n655), .B(new_n785), .C1(new_n703), .C2(new_n634), .ZN(new_n1078));
  AND2_X1   g0878(.A1(new_n1078), .A2(new_n787), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n908), .B(new_n835), .C1(new_n1077), .C2(new_n1079), .ZN(new_n1080));
  AND3_X1   g0880(.A1(new_n1075), .A2(new_n1076), .A3(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1076), .B1(new_n1075), .B2(new_n1080), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n790), .B1(new_n701), .B2(KEYINPUT117), .ZN(new_n1084));
  INV_X1    g0884(.A(G330), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n685), .B2(new_n699), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT117), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1077), .B1(new_n1084), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT118), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1076), .A2(new_n1078), .A3(new_n787), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1089), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n788), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n701), .A2(KEYINPUT117), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n898), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(KEYINPUT118), .B1(new_n1096), .B2(new_n1091), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1076), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n700), .A2(G330), .A3(new_n790), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n1099), .A2(new_n1077), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n893), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1093), .A2(new_n1097), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n620), .A2(new_n1086), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  NOR3_X1   g0904(.A1(new_n1104), .A2(new_n904), .A3(new_n905), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n676), .B1(new_n1083), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1075), .A2(new_n1080), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n1098), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1075), .A2(new_n1076), .A3(new_n1080), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1112));
  AOI21_X1  g0912(.A(KEYINPUT119), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  OAI211_X1 g0913(.A(KEYINPUT119), .B(new_n1112), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1107), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n816), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1050), .B1(new_n370), .B2(new_n731), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(G283), .B2(new_n722), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n935), .A2(new_n566), .B1(new_n738), .B2(new_n950), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(G97), .B2(new_n756), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n285), .B1(new_n742), .B2(G87), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n1121), .A2(new_n800), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n293), .B1(new_n744), .B2(G132), .ZN(new_n1124));
  OR3_X1    g0924(.A1(new_n741), .A2(KEYINPUT53), .A3(new_n796), .ZN(new_n1125));
  OAI21_X1  g0925(.A(KEYINPUT53), .B1(new_n741), .B2(new_n796), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(KEYINPUT54), .B(G143), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n735), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(G125), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n746), .A2(new_n214), .B1(new_n738), .B2(new_n1130), .ZN(new_n1131));
  NOR3_X1   g0931(.A1(new_n1127), .A2(new_n1129), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(G128), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n1133), .A2(new_n721), .B1(new_n731), .B2(new_n797), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(G159), .B2(new_n729), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1119), .A2(new_n1123), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n712), .B1(new_n259), .B2(new_n1117), .C1(new_n1136), .C2(new_n716), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n880), .A2(new_n891), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1137), .B1(new_n1139), .B2(new_n773), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT120), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1141), .B1(new_n1111), .B2(new_n710), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1083), .A2(KEYINPUT120), .A3(new_n711), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1140), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1116), .A2(new_n1144), .ZN(G378));
  NAND2_X1  g0945(.A1(new_n304), .A2(new_n309), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n274), .A2(new_n839), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1146), .B(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1148), .B(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n773), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n756), .A2(G137), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n1153), .B1(new_n741), .B2(new_n1128), .C1(new_n935), .C2(new_n1133), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n731), .A2(new_n801), .B1(new_n728), .B2(new_n796), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n1154), .B(new_n1155), .C1(G125), .C2(new_n722), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  AND2_X1   g0957(.A1(new_n1157), .A2(KEYINPUT59), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1157), .A2(KEYINPUT59), .ZN(new_n1159));
  OR2_X1    g0959(.A1(KEYINPUT121), .A2(G124), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(KEYINPUT121), .A2(G124), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n808), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(G33), .A2(G41), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1162), .B(new_n1163), .C1(new_n397), .C2(new_n746), .ZN(new_n1164));
  NOR3_X1   g0964(.A1(new_n1158), .A2(new_n1159), .A3(new_n1164), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(G97), .A2(new_n938), .B1(new_n722), .B2(G116), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n746), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(G58), .A2(new_n1167), .B1(new_n756), .B2(new_n581), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n744), .A2(G107), .B1(new_n808), .B2(G283), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n293), .A2(new_n276), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n1170), .A2(new_n1003), .A3(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1166), .A2(new_n940), .A3(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT58), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1171), .B(new_n214), .C1(G33), .C2(G41), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n715), .B1(new_n1165), .B2(new_n1178), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1179), .B(KEYINPUT122), .Z(new_n1180));
  AOI211_X1 g0980(.A(new_n764), .B(new_n1180), .C1(new_n214), .C2(new_n816), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1152), .A2(new_n1181), .ZN(new_n1182));
  NOR3_X1   g0982(.A1(new_n870), .A2(new_n879), .A3(new_n836), .ZN(new_n1183));
  AOI21_X1  g0983(.A(KEYINPUT101), .B1(new_n886), .B2(new_n890), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n834), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n923), .A2(G330), .A3(new_n1150), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n921), .A2(new_n922), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n881), .B1(new_n864), .B2(new_n869), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1187), .B(G330), .C1(new_n1188), .C2(new_n916), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n1151), .ZN(new_n1190));
  AND4_X1   g0990(.A1(new_n1185), .A2(new_n901), .A3(new_n1186), .A4(new_n1190), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n1185), .A2(new_n901), .B1(new_n1190), .B2(new_n1186), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1182), .B1(new_n1193), .B2(new_n710), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT57), .ZN(new_n1195));
  OAI21_X1  g0995(.A(KEYINPUT123), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1186), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1150), .B1(new_n923), .B2(G330), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n1197), .A2(new_n1198), .B1(new_n892), .B2(new_n902), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT123), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1195), .B1(new_n1196), .B2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1109), .A2(new_n1106), .A3(new_n1110), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n1105), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n676), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1105), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(new_n1083), .B2(new_n1106), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1195), .B1(new_n1207), .B2(new_n1193), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1194), .B1(new_n1205), .B2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(G375));
  OR2_X1    g1010(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n997), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1211), .A2(new_n1212), .A3(new_n1112), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n712), .B1(G68), .B2(new_n1117), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n898), .A2(new_n774), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT124), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1008), .B1(new_n950), .B2(new_n721), .C1(new_n525), .C2(new_n731), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n735), .A2(new_n370), .B1(new_n738), .B2(new_n812), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(G97), .B2(new_n742), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n285), .B1(new_n744), .B2(G283), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1219), .B(new_n1220), .C1(new_n748), .C2(new_n294), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n729), .A2(G50), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n293), .B1(new_n1167), .B2(G58), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n744), .A2(G137), .B1(new_n808), .B2(G128), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(G159), .A2(new_n742), .B1(new_n756), .B2(G150), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .A4(new_n1225), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n801), .A2(new_n721), .B1(new_n731), .B2(new_n1128), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n1217), .A2(new_n1221), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1214), .B(new_n1216), .C1(new_n715), .C2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n1102), .B2(new_n711), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1213), .A2(new_n1230), .ZN(G381));
  NOR4_X1   g1031(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1232), .A2(new_n1230), .A3(new_n1213), .ZN(new_n1233));
  OR4_X1    g1033(.A1(G387), .A2(new_n1233), .A3(G378), .A4(G375), .ZN(G407));
  INV_X1    g1034(.A(G378), .ZN(new_n1235));
  INV_X1    g1035(.A(G213), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1236), .A2(G343), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1209), .A2(new_n1235), .A3(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(G407), .A2(G213), .A3(new_n1238), .ZN(G409));
  XNOR2_X1  g1039(.A(G393), .B(G396), .ZN(new_n1240));
  AND3_X1   g1040(.A1(new_n1047), .A2(new_n1072), .A3(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1240), .B1(new_n1047), .B2(new_n1072), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(G387), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1243), .B(new_n960), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT61), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1112), .A2(KEYINPUT60), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1249), .A2(new_n1211), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n675), .B1(new_n1249), .B2(new_n1211), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1230), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  OR2_X1    g1052(.A1(new_n1252), .A2(new_n819), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n819), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1237), .A2(G2897), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(new_n1255), .B(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n710), .B1(new_n1196), .B2(new_n1201), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(new_n1152), .B2(new_n1181), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1204), .B(new_n1212), .C1(new_n1192), .C2(new_n1191), .ZN(new_n1260));
  AOI21_X1  g1060(.A(G378), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1201), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1185), .A2(new_n901), .A3(new_n1190), .A4(new_n1186), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1200), .B1(new_n1199), .B2(new_n1263), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1204), .B(KEYINPUT57), .C1(new_n1262), .C2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1208), .A2(new_n1265), .A3(new_n675), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1194), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1266), .A2(G378), .A3(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(KEYINPUT125), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT125), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1266), .A2(G378), .A3(new_n1270), .A4(new_n1267), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1261), .B1(new_n1269), .B2(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1257), .B1(new_n1272), .B2(new_n1237), .ZN(new_n1273));
  NOR3_X1   g1073(.A1(new_n1272), .A2(new_n1237), .A3(new_n1255), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT62), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1248), .B(new_n1273), .C1(new_n1274), .C2(new_n1275), .ZN(new_n1276));
  AND2_X1   g1076(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1247), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT126), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1273), .A2(new_n1279), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1257), .B(KEYINPUT126), .C1(new_n1272), .C2(new_n1237), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1261), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1270), .B1(new_n1209), .B2(G378), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1271), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1283), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1237), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1255), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1288), .A2(KEYINPUT63), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1286), .A2(new_n1287), .A3(new_n1289), .ZN(new_n1290));
  AND3_X1   g1090(.A1(new_n1245), .A2(new_n1246), .A3(new_n1248), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1237), .B1(new_n1293), .B2(new_n1283), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT63), .B1(new_n1294), .B2(new_n1288), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1292), .A2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(KEYINPUT127), .B1(new_n1282), .B2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1290), .B(new_n1291), .C1(new_n1274), .C2(KEYINPUT63), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT127), .ZN(new_n1300));
  NOR3_X1   g1100(.A1(new_n1298), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1278), .B1(new_n1297), .B2(new_n1301), .ZN(G405));
  OAI21_X1  g1102(.A(new_n1293), .B1(G378), .B2(new_n1209), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(new_n1303), .B(new_n1255), .ZN(new_n1304));
  XOR2_X1   g1104(.A(new_n1304), .B(new_n1247), .Z(G402));
endmodule


