//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 1 0 1 1 0 1 0 0 0 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n734, new_n735, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n798, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n879, new_n880, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n995,
    new_n996;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(G1gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT91), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT16), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n202), .B1(new_n205), .B2(G1gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n203), .A2(new_n206), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n204), .A2(new_n207), .A3(G8gat), .ZN(new_n208));
  INV_X1    g007(.A(G8gat), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n203), .B(new_n206), .C1(KEYINPUT91), .C2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT92), .ZN(new_n212));
  XOR2_X1   g011(.A(G43gat), .B(G50gat), .Z(new_n213));
  INV_X1    g012(.A(KEYINPUT15), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G29gat), .ZN(new_n216));
  INV_X1    g015(.A(G36gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(new_n217), .A3(KEYINPUT14), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT14), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(G29gat), .B2(G36gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(G29gat), .A2(G36gat), .ZN(new_n221));
  AND3_X1   g020(.A1(new_n218), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G43gat), .B(G50gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT15), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n215), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT90), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT90), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n215), .A2(new_n222), .A3(new_n227), .A4(new_n224), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n222), .A2(new_n224), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n226), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT17), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n226), .A2(KEYINPUT17), .A3(new_n228), .A4(new_n229), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT92), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n208), .A2(new_n234), .A3(new_n210), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n212), .A2(new_n232), .A3(new_n233), .A4(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G229gat), .A2(G233gat), .ZN(new_n237));
  AND3_X1   g036(.A1(new_n211), .A2(new_n230), .A3(KEYINPUT93), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT93), .B1(new_n211), .B2(new_n230), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n236), .B(new_n237), .C1(new_n238), .C2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT18), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  OR2_X1    g041(.A1(new_n238), .A2(new_n239), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n243), .A2(KEYINPUT18), .A3(new_n237), .A4(new_n236), .ZN(new_n244));
  OAI22_X1  g043(.A1(new_n238), .A2(new_n239), .B1(new_n211), .B2(new_n230), .ZN(new_n245));
  XOR2_X1   g044(.A(new_n237), .B(KEYINPUT13), .Z(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(KEYINPUT94), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT94), .B1(new_n245), .B2(new_n246), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n242), .B(new_n244), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  XOR2_X1   g049(.A(G169gat), .B(G197gat), .Z(new_n251));
  XNOR2_X1  g050(.A(G113gat), .B(G141gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XOR2_X1   g054(.A(new_n255), .B(KEYINPUT12), .Z(new_n256));
  NAND2_X1  g055(.A1(new_n250), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n249), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(new_n247), .ZN(new_n259));
  INV_X1    g058(.A(new_n256), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n259), .A2(new_n260), .A3(new_n242), .A4(new_n244), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT88), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n264), .A2(KEYINPUT35), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT78), .ZN(new_n266));
  INV_X1    g065(.A(G113gat), .ZN(new_n267));
  INV_X1    g066(.A(G120gat), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT1), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n269), .B1(new_n267), .B2(new_n268), .ZN(new_n270));
  INV_X1    g069(.A(G127gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(G134gat), .ZN(new_n272));
  OR2_X1    g071(.A1(KEYINPUT65), .A2(G134gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(KEYINPUT65), .A2(G134gat), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n273), .A2(G127gat), .A3(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n272), .B1(new_n275), .B2(KEYINPUT66), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT66), .ZN(new_n277));
  AND2_X1   g076(.A1(KEYINPUT65), .A2(G134gat), .ZN(new_n278));
  NOR2_X1   g077(.A1(KEYINPUT65), .A2(G134gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n277), .B1(new_n280), .B2(G127gat), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n270), .B1(new_n276), .B2(new_n281), .ZN(new_n282));
  XOR2_X1   g081(.A(G127gat), .B(G134gat), .Z(new_n283));
  NOR2_X1   g082(.A1(new_n270), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  AND2_X1   g085(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n288));
  OAI21_X1  g087(.A(G155gat), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT2), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT74), .ZN(new_n291));
  INV_X1    g090(.A(G148gat), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n291), .B1(new_n292), .B2(G141gat), .ZN(new_n293));
  INV_X1    g092(.A(G141gat), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n294), .A2(KEYINPUT74), .A3(G148gat), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n293), .B(new_n295), .C1(new_n294), .C2(G148gat), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT75), .ZN(new_n297));
  INV_X1    g096(.A(G155gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n298), .A2(G162gat), .ZN(new_n299));
  INV_X1    g098(.A(G162gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n300), .A2(G155gat), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n297), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(G155gat), .B(G162gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT75), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n290), .A2(new_n296), .A3(new_n302), .A4(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT3), .ZN(new_n306));
  XNOR2_X1  g105(.A(G141gat), .B(G148gat), .ZN(new_n307));
  OAI22_X1  g106(.A1(new_n307), .A2(KEYINPUT2), .B1(new_n299), .B2(new_n301), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n305), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n306), .B1(new_n305), .B2(new_n308), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT77), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n286), .B(new_n309), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  AOI211_X1 g111(.A(KEYINPUT77), .B(new_n306), .C1(new_n305), .C2(new_n308), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n266), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  AND2_X1   g113(.A1(new_n286), .A2(new_n309), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n305), .A2(new_n308), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT3), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT77), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n310), .A2(new_n311), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n315), .A2(new_n318), .A3(KEYINPUT78), .A4(new_n319), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n282), .A2(new_n308), .A3(new_n305), .A4(new_n285), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT4), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT79), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n316), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n275), .A2(KEYINPUT66), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n280), .A2(new_n277), .A3(G127gat), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n325), .A2(new_n326), .A3(new_n272), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n284), .B1(new_n327), .B2(new_n270), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT4), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n305), .A2(KEYINPUT79), .A3(new_n308), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n324), .A2(new_n328), .A3(new_n329), .A4(new_n330), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n314), .A2(new_n320), .B1(new_n322), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(G225gat), .A2(G233gat), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n334), .A2(KEYINPUT5), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT80), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n314), .A2(new_n320), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n334), .B1(new_n321), .B2(new_n329), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n324), .A2(new_n328), .A3(KEYINPUT4), .A4(new_n330), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n286), .A2(new_n316), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n321), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(new_n334), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT5), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n337), .B1(new_n343), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n341), .B1(new_n314), .B2(new_n320), .ZN(new_n350));
  NOR3_X1   g149(.A1(new_n350), .A2(KEYINPUT80), .A3(new_n347), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n336), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G1gat), .B(G29gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n353), .B(KEYINPUT0), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(G57gat), .ZN(new_n355));
  INV_X1    g154(.A(G85gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n355), .B(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT6), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(KEYINPUT6), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n352), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n343), .A2(new_n337), .A3(new_n348), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT80), .B1(new_n350), .B2(new_n347), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT6), .ZN(new_n365));
  INV_X1    g164(.A(new_n357), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n364), .A2(new_n365), .A3(new_n336), .A4(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n361), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(G226gat), .A2(G233gat), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT25), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NOR3_X1   g172(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT24), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n376), .A2(G183gat), .A3(G190gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(G169gat), .A2(G176gat), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n379));
  AND2_X1   g178(.A1(G183gat), .A2(G190gat), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n377), .B(new_n378), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n371), .B1(new_n375), .B2(new_n381), .ZN(new_n382));
  OR2_X1    g181(.A1(new_n379), .A2(new_n380), .ZN(new_n383));
  NOR2_X1   g182(.A1(G169gat), .A2(G176gat), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT23), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(new_n372), .ZN(new_n387));
  AOI22_X1  g186(.A1(new_n380), .A2(new_n376), .B1(G169gat), .B2(G176gat), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n383), .A2(new_n387), .A3(new_n388), .A4(KEYINPUT25), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n382), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(G183gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT27), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT27), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(G183gat), .ZN(new_n394));
  INV_X1    g193(.A(G190gat), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n392), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n396), .B1(KEYINPUT64), .B2(KEYINPUT28), .ZN(new_n397));
  XNOR2_X1  g196(.A(KEYINPUT27), .B(G183gat), .ZN(new_n398));
  NOR2_X1   g197(.A1(KEYINPUT64), .A2(KEYINPUT28), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n398), .A2(new_n395), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n380), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT26), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n384), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n403), .B1(new_n384), .B2(new_n404), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n397), .A2(new_n400), .A3(new_n401), .A4(new_n405), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n390), .A2(KEYINPUT72), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT72), .B1(new_n390), .B2(new_n406), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n370), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n396), .B(new_n399), .ZN(new_n410));
  AND2_X1   g209(.A1(new_n405), .A2(new_n401), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n410), .A2(new_n411), .B1(new_n382), .B2(new_n389), .ZN(new_n412));
  OAI211_X1 g211(.A(KEYINPUT71), .B(new_n369), .C1(new_n412), .C2(KEYINPUT29), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT71), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT29), .B1(new_n390), .B2(new_n406), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n414), .B1(new_n415), .B2(new_n370), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n409), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(G204gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(G197gat), .ZN(new_n419));
  INV_X1    g218(.A(G197gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(G204gat), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT69), .ZN(new_n422));
  AND3_X1   g221(.A1(new_n419), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n422), .B1(new_n419), .B2(new_n421), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n425), .A2(KEYINPUT70), .ZN(new_n426));
  NAND2_X1  g225(.A1(G211gat), .A2(G218gat), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT22), .ZN(new_n428));
  AND3_X1   g227(.A1(new_n427), .A2(KEYINPUT70), .A3(new_n428), .ZN(new_n429));
  OAI22_X1  g228(.A1(new_n423), .A2(new_n424), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  XOR2_X1   g229(.A(G211gat), .B(G218gat), .Z(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n431), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n419), .A2(new_n421), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT69), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n419), .A2(new_n421), .A3(new_n422), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n425), .B(KEYINPUT70), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n433), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n432), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n417), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n440), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT73), .B1(new_n412), .B2(new_n369), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n390), .A2(new_n406), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT73), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(new_n445), .A3(new_n370), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT72), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n390), .A2(KEYINPUT72), .A3(new_n406), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT29), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n442), .B(new_n447), .C1(new_n451), .C2(new_n370), .ZN(new_n452));
  XNOR2_X1  g251(.A(G8gat), .B(G36gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n453), .B(G64gat), .ZN(new_n454));
  INV_X1    g253(.A(G92gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n441), .A2(new_n452), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT30), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n441), .A2(KEYINPUT30), .A3(new_n452), .A4(new_n456), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n441), .A2(new_n452), .ZN(new_n461));
  INV_X1    g260(.A(new_n456), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n459), .A2(new_n460), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n264), .A2(KEYINPUT35), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n368), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(G227gat), .A2(G233gat), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n412), .A2(new_n328), .ZN(new_n470));
  AOI22_X1  g269(.A1(new_n390), .A2(new_n406), .B1(new_n282), .B2(new_n285), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT67), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n444), .A2(new_n286), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n474), .A2(KEYINPUT67), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n469), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT32), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT33), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  XOR2_X1   g278(.A(G15gat), .B(G43gat), .Z(new_n480));
  XNOR2_X1  g279(.A(G71gat), .B(G99gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n480), .B(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n477), .A2(new_n479), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n482), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n476), .B(KEYINPUT32), .C1(new_n478), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n474), .A2(KEYINPUT67), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n487), .A2(new_n488), .A3(new_n468), .A4(new_n470), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT34), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n444), .A2(new_n286), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n492), .B1(KEYINPUT67), .B2(new_n474), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n493), .A2(KEYINPUT34), .A3(new_n468), .A4(new_n488), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT68), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n486), .A2(new_n496), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n491), .A2(new_n494), .A3(KEYINPUT68), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n483), .B(new_n485), .C1(new_n498), .C2(new_n495), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT83), .ZN(new_n501));
  NAND2_X1  g300(.A1(G228gat), .A2(G233gat), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT29), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n503), .B1(new_n432), .B2(new_n439), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n306), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n502), .B1(new_n505), .B2(new_n316), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n309), .A2(new_n503), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT81), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT81), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n309), .A2(new_n509), .A3(new_n503), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n508), .A2(new_n440), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n430), .A2(new_n431), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n437), .A2(new_n433), .A3(new_n438), .ZN(new_n514));
  AOI21_X1  g313(.A(KEYINPUT29), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n305), .A2(KEYINPUT79), .A3(new_n308), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT79), .B1(new_n305), .B2(new_n308), .ZN(new_n517));
  OAI22_X1  g316(.A1(new_n515), .A2(KEYINPUT3), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n507), .A2(new_n440), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(new_n502), .ZN(new_n521));
  INV_X1    g320(.A(G22gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n512), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT82), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G78gat), .B(G106gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(KEYINPUT31), .B(G50gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n501), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n528), .ZN(new_n530));
  AOI211_X1 g329(.A(KEYINPUT83), .B(new_n530), .C1(new_n523), .C2(new_n524), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n512), .A2(new_n521), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(G22gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(new_n523), .ZN(new_n534));
  NOR3_X1   g333(.A1(new_n529), .A2(new_n531), .A3(new_n534), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n533), .A2(new_n523), .ZN(new_n536));
  AOI22_X1  g335(.A1(new_n511), .A2(new_n506), .B1(new_n520), .B2(new_n502), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT82), .B1(new_n537), .B2(new_n522), .ZN(new_n538));
  OAI21_X1  g337(.A(KEYINPUT83), .B1(new_n538), .B2(new_n530), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n525), .A2(new_n501), .A3(new_n528), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n536), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n500), .B1(new_n535), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n265), .B1(new_n467), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n497), .A2(new_n499), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n534), .B1(new_n529), .B2(new_n531), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n539), .A2(new_n536), .A3(new_n540), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n464), .B1(new_n361), .B2(new_n367), .ZN(new_n548));
  INV_X1    g347(.A(new_n265), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n547), .A2(new_n548), .A3(new_n549), .A4(new_n466), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n543), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n544), .A2(KEYINPUT36), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT36), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n497), .A2(new_n499), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n545), .A2(new_n546), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n368), .A2(new_n465), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n555), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT37), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n441), .A2(new_n560), .A3(new_n452), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n462), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n560), .B1(new_n441), .B2(new_n452), .ZN(new_n563));
  OAI21_X1  g362(.A(KEYINPUT38), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n457), .ZN(new_n565));
  AND2_X1   g364(.A1(new_n561), .A2(new_n462), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n503), .B1(new_n407), .B2(new_n408), .ZN(new_n567));
  AOI22_X1  g366(.A1(new_n567), .A2(new_n369), .B1(new_n443), .B2(new_n446), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n560), .B1(new_n568), .B2(new_n440), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n417), .A2(new_n442), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT38), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n565), .B1(new_n566), .B2(new_n571), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n361), .A2(new_n367), .A3(new_n564), .A4(new_n572), .ZN(new_n573));
  AOI22_X1  g372(.A1(new_n362), .A2(new_n363), .B1(new_n332), .B2(new_n335), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n464), .B1(new_n574), .B2(new_n357), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n331), .A2(new_n322), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n333), .B1(new_n338), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n344), .A2(new_n333), .A3(new_n321), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(KEYINPUT39), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT85), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n578), .A2(KEYINPUT85), .A3(KEYINPUT39), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n357), .B1(new_n577), .B2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(KEYINPUT84), .B(KEYINPUT39), .ZN(new_n585));
  NOR3_X1   g384(.A1(new_n332), .A2(new_n333), .A3(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(KEYINPUT86), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT40), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI211_X1 g388(.A(KEYINPUT86), .B(KEYINPUT40), .C1(new_n584), .C2(new_n586), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n575), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  OAI211_X1 g390(.A(new_n556), .B(new_n573), .C1(new_n591), .C2(KEYINPUT87), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n589), .A2(new_n590), .ZN(new_n593));
  INV_X1    g392(.A(new_n575), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n593), .A2(KEYINPUT87), .A3(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n559), .B1(new_n592), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n263), .B1(new_n551), .B2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G57gat), .B(G64gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(G71gat), .A2(G78gat), .ZN(new_n600));
  INV_X1    g399(.A(G71gat), .ZN(new_n601));
  INV_X1    g400(.A(G78gat), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n601), .A2(new_n602), .A3(KEYINPUT9), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n599), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(G57gat), .B(G64gat), .Z(new_n605));
  INV_X1    g404(.A(KEYINPUT96), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT9), .ZN(new_n607));
  AOI22_X1  g406(.A1(new_n605), .A2(new_n606), .B1(new_n607), .B2(new_n600), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n599), .A2(KEYINPUT96), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n600), .A2(KEYINPUT95), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n600), .A2(KEYINPUT95), .ZN(new_n612));
  AOI22_X1  g411(.A1(new_n611), .A2(new_n612), .B1(new_n601), .B2(new_n602), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n604), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT97), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI211_X1 g415(.A(KEYINPUT97), .B(new_n604), .C1(new_n610), .C2(new_n613), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OR2_X1    g417(.A1(new_n618), .A2(KEYINPUT21), .ZN(new_n619));
  XNOR2_X1  g418(.A(G127gat), .B(G155gat), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n618), .A2(KEYINPUT21), .ZN(new_n624));
  INV_X1    g423(.A(new_n211), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n391), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AOI211_X1 g425(.A(G183gat), .B(new_n211), .C1(new_n618), .C2(KEYINPUT21), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n621), .B(new_n622), .C1(new_n626), .C2(new_n627), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT98), .ZN(new_n633));
  NAND2_X1  g432(.A1(G231gat), .A2(G233gat), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n633), .B(new_n634), .Z(new_n635));
  XOR2_X1   g434(.A(KEYINPUT99), .B(G211gat), .Z(new_n636));
  XOR2_X1   g435(.A(new_n635), .B(new_n636), .Z(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n631), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n629), .A2(new_n630), .A3(new_n637), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G134gat), .B(G162gat), .ZN(new_n643));
  NAND2_X1  g442(.A1(G232gat), .A2(G233gat), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT41), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n643), .B(new_n646), .Z(new_n647));
  XNOR2_X1  g446(.A(G190gat), .B(G218gat), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  OAI22_X1  g448(.A1(new_n649), .A2(KEYINPUT105), .B1(new_n645), .B2(new_n644), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT100), .ZN(new_n651));
  OAI211_X1 g450(.A(new_n651), .B(KEYINPUT7), .C1(new_n356), .C2(new_n455), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT7), .ZN(new_n653));
  OAI211_X1 g452(.A(G85gat), .B(G92gat), .C1(new_n653), .C2(KEYINPUT100), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(G99gat), .A2(G106gat), .ZN(new_n656));
  AOI22_X1  g455(.A1(KEYINPUT8), .A2(new_n656), .B1(new_n356), .B2(new_n455), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT101), .ZN(new_n659));
  XOR2_X1   g458(.A(G99gat), .B(G106gat), .Z(new_n660));
  OR3_X1    g459(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n659), .B1(new_n658), .B2(new_n660), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n658), .A2(new_n660), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT102), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n658), .A2(KEYINPUT102), .A3(new_n660), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n663), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(KEYINPUT103), .ZN(new_n670));
  AOI22_X1  g469(.A1(new_n662), .A2(new_n661), .B1(new_n666), .B2(new_n667), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT103), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n650), .B1(new_n675), .B2(new_n230), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT104), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n232), .A2(new_n233), .ZN(new_n678));
  AND3_X1   g477(.A1(new_n674), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n677), .B1(new_n674), .B2(new_n678), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n676), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n649), .A2(KEYINPUT105), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n676), .B(new_n682), .C1(new_n679), .C2(new_n680), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n647), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n684), .A2(new_n647), .A3(new_n685), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n663), .A2(new_n614), .A3(new_n664), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT10), .ZN(new_n691));
  OAI211_X1 g490(.A(new_n690), .B(new_n691), .C1(new_n618), .C2(new_n671), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n670), .A2(new_n618), .A3(new_n673), .A4(KEYINPUT10), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(G230gat), .A2(G233gat), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n690), .B1(new_n618), .B2(new_n671), .ZN(new_n697));
  INV_X1    g496(.A(new_n695), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(G120gat), .B(G148gat), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(G176gat), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(new_n418), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n696), .A2(new_n699), .A3(new_n703), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n642), .A2(new_n689), .A3(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n709), .A2(KEYINPUT106), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT106), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n684), .A2(new_n647), .A3(new_n685), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(new_n686), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n713), .A2(new_n641), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n711), .B1(new_n714), .B2(new_n708), .ZN(new_n715));
  OR2_X1    g514(.A1(new_n710), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n598), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n368), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g520(.A1(new_n718), .A2(new_n464), .ZN(new_n722));
  XNOR2_X1  g521(.A(KEYINPUT16), .B(G8gat), .ZN(new_n723));
  OR2_X1    g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT42), .ZN(new_n725));
  OR2_X1    g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n722), .A2(G8gat), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n724), .A2(new_n725), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(G1325gat));
  INV_X1    g528(.A(G15gat), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n718), .A2(new_n730), .A3(new_n500), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n717), .B1(new_n552), .B2(new_n554), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n731), .B1(new_n732), .B2(new_n730), .ZN(G1326gat));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n556), .ZN(new_n734));
  XOR2_X1   g533(.A(KEYINPUT43), .B(G22gat), .Z(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1327gat));
  OAI211_X1 g535(.A(new_n552), .B(new_n554), .C1(new_n548), .C2(new_n556), .ZN(new_n737));
  AOI21_X1  g536(.A(KEYINPUT87), .B1(new_n593), .B2(new_n594), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n573), .A2(new_n556), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n737), .B1(new_n740), .B2(new_n595), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n543), .A2(new_n550), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n713), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(KEYINPUT44), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n551), .A2(new_n597), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT44), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n745), .A2(new_n746), .A3(new_n713), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n642), .A2(new_n707), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n750), .A2(new_n263), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(G29gat), .B1(new_n753), .B2(new_n368), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n750), .A2(new_n689), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n598), .A2(new_n755), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n756), .A2(G29gat), .A3(new_n368), .ZN(new_n757));
  XNOR2_X1  g556(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n754), .A2(new_n759), .ZN(G1328gat));
  OAI21_X1  g559(.A(G36gat), .B1(new_n753), .B2(new_n465), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n756), .A2(G36gat), .A3(new_n465), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT46), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(G1329gat));
  NAND3_X1  g563(.A1(new_n752), .A2(G43gat), .A3(new_n555), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT108), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n598), .A2(new_n500), .A3(new_n755), .ZN(new_n767));
  INV_X1    g566(.A(G43gat), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  AND3_X1   g568(.A1(new_n765), .A2(KEYINPUT47), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT47), .B1(new_n765), .B2(new_n769), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n770), .A2(new_n771), .ZN(G1330gat));
  INV_X1    g571(.A(G50gat), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n773), .B1(new_n752), .B2(new_n557), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n598), .A2(new_n773), .A3(new_n557), .A4(new_n755), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT110), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  XOR2_X1   g576(.A(KEYINPUT109), .B(KEYINPUT48), .Z(new_n778));
  NAND2_X1  g577(.A1(new_n775), .A2(KEYINPUT48), .ZN(new_n779));
  OAI22_X1  g578(.A1(new_n777), .A2(new_n778), .B1(new_n774), .B2(new_n779), .ZN(G1331gat));
  NAND3_X1  g579(.A1(new_n714), .A2(new_n263), .A3(new_n707), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n781), .B1(new_n551), .B2(new_n597), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n719), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g583(.A(new_n464), .B(KEYINPUT111), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n786), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n782), .A2(new_n787), .ZN(new_n788));
  XOR2_X1   g587(.A(new_n788), .B(KEYINPUT112), .Z(new_n789));
  NOR2_X1   g588(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n789), .B(new_n790), .ZN(G1333gat));
  NAND2_X1  g590(.A1(new_n782), .A2(new_n500), .ZN(new_n792));
  AOI21_X1  g591(.A(G71gat), .B1(new_n792), .B2(KEYINPUT113), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n793), .B1(KEYINPUT113), .B2(new_n792), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n782), .A2(G71gat), .A3(new_n555), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n557), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g598(.A1(new_n642), .A2(new_n262), .A3(new_n708), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n748), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(G85gat), .B1(new_n801), .B2(new_n368), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n803), .B(new_n713), .C1(new_n741), .C2(new_n742), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n642), .A2(new_n262), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n803), .B1(new_n745), .B2(new_n713), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT51), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n743), .A2(KEYINPUT114), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n809), .A2(new_n810), .A3(new_n805), .A4(new_n804), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n808), .A2(new_n707), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n719), .A2(new_n356), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n802), .B1(new_n812), .B2(new_n813), .ZN(G1336gat));
  OAI21_X1  g613(.A(G92gat), .B1(new_n801), .B2(new_n786), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n786), .A2(G92gat), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n808), .A2(new_n811), .A3(new_n707), .A4(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n815), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(G92gat), .B1(new_n801), .B2(new_n465), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n820), .A2(new_n818), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n819), .B1(new_n821), .B2(new_n816), .ZN(G1337gat));
  INV_X1    g621(.A(G99gat), .ZN(new_n823));
  AOI211_X1 g622(.A(new_n823), .B(new_n801), .C1(new_n552), .C2(new_n554), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n812), .A2(new_n544), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n824), .B1(new_n823), .B2(new_n825), .ZN(G1338gat));
  AOI21_X1  g625(.A(new_n746), .B1(new_n745), .B2(new_n713), .ZN(new_n827));
  AOI211_X1 g626(.A(KEYINPUT44), .B(new_n689), .C1(new_n551), .C2(new_n597), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n557), .B(new_n800), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(G106gat), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT53), .B1(new_n830), .B2(KEYINPUT115), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n556), .A2(G106gat), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n808), .A2(new_n811), .A3(new_n707), .A4(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n830), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n833), .B(new_n830), .C1(KEYINPUT115), .C2(KEYINPUT53), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n835), .A2(new_n836), .ZN(G1339gat));
  NAND3_X1  g636(.A1(new_n692), .A2(new_n693), .A3(new_n698), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n696), .A2(KEYINPUT54), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n698), .B1(new_n692), .B2(new_n693), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n703), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n839), .A2(KEYINPUT55), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n706), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(KEYINPUT116), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n843), .A2(new_n846), .A3(new_n706), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n839), .A2(new_n842), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT55), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n845), .A2(new_n262), .A3(new_n847), .A4(new_n850), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n245), .A2(new_n246), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n237), .B1(new_n243), .B2(new_n236), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n255), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n261), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n707), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n713), .B1(new_n851), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n845), .A2(new_n847), .A3(new_n850), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n687), .A2(new_n856), .A3(new_n688), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n641), .B1(new_n858), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n709), .A2(new_n262), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n557), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n785), .A2(new_n368), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n865), .A2(new_n500), .A3(new_n866), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n867), .A2(new_n267), .A3(new_n263), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n368), .B1(new_n862), .B2(new_n864), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n869), .A2(new_n547), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n870), .A2(new_n786), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n262), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n868), .B1(new_n872), .B2(new_n267), .ZN(G1340gat));
  NAND2_X1  g672(.A1(new_n707), .A2(G120gat), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n867), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n869), .A2(new_n547), .A3(new_n707), .A4(new_n786), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n875), .B1(new_n268), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT117), .ZN(G1341gat));
  NAND3_X1  g677(.A1(new_n871), .A2(new_n271), .A3(new_n642), .ZN(new_n879));
  OAI21_X1  g678(.A(G127gat), .B1(new_n867), .B2(new_n641), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(G1342gat));
  NOR2_X1   g680(.A1(new_n689), .A2(new_n464), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT118), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT56), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n870), .A2(new_n280), .A3(new_n882), .A4(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n883), .A2(KEYINPUT56), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n885), .B(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(G134gat), .B1(new_n867), .B2(new_n689), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(KEYINPUT119), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(new_n889), .ZN(G1343gat));
  NOR2_X1   g689(.A1(new_n555), .A2(new_n556), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(KEYINPUT121), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n263), .A2(G141gat), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n869), .A2(new_n786), .A3(new_n892), .A4(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT58), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n894), .B1(KEYINPUT122), .B2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(new_n866), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n897), .A2(new_n555), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n557), .A2(KEYINPUT57), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n262), .A2(new_n850), .A3(new_n706), .A4(new_n843), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n713), .B1(new_n900), .B2(new_n857), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n641), .B1(new_n861), .B2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT120), .ZN(new_n903));
  OR2_X1    g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n863), .B1(new_n902), .B2(new_n903), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n899), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n862), .A2(new_n864), .ZN(new_n907));
  AOI21_X1  g706(.A(KEYINPUT57), .B1(new_n907), .B2(new_n557), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n262), .B(new_n898), .C1(new_n906), .C2(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n896), .B1(new_n909), .B2(G141gat), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n895), .A2(KEYINPUT122), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n910), .B(new_n911), .ZN(G1344gat));
  INV_X1    g711(.A(KEYINPUT57), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n913), .B1(new_n907), .B2(new_n557), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n557), .A2(new_n913), .ZN(new_n915));
  OAI21_X1  g714(.A(KEYINPUT124), .B1(new_n861), .B2(new_n901), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n917));
  AOI22_X1  g716(.A1(new_n844), .A2(KEYINPUT116), .B1(new_n849), .B2(new_n848), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n918), .A2(new_n713), .A3(new_n856), .A4(new_n847), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n900), .A2(new_n857), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n917), .B(new_n919), .C1(new_n920), .C2(new_n713), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n916), .A2(new_n921), .A3(new_n641), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n263), .B1(new_n710), .B2(new_n715), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n915), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(new_n898), .ZN(new_n925));
  NOR4_X1   g724(.A1(new_n914), .A2(new_n924), .A3(new_n708), .A4(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(KEYINPUT59), .B1(new_n926), .B2(new_n292), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n707), .B(new_n898), .C1(new_n906), .C2(new_n908), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT123), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n292), .A2(KEYINPUT59), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n929), .B1(new_n928), .B2(new_n930), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n927), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n869), .A2(new_n892), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n934), .A2(new_n785), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(new_n292), .A3(new_n707), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n933), .A2(new_n936), .ZN(G1345gat));
  OAI21_X1  g736(.A(new_n898), .B1(new_n906), .B2(new_n908), .ZN(new_n938));
  OAI21_X1  g737(.A(G155gat), .B1(new_n938), .B2(new_n641), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n935), .A2(new_n298), .A3(new_n642), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(G1346gat));
  OAI22_X1  g740(.A1(new_n938), .A2(new_n689), .B1(new_n288), .B2(new_n287), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n287), .A2(new_n288), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n882), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n942), .B1(new_n934), .B2(new_n944), .ZN(G1347gat));
  AOI21_X1  g744(.A(new_n719), .B1(new_n862), .B2(new_n864), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n786), .A2(new_n542), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(G169gat), .B1(new_n949), .B2(new_n262), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT126), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n368), .A2(new_n464), .A3(new_n500), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT125), .ZN(new_n953));
  AND3_X1   g752(.A1(new_n865), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n951), .B1(new_n865), .B2(new_n953), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n262), .A2(G169gat), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n950), .B1(new_n956), .B2(new_n957), .ZN(G1348gat));
  INV_X1    g757(.A(G176gat), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n949), .A2(new_n959), .A3(new_n707), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n954), .A2(new_n955), .A3(new_n708), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n960), .B1(new_n961), .B2(new_n959), .ZN(G1349gat));
  NAND3_X1  g761(.A1(new_n949), .A2(new_n398), .A3(new_n642), .ZN(new_n963));
  NOR3_X1   g762(.A1(new_n954), .A2(new_n955), .A3(new_n641), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n963), .B1(new_n964), .B2(new_n391), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(KEYINPUT60), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT60), .ZN(new_n967));
  OAI211_X1 g766(.A(new_n963), .B(new_n967), .C1(new_n964), .C2(new_n391), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n966), .A2(new_n968), .ZN(G1350gat));
  NAND3_X1  g768(.A1(new_n949), .A2(new_n395), .A3(new_n713), .ZN(new_n970));
  XOR2_X1   g769(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n971));
  INV_X1    g770(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n713), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n972), .B1(new_n973), .B2(G190gat), .ZN(new_n974));
  AOI211_X1 g773(.A(new_n395), .B(new_n971), .C1(new_n956), .C2(new_n713), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n970), .B1(new_n974), .B2(new_n975), .ZN(G1351gat));
  NOR3_X1   g775(.A1(new_n786), .A2(new_n555), .A3(new_n556), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n946), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g777(.A(G197gat), .B1(new_n978), .B2(new_n262), .ZN(new_n979));
  NOR3_X1   g778(.A1(new_n555), .A2(new_n719), .A3(new_n465), .ZN(new_n980));
  INV_X1    g779(.A(new_n980), .ZN(new_n981));
  NOR3_X1   g780(.A1(new_n914), .A2(new_n924), .A3(new_n981), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n263), .A2(new_n420), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n979), .B1(new_n982), .B2(new_n983), .ZN(G1352gat));
  NAND3_X1  g783(.A1(new_n978), .A2(new_n418), .A3(new_n707), .ZN(new_n985));
  XOR2_X1   g784(.A(new_n985), .B(KEYINPUT62), .Z(new_n986));
  NOR4_X1   g785(.A1(new_n914), .A2(new_n924), .A3(new_n708), .A4(new_n981), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n986), .B1(new_n987), .B2(new_n418), .ZN(G1353gat));
  INV_X1    g787(.A(G211gat), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n978), .A2(new_n989), .A3(new_n642), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n982), .A2(new_n642), .ZN(new_n991));
  AND3_X1   g790(.A1(new_n991), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n992));
  AOI21_X1  g791(.A(KEYINPUT63), .B1(new_n991), .B2(G211gat), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n990), .B1(new_n992), .B2(new_n993), .ZN(G1354gat));
  AOI21_X1  g793(.A(G218gat), .B1(new_n978), .B2(new_n713), .ZN(new_n995));
  AND2_X1   g794(.A1(new_n713), .A2(G218gat), .ZN(new_n996));
  AOI21_X1  g795(.A(new_n995), .B1(new_n982), .B2(new_n996), .ZN(G1355gat));
endmodule


