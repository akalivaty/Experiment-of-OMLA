

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578;

  XNOR2_X2 U321 ( .A(KEYINPUT110), .B(n490), .ZN(n496) );
  XOR2_X1 U322 ( .A(n310), .B(n406), .Z(n524) );
  XNOR2_X1 U323 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U324 ( .A(n368), .B(n367), .ZN(n370) );
  XNOR2_X1 U325 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n392) );
  XNOR2_X1 U326 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U327 ( .A(n393), .B(n392), .ZN(n539) );
  XNOR2_X1 U328 ( .A(n378), .B(n377), .ZN(n387) );
  NOR2_X1 U329 ( .A1(n524), .A2(n450), .ZN(n558) );
  XOR2_X1 U330 ( .A(n568), .B(n379), .Z(n545) );
  XNOR2_X1 U331 ( .A(n452), .B(G176GAT), .ZN(n453) );
  XNOR2_X1 U332 ( .A(n454), .B(n453), .ZN(G1349GAT) );
  XOR2_X1 U333 ( .A(G176GAT), .B(KEYINPUT91), .Z(n290) );
  XNOR2_X1 U334 ( .A(KEYINPUT88), .B(KEYINPUT92), .ZN(n289) );
  XNOR2_X1 U335 ( .A(n290), .B(n289), .ZN(n294) );
  XOR2_X1 U336 ( .A(G183GAT), .B(KEYINPUT87), .Z(n292) );
  XNOR2_X1 U337 ( .A(G169GAT), .B(KEYINPUT20), .ZN(n291) );
  XNOR2_X1 U338 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U339 ( .A(n294), .B(n293), .Z(n306) );
  XNOR2_X1 U340 ( .A(G127GAT), .B(KEYINPUT86), .ZN(n295) );
  XNOR2_X1 U341 ( .A(n295), .B(KEYINPUT0), .ZN(n296) );
  XOR2_X1 U342 ( .A(n296), .B(KEYINPUT85), .Z(n298) );
  XNOR2_X1 U343 ( .A(G113GAT), .B(G134GAT), .ZN(n297) );
  XNOR2_X1 U344 ( .A(n298), .B(n297), .ZN(n432) );
  XOR2_X1 U345 ( .A(G120GAT), .B(G71GAT), .Z(n363) );
  XOR2_X1 U346 ( .A(G99GAT), .B(G190GAT), .Z(n300) );
  XNOR2_X1 U347 ( .A(G43GAT), .B(G15GAT), .ZN(n299) );
  XNOR2_X1 U348 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U349 ( .A(n363), .B(n301), .Z(n303) );
  NAND2_X1 U350 ( .A1(G227GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U351 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U352 ( .A(n432), .B(n304), .ZN(n305) );
  XNOR2_X1 U353 ( .A(n306), .B(n305), .ZN(n310) );
  XOR2_X1 U354 ( .A(KEYINPUT90), .B(KEYINPUT19), .Z(n308) );
  XNOR2_X1 U355 ( .A(KEYINPUT89), .B(KEYINPUT17), .ZN(n307) );
  XNOR2_X1 U356 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U357 ( .A(KEYINPUT18), .B(n309), .Z(n406) );
  XOR2_X1 U358 ( .A(G183GAT), .B(KEYINPUT78), .Z(n394) );
  XNOR2_X1 U359 ( .A(G15GAT), .B(G1GAT), .ZN(n311) );
  XNOR2_X1 U360 ( .A(n311), .B(KEYINPUT70), .ZN(n354) );
  XOR2_X1 U361 ( .A(n354), .B(KEYINPUT15), .Z(n313) );
  NAND2_X1 U362 ( .A1(G231GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U364 ( .A(n394), .B(n314), .Z(n317) );
  XOR2_X1 U365 ( .A(G22GAT), .B(G155GAT), .Z(n434) );
  XNOR2_X1 U366 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n315) );
  XNOR2_X1 U367 ( .A(n315), .B(KEYINPUT72), .ZN(n364) );
  XNOR2_X1 U368 ( .A(n434), .B(n364), .ZN(n316) );
  XNOR2_X1 U369 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U370 ( .A(G78GAT), .B(G211GAT), .Z(n319) );
  XNOR2_X1 U371 ( .A(G127GAT), .B(G71GAT), .ZN(n318) );
  XNOR2_X1 U372 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U373 ( .A(n321), .B(n320), .Z(n329) );
  XOR2_X1 U374 ( .A(KEYINPUT79), .B(KEYINPUT82), .Z(n323) );
  XNOR2_X1 U375 ( .A(KEYINPUT14), .B(KEYINPUT81), .ZN(n322) );
  XNOR2_X1 U376 ( .A(n323), .B(n322), .ZN(n327) );
  XOR2_X1 U377 ( .A(KEYINPUT80), .B(KEYINPUT12), .Z(n325) );
  XNOR2_X1 U378 ( .A(G8GAT), .B(G64GAT), .ZN(n324) );
  XNOR2_X1 U379 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U380 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U381 ( .A(n329), .B(n328), .Z(n571) );
  INV_X1 U382 ( .A(n571), .ZN(n549) );
  XOR2_X1 U383 ( .A(G36GAT), .B(G190GAT), .Z(n401) );
  XOR2_X1 U384 ( .A(KEYINPUT9), .B(G106GAT), .Z(n331) );
  XNOR2_X1 U385 ( .A(G134GAT), .B(G218GAT), .ZN(n330) );
  XNOR2_X1 U386 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U387 ( .A(n401), .B(n332), .Z(n336) );
  XOR2_X1 U388 ( .A(G50GAT), .B(G162GAT), .Z(n435) );
  XOR2_X1 U389 ( .A(G92GAT), .B(KEYINPUT73), .Z(n334) );
  XNOR2_X1 U390 ( .A(G99GAT), .B(G85GAT), .ZN(n333) );
  XNOR2_X1 U391 ( .A(n334), .B(n333), .ZN(n372) );
  XNOR2_X1 U392 ( .A(n435), .B(n372), .ZN(n335) );
  XNOR2_X1 U393 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U394 ( .A(KEYINPUT11), .B(KEYINPUT77), .Z(n338) );
  NAND2_X1 U395 ( .A1(G232GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U396 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U397 ( .A(n340), .B(n339), .Z(n345) );
  XOR2_X1 U398 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n342) );
  XNOR2_X1 U399 ( .A(G43GAT), .B(G29GAT), .ZN(n341) );
  XNOR2_X1 U400 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U401 ( .A(KEYINPUT69), .B(n343), .Z(n358) );
  XNOR2_X1 U402 ( .A(n358), .B(KEYINPUT10), .ZN(n344) );
  XOR2_X1 U403 ( .A(n345), .B(n344), .Z(n552) );
  INV_X1 U404 ( .A(n552), .ZN(n557) );
  XNOR2_X1 U405 ( .A(KEYINPUT119), .B(KEYINPUT46), .ZN(n381) );
  XOR2_X1 U406 ( .A(KEYINPUT29), .B(KEYINPUT66), .Z(n347) );
  XNOR2_X1 U407 ( .A(KEYINPUT68), .B(KEYINPUT67), .ZN(n346) );
  XNOR2_X1 U408 ( .A(n347), .B(n346), .ZN(n362) );
  XOR2_X1 U409 ( .A(G22GAT), .B(G197GAT), .Z(n349) );
  XNOR2_X1 U410 ( .A(G36GAT), .B(G50GAT), .ZN(n348) );
  XNOR2_X1 U411 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U412 ( .A(KEYINPUT71), .B(KEYINPUT30), .Z(n351) );
  XNOR2_X1 U413 ( .A(G141GAT), .B(G113GAT), .ZN(n350) );
  XNOR2_X1 U414 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U415 ( .A(n353), .B(n352), .Z(n360) );
  XOR2_X1 U416 ( .A(G169GAT), .B(G8GAT), .Z(n407) );
  XOR2_X1 U417 ( .A(n407), .B(n354), .Z(n356) );
  NAND2_X1 U418 ( .A1(G229GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U419 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U420 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U421 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U422 ( .A(n362), .B(n361), .ZN(n563) );
  INV_X1 U423 ( .A(n563), .ZN(n542) );
  XNOR2_X1 U424 ( .A(n364), .B(n363), .ZN(n368) );
  AND2_X1 U425 ( .A1(G230GAT), .A2(G233GAT), .ZN(n366) );
  INV_X1 U426 ( .A(KEYINPUT74), .ZN(n365) );
  XOR2_X1 U427 ( .A(G176GAT), .B(G64GAT), .Z(n400) );
  XNOR2_X1 U428 ( .A(G204GAT), .B(n400), .ZN(n369) );
  XNOR2_X1 U429 ( .A(n370), .B(n369), .ZN(n378) );
  XNOR2_X1 U430 ( .A(G106GAT), .B(G78GAT), .ZN(n371) );
  XNOR2_X1 U431 ( .A(n371), .B(G148GAT), .ZN(n439) );
  XOR2_X1 U432 ( .A(n439), .B(n372), .Z(n376) );
  XOR2_X1 U433 ( .A(KEYINPUT32), .B(KEYINPUT75), .Z(n374) );
  XNOR2_X1 U434 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n373) );
  XNOR2_X1 U435 ( .A(n374), .B(n373), .ZN(n375) );
  INV_X1 U436 ( .A(n387), .ZN(n568) );
  XNOR2_X1 U437 ( .A(KEYINPUT41), .B(KEYINPUT65), .ZN(n379) );
  NOR2_X1 U438 ( .A1(n542), .A2(n545), .ZN(n380) );
  XOR2_X1 U439 ( .A(n381), .B(n380), .Z(n382) );
  NOR2_X1 U440 ( .A1(n557), .A2(n382), .ZN(n383) );
  NAND2_X1 U441 ( .A1(n549), .A2(n383), .ZN(n384) );
  XNOR2_X1 U442 ( .A(n384), .B(KEYINPUT47), .ZN(n391) );
  XOR2_X1 U443 ( .A(n552), .B(KEYINPUT109), .Z(n385) );
  XNOR2_X1 U444 ( .A(n385), .B(KEYINPUT36), .ZN(n575) );
  NOR2_X1 U445 ( .A1(n575), .A2(n549), .ZN(n386) );
  XNOR2_X1 U446 ( .A(KEYINPUT45), .B(n386), .ZN(n388) );
  NAND2_X1 U447 ( .A1(n388), .A2(n387), .ZN(n389) );
  NOR2_X1 U448 ( .A1(n563), .A2(n389), .ZN(n390) );
  NOR2_X1 U449 ( .A1(n391), .A2(n390), .ZN(n393) );
  XOR2_X1 U450 ( .A(KEYINPUT101), .B(n394), .Z(n399) );
  XOR2_X1 U451 ( .A(G211GAT), .B(G218GAT), .Z(n396) );
  XNOR2_X1 U452 ( .A(KEYINPUT21), .B(G204GAT), .ZN(n395) );
  XNOR2_X1 U453 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U454 ( .A(G197GAT), .B(n397), .Z(n446) );
  XNOR2_X1 U455 ( .A(n446), .B(G92GAT), .ZN(n398) );
  XNOR2_X1 U456 ( .A(n399), .B(n398), .ZN(n405) );
  XOR2_X1 U457 ( .A(n401), .B(n400), .Z(n403) );
  NAND2_X1 U458 ( .A1(G226GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U459 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U460 ( .A(n405), .B(n404), .Z(n409) );
  XNOR2_X1 U461 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U462 ( .A(n409), .B(n408), .ZN(n517) );
  NOR2_X1 U463 ( .A1(n539), .A2(n517), .ZN(n410) );
  XNOR2_X1 U464 ( .A(n410), .B(KEYINPUT54), .ZN(n433) );
  XOR2_X1 U465 ( .A(G85GAT), .B(KEYINPUT6), .Z(n412) );
  XNOR2_X1 U466 ( .A(G162GAT), .B(KEYINPUT1), .ZN(n411) );
  XNOR2_X1 U467 ( .A(n412), .B(n411), .ZN(n428) );
  XOR2_X1 U468 ( .A(KEYINPUT97), .B(KEYINPUT100), .Z(n414) );
  XNOR2_X1 U469 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n413) );
  XNOR2_X1 U470 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U471 ( .A(G155GAT), .B(G148GAT), .Z(n416) );
  XNOR2_X1 U472 ( .A(G29GAT), .B(G120GAT), .ZN(n415) );
  XNOR2_X1 U473 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U474 ( .A(n418), .B(n417), .Z(n426) );
  XOR2_X1 U475 ( .A(KEYINPUT95), .B(KEYINPUT2), .Z(n420) );
  XNOR2_X1 U476 ( .A(KEYINPUT3), .B(KEYINPUT96), .ZN(n419) );
  XNOR2_X1 U477 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U478 ( .A(G141GAT), .B(n421), .Z(n447) );
  XOR2_X1 U479 ( .A(KEYINPUT4), .B(KEYINPUT99), .Z(n423) );
  XNOR2_X1 U480 ( .A(KEYINPUT98), .B(G57GAT), .ZN(n422) );
  XNOR2_X1 U481 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U482 ( .A(n447), .B(n424), .ZN(n425) );
  XNOR2_X1 U483 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U484 ( .A(n428), .B(n427), .Z(n430) );
  NAND2_X1 U485 ( .A1(G225GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U486 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U487 ( .A(n432), .B(n431), .ZN(n538) );
  NAND2_X1 U488 ( .A1(n433), .A2(n538), .ZN(n561) );
  XOR2_X1 U489 ( .A(KEYINPUT94), .B(KEYINPUT22), .Z(n437) );
  XNOR2_X1 U490 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U492 ( .A(n438), .B(KEYINPUT93), .Z(n444) );
  XOR2_X1 U493 ( .A(n439), .B(KEYINPUT24), .Z(n441) );
  NAND2_X1 U494 ( .A1(G228GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U495 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U496 ( .A(n442), .B(KEYINPUT23), .ZN(n443) );
  XNOR2_X1 U497 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U498 ( .A(n446), .B(n445), .ZN(n448) );
  XOR2_X1 U499 ( .A(n448), .B(n447), .Z(n462) );
  NOR2_X1 U500 ( .A1(n561), .A2(n462), .ZN(n449) );
  XNOR2_X1 U501 ( .A(n449), .B(KEYINPUT55), .ZN(n450) );
  INV_X1 U502 ( .A(n545), .ZN(n451) );
  NAND2_X1 U503 ( .A1(n558), .A2(n451), .ZN(n454) );
  XOR2_X1 U504 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n452) );
  NOR2_X1 U505 ( .A1(n568), .A2(n542), .ZN(n455) );
  XNOR2_X1 U506 ( .A(n455), .B(KEYINPUT76), .ZN(n488) );
  XNOR2_X1 U507 ( .A(n517), .B(KEYINPUT27), .ZN(n460) );
  INV_X1 U508 ( .A(n460), .ZN(n456) );
  XOR2_X1 U509 ( .A(KEYINPUT28), .B(n462), .Z(n520) );
  NAND2_X1 U510 ( .A1(n456), .A2(n520), .ZN(n457) );
  NOR2_X1 U511 ( .A1(n538), .A2(n457), .ZN(n526) );
  XNOR2_X1 U512 ( .A(KEYINPUT102), .B(n526), .ZN(n458) );
  NAND2_X1 U513 ( .A1(n458), .A2(n524), .ZN(n468) );
  NAND2_X1 U514 ( .A1(n462), .A2(n524), .ZN(n459) );
  XNOR2_X1 U515 ( .A(n459), .B(KEYINPUT26), .ZN(n562) );
  NOR2_X1 U516 ( .A1(n562), .A2(n460), .ZN(n541) );
  NOR2_X1 U517 ( .A1(n524), .A2(n517), .ZN(n461) );
  NOR2_X1 U518 ( .A1(n462), .A2(n461), .ZN(n463) );
  XOR2_X1 U519 ( .A(KEYINPUT25), .B(n463), .Z(n464) );
  NOR2_X1 U520 ( .A1(n541), .A2(n464), .ZN(n465) );
  XNOR2_X1 U521 ( .A(n465), .B(KEYINPUT103), .ZN(n466) );
  NAND2_X1 U522 ( .A1(n466), .A2(n538), .ZN(n467) );
  NAND2_X1 U523 ( .A1(n468), .A2(n467), .ZN(n485) );
  XNOR2_X1 U524 ( .A(KEYINPUT16), .B(KEYINPUT84), .ZN(n469) );
  XNOR2_X1 U525 ( .A(n469), .B(KEYINPUT83), .ZN(n471) );
  NOR2_X1 U526 ( .A1(n557), .A2(n549), .ZN(n470) );
  XOR2_X1 U527 ( .A(n471), .B(n470), .Z(n472) );
  NAND2_X1 U528 ( .A1(n485), .A2(n472), .ZN(n473) );
  XOR2_X1 U529 ( .A(KEYINPUT104), .B(n473), .Z(n499) );
  NAND2_X1 U530 ( .A1(n488), .A2(n499), .ZN(n483) );
  NOR2_X1 U531 ( .A1(n538), .A2(n483), .ZN(n475) );
  XNOR2_X1 U532 ( .A(KEYINPUT34), .B(KEYINPUT105), .ZN(n474) );
  XNOR2_X1 U533 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U534 ( .A(G1GAT), .B(n476), .ZN(G1324GAT) );
  NOR2_X1 U535 ( .A1(n517), .A2(n483), .ZN(n478) );
  XNOR2_X1 U536 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n477) );
  XNOR2_X1 U537 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U538 ( .A(G8GAT), .B(n479), .ZN(G1325GAT) );
  NOR2_X1 U539 ( .A1(n524), .A2(n483), .ZN(n481) );
  XNOR2_X1 U540 ( .A(KEYINPUT35), .B(KEYINPUT108), .ZN(n480) );
  XNOR2_X1 U541 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U542 ( .A(G15GAT), .B(n482), .ZN(G1326GAT) );
  NOR2_X1 U543 ( .A1(n520), .A2(n483), .ZN(n484) );
  XOR2_X1 U544 ( .A(G22GAT), .B(n484), .Z(G1327GAT) );
  NOR2_X1 U545 ( .A1(n575), .A2(n571), .ZN(n486) );
  NAND2_X1 U546 ( .A1(n486), .A2(n485), .ZN(n487) );
  XNOR2_X1 U547 ( .A(KEYINPUT37), .B(n487), .ZN(n511) );
  NAND2_X1 U548 ( .A1(n488), .A2(n511), .ZN(n489) );
  XNOR2_X1 U549 ( .A(n489), .B(KEYINPUT38), .ZN(n490) );
  NOR2_X1 U550 ( .A1(n538), .A2(n496), .ZN(n492) );
  XNOR2_X1 U551 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n492), .B(n491), .ZN(G1328GAT) );
  NOR2_X1 U553 ( .A1(n517), .A2(n496), .ZN(n493) );
  XOR2_X1 U554 ( .A(G36GAT), .B(n493), .Z(G1329GAT) );
  NOR2_X1 U555 ( .A1(n524), .A2(n496), .ZN(n494) );
  XOR2_X1 U556 ( .A(KEYINPUT40), .B(n494), .Z(n495) );
  XNOR2_X1 U557 ( .A(G43GAT), .B(n495), .ZN(G1330GAT) );
  NOR2_X1 U558 ( .A1(n520), .A2(n496), .ZN(n498) );
  XNOR2_X1 U559 ( .A(G50GAT), .B(KEYINPUT111), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(G1331GAT) );
  NOR2_X1 U561 ( .A1(n545), .A2(n563), .ZN(n512) );
  NAND2_X1 U562 ( .A1(n499), .A2(n512), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n500), .B(KEYINPUT112), .ZN(n508) );
  NOR2_X1 U564 ( .A1(n508), .A2(n538), .ZN(n501) );
  XOR2_X1 U565 ( .A(KEYINPUT42), .B(n501), .Z(n502) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(n502), .ZN(G1332GAT) );
  XNOR2_X1 U567 ( .A(G64GAT), .B(KEYINPUT113), .ZN(n504) );
  NOR2_X1 U568 ( .A1(n517), .A2(n508), .ZN(n503) );
  XNOR2_X1 U569 ( .A(n504), .B(n503), .ZN(G1333GAT) );
  XNOR2_X1 U570 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n506) );
  NOR2_X1 U571 ( .A1(n524), .A2(n508), .ZN(n505) );
  XNOR2_X1 U572 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U573 ( .A(G71GAT), .B(n507), .ZN(G1334GAT) );
  NOR2_X1 U574 ( .A1(n508), .A2(n520), .ZN(n510) );
  XNOR2_X1 U575 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(G1335GAT) );
  NAND2_X1 U577 ( .A1(n512), .A2(n511), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n513), .B(KEYINPUT116), .ZN(n521) );
  NOR2_X1 U579 ( .A1(n521), .A2(n538), .ZN(n515) );
  XNOR2_X1 U580 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U582 ( .A(G85GAT), .B(n516), .ZN(G1336GAT) );
  NOR2_X1 U583 ( .A1(n517), .A2(n521), .ZN(n518) );
  XOR2_X1 U584 ( .A(G92GAT), .B(n518), .Z(G1337GAT) );
  NOR2_X1 U585 ( .A1(n524), .A2(n521), .ZN(n519) );
  XOR2_X1 U586 ( .A(G99GAT), .B(n519), .Z(G1338GAT) );
  NOR2_X1 U587 ( .A1(n521), .A2(n520), .ZN(n522) );
  XOR2_X1 U588 ( .A(KEYINPUT44), .B(n522), .Z(n523) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n523), .ZN(G1339GAT) );
  NOR2_X1 U590 ( .A1(n524), .A2(n539), .ZN(n525) );
  NAND2_X1 U591 ( .A1(n526), .A2(n525), .ZN(n535) );
  NOR2_X1 U592 ( .A1(n542), .A2(n535), .ZN(n527) );
  XOR2_X1 U593 ( .A(G113GAT), .B(n527), .Z(G1340GAT) );
  NOR2_X1 U594 ( .A1(n535), .A2(n545), .ZN(n531) );
  XOR2_X1 U595 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n529) );
  XNOR2_X1 U596 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n528) );
  XNOR2_X1 U597 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U598 ( .A(n531), .B(n530), .ZN(G1341GAT) );
  NOR2_X1 U599 ( .A1(n549), .A2(n535), .ZN(n533) );
  XNOR2_X1 U600 ( .A(KEYINPUT122), .B(KEYINPUT50), .ZN(n532) );
  XNOR2_X1 U601 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U602 ( .A(G127GAT), .B(n534), .Z(G1342GAT) );
  NOR2_X1 U603 ( .A1(n552), .A2(n535), .ZN(n537) );
  XNOR2_X1 U604 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n536) );
  XNOR2_X1 U605 ( .A(n537), .B(n536), .ZN(G1343GAT) );
  NOR2_X1 U606 ( .A1(n539), .A2(n538), .ZN(n540) );
  NAND2_X1 U607 ( .A1(n541), .A2(n540), .ZN(n551) );
  NOR2_X1 U608 ( .A1(n542), .A2(n551), .ZN(n544) );
  XNOR2_X1 U609 ( .A(G141GAT), .B(KEYINPUT123), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(G1344GAT) );
  NOR2_X1 U611 ( .A1(n545), .A2(n551), .ZN(n547) );
  XNOR2_X1 U612 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(n548), .ZN(G1345GAT) );
  NOR2_X1 U615 ( .A1(n549), .A2(n551), .ZN(n550) );
  XOR2_X1 U616 ( .A(G155GAT), .B(n550), .Z(G1346GAT) );
  NOR2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U618 ( .A(KEYINPUT124), .B(n553), .Z(n554) );
  XNOR2_X1 U619 ( .A(G162GAT), .B(n554), .ZN(G1347GAT) );
  NAND2_X1 U620 ( .A1(n563), .A2(n558), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n555), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U622 ( .A1(n571), .A2(n558), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(KEYINPUT58), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G190GAT), .B(n560), .ZN(G1351GAT) );
  XOR2_X1 U627 ( .A(G197GAT), .B(KEYINPUT59), .Z(n565) );
  NOR2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n573) );
  NAND2_X1 U629 ( .A1(n573), .A2(n563), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(n567) );
  XOR2_X1 U631 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(G1352GAT) );
  XOR2_X1 U633 ( .A(G204GAT), .B(KEYINPUT61), .Z(n570) );
  NAND2_X1 U634 ( .A1(n573), .A2(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1353GAT) );
  NAND2_X1 U636 ( .A1(n571), .A2(n573), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n572), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U638 ( .A(n573), .ZN(n574) );
  NOR2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n577) );
  XNOR2_X1 U640 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n577), .B(n576), .ZN(n578) );
  XOR2_X1 U642 ( .A(G218GAT), .B(n578), .Z(G1355GAT) );
endmodule

