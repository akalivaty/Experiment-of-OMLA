

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XNOR2_X1 U322 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U323 ( .A(KEYINPUT45), .B(KEYINPUT112), .ZN(n364) );
  XNOR2_X1 U324 ( .A(n365), .B(n364), .ZN(n367) );
  XNOR2_X1 U325 ( .A(n376), .B(n298), .ZN(n299) );
  XNOR2_X1 U326 ( .A(n418), .B(n299), .ZN(n300) );
  XNOR2_X1 U327 ( .A(n427), .B(KEYINPUT120), .ZN(n428) );
  XNOR2_X1 U328 ( .A(n429), .B(n428), .ZN(n450) );
  XNOR2_X1 U329 ( .A(n312), .B(n311), .ZN(n362) );
  XNOR2_X1 U330 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U331 ( .A(n456), .B(n455), .ZN(G1351GAT) );
  XOR2_X1 U332 ( .A(KEYINPUT65), .B(KEYINPUT9), .Z(n291) );
  XNOR2_X1 U333 ( .A(KEYINPUT67), .B(KEYINPUT79), .ZN(n290) );
  XNOR2_X1 U334 ( .A(n291), .B(n290), .ZN(n292) );
  XNOR2_X1 U335 ( .A(KEYINPUT10), .B(n292), .ZN(n294) );
  AND2_X1 U336 ( .A1(G232GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U337 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U338 ( .A(KEYINPUT68), .B(n295), .Z(n302) );
  XOR2_X1 U339 ( .A(G162GAT), .B(KEYINPUT77), .Z(n297) );
  XNOR2_X1 U340 ( .A(G50GAT), .B(G218GAT), .ZN(n296) );
  XNOR2_X1 U341 ( .A(n297), .B(n296), .ZN(n418) );
  XOR2_X1 U342 ( .A(G36GAT), .B(G190GAT), .Z(n376) );
  XOR2_X1 U343 ( .A(KEYINPUT11), .B(KEYINPUT78), .Z(n298) );
  XNOR2_X1 U344 ( .A(n300), .B(G134GAT), .ZN(n301) );
  XNOR2_X1 U345 ( .A(n302), .B(n301), .ZN(n312) );
  XOR2_X1 U346 ( .A(KEYINPUT74), .B(G85GAT), .Z(n304) );
  XNOR2_X1 U347 ( .A(G99GAT), .B(G92GAT), .ZN(n303) );
  XNOR2_X1 U348 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U349 ( .A(G106GAT), .B(n305), .Z(n323) );
  INV_X1 U350 ( .A(n323), .ZN(n310) );
  XOR2_X1 U351 ( .A(KEYINPUT70), .B(KEYINPUT7), .Z(n307) );
  XNOR2_X1 U352 ( .A(G43GAT), .B(G29GAT), .ZN(n306) );
  XNOR2_X1 U353 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U354 ( .A(KEYINPUT8), .B(n308), .Z(n330) );
  INV_X1 U355 ( .A(n330), .ZN(n309) );
  XOR2_X1 U356 ( .A(KEYINPUT75), .B(KEYINPUT32), .Z(n318) );
  XNOR2_X1 U357 ( .A(G78GAT), .B(KEYINPUT73), .ZN(n313) );
  XNOR2_X1 U358 ( .A(n313), .B(G148GAT), .ZN(n423) );
  XOR2_X1 U359 ( .A(KEYINPUT72), .B(KEYINPUT33), .Z(n315) );
  XNOR2_X1 U360 ( .A(G204GAT), .B(KEYINPUT31), .ZN(n314) );
  XNOR2_X1 U361 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U362 ( .A(n423), .B(n316), .ZN(n317) );
  XNOR2_X1 U363 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U364 ( .A(KEYINPUT13), .B(G57GAT), .Z(n348) );
  XOR2_X1 U365 ( .A(G176GAT), .B(G64GAT), .Z(n379) );
  XOR2_X1 U366 ( .A(n348), .B(n379), .Z(n320) );
  NAND2_X1 U367 ( .A1(G230GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U368 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U369 ( .A(n322), .B(n321), .Z(n325) );
  XOR2_X1 U370 ( .A(G120GAT), .B(G71GAT), .Z(n433) );
  XNOR2_X1 U371 ( .A(n433), .B(n323), .ZN(n324) );
  XNOR2_X1 U372 ( .A(n325), .B(n324), .ZN(n575) );
  XNOR2_X1 U373 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n326) );
  XNOR2_X1 U374 ( .A(n575), .B(n326), .ZN(n550) );
  XOR2_X1 U375 ( .A(G15GAT), .B(G197GAT), .Z(n328) );
  XNOR2_X1 U376 ( .A(G141GAT), .B(G22GAT), .ZN(n327) );
  XNOR2_X1 U377 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U378 ( .A(n330), .B(n329), .ZN(n340) );
  XOR2_X1 U379 ( .A(KEYINPUT71), .B(KEYINPUT30), .Z(n332) );
  XNOR2_X1 U380 ( .A(KEYINPUT29), .B(KEYINPUT69), .ZN(n331) );
  XNOR2_X1 U381 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U382 ( .A(G50GAT), .B(G36GAT), .Z(n334) );
  XOR2_X1 U383 ( .A(G169GAT), .B(G8GAT), .Z(n385) );
  XOR2_X1 U384 ( .A(G113GAT), .B(G1GAT), .Z(n395) );
  XNOR2_X1 U385 ( .A(n385), .B(n395), .ZN(n333) );
  XNOR2_X1 U386 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U387 ( .A(n336), .B(n335), .Z(n338) );
  NAND2_X1 U388 ( .A1(G229GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U389 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U390 ( .A(n340), .B(n339), .ZN(n570) );
  INV_X1 U391 ( .A(n570), .ZN(n547) );
  NAND2_X1 U392 ( .A1(n550), .A2(n547), .ZN(n341) );
  XNOR2_X1 U393 ( .A(KEYINPUT46), .B(n341), .ZN(n359) );
  XOR2_X1 U394 ( .A(G64GAT), .B(G71GAT), .Z(n343) );
  XNOR2_X1 U395 ( .A(G8GAT), .B(G183GAT), .ZN(n342) );
  XNOR2_X1 U396 ( .A(n343), .B(n342), .ZN(n347) );
  XOR2_X1 U397 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n345) );
  XNOR2_X1 U398 ( .A(G1GAT), .B(KEYINPUT12), .ZN(n344) );
  XNOR2_X1 U399 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U400 ( .A(n347), .B(n346), .ZN(n358) );
  XOR2_X1 U401 ( .A(G22GAT), .B(G155GAT), .Z(n414) );
  XOR2_X1 U402 ( .A(n348), .B(n414), .Z(n350) );
  XNOR2_X1 U403 ( .A(G211GAT), .B(G78GAT), .ZN(n349) );
  XNOR2_X1 U404 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U405 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n352) );
  NAND2_X1 U406 ( .A1(G231GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U407 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U408 ( .A(n354), .B(n353), .Z(n356) );
  XOR2_X1 U409 ( .A(G15GAT), .B(G127GAT), .Z(n443) );
  XNOR2_X1 U410 ( .A(n443), .B(KEYINPUT81), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U412 ( .A(n358), .B(n357), .ZN(n578) );
  NAND2_X1 U413 ( .A1(n359), .A2(n578), .ZN(n360) );
  NOR2_X1 U414 ( .A1(n362), .A2(n360), .ZN(n361) );
  XNOR2_X1 U415 ( .A(KEYINPUT47), .B(n361), .ZN(n370) );
  XNOR2_X1 U416 ( .A(KEYINPUT36), .B(KEYINPUT99), .ZN(n363) );
  XNOR2_X1 U417 ( .A(KEYINPUT80), .B(n362), .ZN(n540) );
  XNOR2_X1 U418 ( .A(n363), .B(n540), .ZN(n484) );
  NOR2_X1 U419 ( .A1(n578), .A2(n484), .ZN(n365) );
  AND2_X1 U420 ( .A1(n575), .A2(n570), .ZN(n366) );
  AND2_X1 U421 ( .A1(n367), .A2(n366), .ZN(n368) );
  XNOR2_X1 U422 ( .A(n368), .B(KEYINPUT113), .ZN(n369) );
  NAND2_X1 U423 ( .A1(n370), .A2(n369), .ZN(n371) );
  XNOR2_X1 U424 ( .A(KEYINPUT48), .B(n371), .ZN(n529) );
  XOR2_X1 U425 ( .A(G183GAT), .B(KEYINPUT18), .Z(n373) );
  XNOR2_X1 U426 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n372) );
  XNOR2_X1 U427 ( .A(n373), .B(n372), .ZN(n442) );
  XNOR2_X1 U428 ( .A(n442), .B(G218GAT), .ZN(n374) );
  XNOR2_X1 U429 ( .A(n374), .B(G92GAT), .ZN(n375) );
  XOR2_X1 U430 ( .A(n376), .B(n375), .Z(n378) );
  NAND2_X1 U431 ( .A1(G226GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U432 ( .A(n378), .B(n377), .ZN(n380) );
  XOR2_X1 U433 ( .A(n380), .B(n379), .Z(n387) );
  XNOR2_X1 U434 ( .A(G211GAT), .B(KEYINPUT91), .ZN(n381) );
  XNOR2_X1 U435 ( .A(n381), .B(KEYINPUT92), .ZN(n382) );
  XOR2_X1 U436 ( .A(n382), .B(KEYINPUT21), .Z(n384) );
  XNOR2_X1 U437 ( .A(G197GAT), .B(G204GAT), .ZN(n383) );
  XNOR2_X1 U438 ( .A(n384), .B(n383), .ZN(n424) );
  XNOR2_X1 U439 ( .A(n385), .B(n424), .ZN(n386) );
  XNOR2_X1 U440 ( .A(n387), .B(n386), .ZN(n476) );
  NAND2_X1 U441 ( .A1(n529), .A2(n476), .ZN(n389) );
  XOR2_X1 U442 ( .A(KEYINPUT119), .B(KEYINPUT54), .Z(n388) );
  XNOR2_X1 U443 ( .A(n389), .B(n388), .ZN(n410) );
  XOR2_X1 U444 ( .A(KEYINPUT5), .B(KEYINPUT6), .Z(n391) );
  XNOR2_X1 U445 ( .A(G120GAT), .B(G57GAT), .ZN(n390) );
  XNOR2_X1 U446 ( .A(n391), .B(n390), .ZN(n399) );
  XOR2_X1 U447 ( .A(G155GAT), .B(G162GAT), .Z(n393) );
  XNOR2_X1 U448 ( .A(G127GAT), .B(G148GAT), .ZN(n392) );
  XNOR2_X1 U449 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U450 ( .A(n394), .B(G85GAT), .Z(n397) );
  XNOR2_X1 U451 ( .A(G29GAT), .B(n395), .ZN(n396) );
  XNOR2_X1 U452 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U453 ( .A(n399), .B(n398), .ZN(n409) );
  XOR2_X1 U454 ( .A(KEYINPUT1), .B(KEYINPUT94), .Z(n401) );
  NAND2_X1 U455 ( .A1(G225GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U456 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U457 ( .A(n402), .B(KEYINPUT4), .Z(n407) );
  XOR2_X1 U458 ( .A(KEYINPUT85), .B(KEYINPUT0), .Z(n404) );
  XNOR2_X1 U459 ( .A(G134GAT), .B(KEYINPUT84), .ZN(n403) );
  XNOR2_X1 U460 ( .A(n404), .B(n403), .ZN(n436) );
  XNOR2_X1 U461 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n405) );
  XNOR2_X1 U462 ( .A(n405), .B(KEYINPUT2), .ZN(n421) );
  XNOR2_X1 U463 ( .A(n436), .B(n421), .ZN(n406) );
  XNOR2_X1 U464 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U465 ( .A(n409), .B(n408), .ZN(n464) );
  NOR2_X1 U466 ( .A1(n410), .A2(n464), .ZN(n569) );
  XOR2_X1 U467 ( .A(KEYINPUT22), .B(KEYINPUT93), .Z(n412) );
  XNOR2_X1 U468 ( .A(G106GAT), .B(KEYINPUT23), .ZN(n411) );
  XNOR2_X1 U469 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U470 ( .A(n414), .B(n413), .Z(n416) );
  NAND2_X1 U471 ( .A1(G228GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U472 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U473 ( .A(n417), .B(KEYINPUT90), .Z(n420) );
  XNOR2_X1 U474 ( .A(n418), .B(KEYINPUT24), .ZN(n419) );
  XNOR2_X1 U475 ( .A(n420), .B(n419), .ZN(n422) );
  XOR2_X1 U476 ( .A(n422), .B(n421), .Z(n426) );
  XNOR2_X1 U477 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U478 ( .A(n426), .B(n425), .ZN(n466) );
  NAND2_X1 U479 ( .A1(n569), .A2(n466), .ZN(n429) );
  XOR2_X1 U480 ( .A(KEYINPUT121), .B(KEYINPUT55), .Z(n427) );
  XOR2_X1 U481 ( .A(KEYINPUT89), .B(KEYINPUT88), .Z(n431) );
  XNOR2_X1 U482 ( .A(G190GAT), .B(KEYINPUT86), .ZN(n430) );
  XNOR2_X1 U483 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U484 ( .A(n432), .B(G99GAT), .Z(n435) );
  XNOR2_X1 U485 ( .A(G43GAT), .B(n433), .ZN(n434) );
  XNOR2_X1 U486 ( .A(n435), .B(n434), .ZN(n437) );
  XOR2_X1 U487 ( .A(n437), .B(n436), .Z(n439) );
  XNOR2_X1 U488 ( .A(G169GAT), .B(G113GAT), .ZN(n438) );
  XNOR2_X1 U489 ( .A(n439), .B(n438), .ZN(n449) );
  XOR2_X1 U490 ( .A(G176GAT), .B(KEYINPUT20), .Z(n441) );
  XNOR2_X1 U491 ( .A(KEYINPUT66), .B(KEYINPUT87), .ZN(n440) );
  XNOR2_X1 U492 ( .A(n441), .B(n440), .ZN(n447) );
  XOR2_X1 U493 ( .A(n443), .B(n442), .Z(n445) );
  NAND2_X1 U494 ( .A1(G227GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U495 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U496 ( .A(n447), .B(n446), .Z(n448) );
  XNOR2_X1 U497 ( .A(n449), .B(n448), .ZN(n531) );
  NAND2_X1 U498 ( .A1(n450), .A2(n531), .ZN(n452) );
  INV_X1 U499 ( .A(KEYINPUT122), .ZN(n451) );
  XNOR2_X1 U500 ( .A(n452), .B(n451), .ZN(n559) );
  NAND2_X1 U501 ( .A1(n559), .A2(n540), .ZN(n456) );
  XOR2_X1 U502 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n454) );
  INV_X1 U503 ( .A(G190GAT), .ZN(n453) );
  INV_X1 U504 ( .A(n464), .ZN(n516) );
  NAND2_X1 U505 ( .A1(n476), .A2(n531), .ZN(n457) );
  XOR2_X1 U506 ( .A(KEYINPUT95), .B(n457), .Z(n458) );
  NAND2_X1 U507 ( .A1(n466), .A2(n458), .ZN(n459) );
  XNOR2_X1 U508 ( .A(n459), .B(KEYINPUT25), .ZN(n462) );
  NOR2_X1 U509 ( .A1(n531), .A2(n466), .ZN(n460) );
  XNOR2_X1 U510 ( .A(n460), .B(KEYINPUT26), .ZN(n568) );
  INV_X1 U511 ( .A(n568), .ZN(n544) );
  XOR2_X1 U512 ( .A(n476), .B(KEYINPUT27), .Z(n465) );
  NOR2_X1 U513 ( .A1(n544), .A2(n465), .ZN(n461) );
  NOR2_X1 U514 ( .A1(n462), .A2(n461), .ZN(n463) );
  NOR2_X1 U515 ( .A1(n464), .A2(n463), .ZN(n469) );
  NOR2_X1 U516 ( .A1(n465), .A2(n516), .ZN(n528) );
  XNOR2_X1 U517 ( .A(n466), .B(KEYINPUT28), .ZN(n530) );
  NAND2_X1 U518 ( .A1(n528), .A2(n530), .ZN(n467) );
  NOR2_X1 U519 ( .A1(n467), .A2(n531), .ZN(n468) );
  NOR2_X1 U520 ( .A1(n469), .A2(n468), .ZN(n485) );
  NOR2_X1 U521 ( .A1(n578), .A2(n540), .ZN(n470) );
  XOR2_X1 U522 ( .A(KEYINPUT16), .B(n470), .Z(n471) );
  NOR2_X1 U523 ( .A1(n485), .A2(n471), .ZN(n502) );
  NAND2_X1 U524 ( .A1(n547), .A2(n575), .ZN(n472) );
  XOR2_X1 U525 ( .A(KEYINPUT76), .B(n472), .Z(n489) );
  NAND2_X1 U526 ( .A1(n502), .A2(n489), .ZN(n481) );
  NOR2_X1 U527 ( .A1(n516), .A2(n481), .ZN(n474) );
  XNOR2_X1 U528 ( .A(KEYINPUT34), .B(KEYINPUT96), .ZN(n473) );
  XNOR2_X1 U529 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U530 ( .A(G1GAT), .B(n475), .Z(G1324GAT) );
  INV_X1 U531 ( .A(n476), .ZN(n519) );
  NOR2_X1 U532 ( .A1(n519), .A2(n481), .ZN(n477) );
  XOR2_X1 U533 ( .A(G8GAT), .B(n477), .Z(G1325GAT) );
  INV_X1 U534 ( .A(n531), .ZN(n522) );
  NOR2_X1 U535 ( .A1(n522), .A2(n481), .ZN(n479) );
  XNOR2_X1 U536 ( .A(KEYINPUT97), .B(KEYINPUT35), .ZN(n478) );
  XNOR2_X1 U537 ( .A(n479), .B(n478), .ZN(n480) );
  XOR2_X1 U538 ( .A(G15GAT), .B(n480), .Z(G1326GAT) );
  NOR2_X1 U539 ( .A1(n530), .A2(n481), .ZN(n482) );
  XOR2_X1 U540 ( .A(KEYINPUT98), .B(n482), .Z(n483) );
  XNOR2_X1 U541 ( .A(G22GAT), .B(n483), .ZN(G1327GAT) );
  NOR2_X1 U542 ( .A1(n484), .A2(n485), .ZN(n486) );
  NAND2_X1 U543 ( .A1(n578), .A2(n486), .ZN(n487) );
  XNOR2_X1 U544 ( .A(KEYINPUT37), .B(n487), .ZN(n488) );
  XNOR2_X1 U545 ( .A(KEYINPUT100), .B(n488), .ZN(n514) );
  NAND2_X1 U546 ( .A1(n514), .A2(n489), .ZN(n490) );
  XNOR2_X1 U547 ( .A(KEYINPUT38), .B(n490), .ZN(n499) );
  NOR2_X1 U548 ( .A1(n499), .A2(n516), .ZN(n493) );
  XOR2_X1 U549 ( .A(G29GAT), .B(KEYINPUT101), .Z(n491) );
  XNOR2_X1 U550 ( .A(KEYINPUT39), .B(n491), .ZN(n492) );
  XNOR2_X1 U551 ( .A(n493), .B(n492), .ZN(G1328GAT) );
  NOR2_X1 U552 ( .A1(n499), .A2(n519), .ZN(n494) );
  XOR2_X1 U553 ( .A(G36GAT), .B(n494), .Z(n495) );
  XNOR2_X1 U554 ( .A(KEYINPUT102), .B(n495), .ZN(G1329GAT) );
  XNOR2_X1 U555 ( .A(KEYINPUT40), .B(KEYINPUT103), .ZN(n497) );
  NOR2_X1 U556 ( .A1(n522), .A2(n499), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U558 ( .A(G43GAT), .B(n498), .ZN(G1330GAT) );
  NOR2_X1 U559 ( .A1(n499), .A2(n530), .ZN(n500) );
  XOR2_X1 U560 ( .A(KEYINPUT104), .B(n500), .Z(n501) );
  XNOR2_X1 U561 ( .A(G50GAT), .B(n501), .ZN(G1331GAT) );
  INV_X1 U562 ( .A(n550), .ZN(n561) );
  NOR2_X1 U563 ( .A1(n547), .A2(n561), .ZN(n515) );
  NAND2_X1 U564 ( .A1(n515), .A2(n502), .ZN(n510) );
  NOR2_X1 U565 ( .A1(n516), .A2(n510), .ZN(n504) );
  XNOR2_X1 U566 ( .A(KEYINPUT105), .B(KEYINPUT42), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(n505), .ZN(G1332GAT) );
  NOR2_X1 U569 ( .A1(n519), .A2(n510), .ZN(n507) );
  XNOR2_X1 U570 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U572 ( .A(G64GAT), .B(n508), .ZN(G1333GAT) );
  NOR2_X1 U573 ( .A1(n522), .A2(n510), .ZN(n509) );
  XOR2_X1 U574 ( .A(G71GAT), .B(n509), .Z(G1334GAT) );
  NOR2_X1 U575 ( .A1(n530), .A2(n510), .ZN(n512) );
  XNOR2_X1 U576 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U578 ( .A(G78GAT), .B(n513), .ZN(G1335GAT) );
  NAND2_X1 U579 ( .A1(n515), .A2(n514), .ZN(n524) );
  NOR2_X1 U580 ( .A1(n516), .A2(n524), .ZN(n518) );
  XNOR2_X1 U581 ( .A(G85GAT), .B(KEYINPUT109), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n518), .B(n517), .ZN(G1336GAT) );
  NOR2_X1 U583 ( .A1(n519), .A2(n524), .ZN(n520) );
  XOR2_X1 U584 ( .A(KEYINPUT110), .B(n520), .Z(n521) );
  XNOR2_X1 U585 ( .A(G92GAT), .B(n521), .ZN(G1337GAT) );
  NOR2_X1 U586 ( .A1(n522), .A2(n524), .ZN(n523) );
  XOR2_X1 U587 ( .A(G99GAT), .B(n523), .Z(G1338GAT) );
  NOR2_X1 U588 ( .A1(n530), .A2(n524), .ZN(n526) );
  XNOR2_X1 U589 ( .A(KEYINPUT44), .B(KEYINPUT111), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n527), .ZN(G1339GAT) );
  NAND2_X1 U592 ( .A1(n529), .A2(n528), .ZN(n545) );
  NAND2_X1 U593 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U594 ( .A1(n545), .A2(n532), .ZN(n533) );
  XNOR2_X1 U595 ( .A(KEYINPUT114), .B(n533), .ZN(n541) );
  NAND2_X1 U596 ( .A1(n541), .A2(n547), .ZN(n534) );
  XNOR2_X1 U597 ( .A(n534), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT49), .Z(n536) );
  NAND2_X1 U599 ( .A1(n550), .A2(n541), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n536), .B(n535), .ZN(G1341GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n538) );
  INV_X1 U602 ( .A(n578), .ZN(n555) );
  NAND2_X1 U603 ( .A1(n541), .A2(n555), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(n539), .ZN(G1342GAT) );
  XOR2_X1 U606 ( .A(G134GAT), .B(KEYINPUT51), .Z(n543) );
  NAND2_X1 U607 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(G1343GAT) );
  XOR2_X1 U609 ( .A(G141GAT), .B(KEYINPUT117), .Z(n549) );
  NOR2_X1 U610 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n546), .B(KEYINPUT116), .ZN(n557) );
  NAND2_X1 U612 ( .A1(n557), .A2(n547), .ZN(n548) );
  XNOR2_X1 U613 ( .A(n549), .B(n548), .ZN(G1344GAT) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n554) );
  XOR2_X1 U615 ( .A(KEYINPUT118), .B(KEYINPUT52), .Z(n552) );
  NAND2_X1 U616 ( .A1(n550), .A2(n557), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n554), .B(n553), .ZN(G1345GAT) );
  NAND2_X1 U619 ( .A1(n557), .A2(n555), .ZN(n556) );
  XNOR2_X1 U620 ( .A(n556), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U621 ( .A1(n557), .A2(n362), .ZN(n558) );
  XNOR2_X1 U622 ( .A(n558), .B(G162GAT), .ZN(G1347GAT) );
  INV_X1 U623 ( .A(n559), .ZN(n566) );
  NOR2_X1 U624 ( .A1(n566), .A2(n570), .ZN(n560) );
  XOR2_X1 U625 ( .A(n560), .B(G169GAT), .Z(G1348GAT) );
  NOR2_X1 U626 ( .A1(n561), .A2(n566), .ZN(n565) );
  XOR2_X1 U627 ( .A(KEYINPUT123), .B(KEYINPUT56), .Z(n563) );
  XNOR2_X1 U628 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(G1349GAT) );
  NOR2_X1 U631 ( .A1(n566), .A2(n578), .ZN(n567) );
  XOR2_X1 U632 ( .A(n567), .B(G183GAT), .Z(G1350GAT) );
  NAND2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n581) );
  NOR2_X1 U634 ( .A1(n581), .A2(n570), .ZN(n574) );
  XOR2_X1 U635 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n572) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  NOR2_X1 U639 ( .A1(n575), .A2(n581), .ZN(n577) );
  XNOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NOR2_X1 U642 ( .A1(n578), .A2(n581), .ZN(n579) );
  XOR2_X1 U643 ( .A(KEYINPUT126), .B(n579), .Z(n580) );
  XNOR2_X1 U644 ( .A(G211GAT), .B(n580), .ZN(G1354GAT) );
  NOR2_X1 U645 ( .A1(n484), .A2(n581), .ZN(n583) );
  XNOR2_X1 U646 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

