

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U553 ( .A1(G651), .A2(n564), .ZN(n794) );
  NOR2_X1 U554 ( .A1(n564), .A2(n532), .ZN(n788) );
  NOR2_X1 U555 ( .A1(G1384), .A2(G164), .ZN(n700) );
  OR2_X1 U556 ( .A1(n611), .A2(n986), .ZN(n614) );
  NOR2_X1 U557 ( .A1(n614), .A2(n613), .ZN(n625) );
  INV_X1 U558 ( .A(KEYINPUT100), .ZN(n623) );
  XNOR2_X1 U559 ( .A(n624), .B(n623), .ZN(n632) );
  NAND2_X1 U560 ( .A1(n598), .A2(n700), .ZN(n626) );
  INV_X1 U561 ( .A(KEYINPUT65), .ZN(n593) );
  INV_X1 U562 ( .A(G2104), .ZN(n525) );
  NOR2_X1 U563 ( .A1(G2105), .A2(n525), .ZN(n589) );
  BUF_X1 U564 ( .A(n589), .Z(n898) );
  NAND2_X1 U565 ( .A1(G102), .A2(n898), .ZN(n524) );
  NOR2_X1 U566 ( .A1(G2105), .A2(G2104), .ZN(n522) );
  XOR2_X2 U567 ( .A(KEYINPUT17), .B(n522), .Z(n895) );
  NAND2_X1 U568 ( .A1(G138), .A2(n895), .ZN(n523) );
  NAND2_X1 U569 ( .A1(n524), .A2(n523), .ZN(n530) );
  INV_X1 U570 ( .A(G2105), .ZN(n526) );
  NOR2_X1 U571 ( .A1(n526), .A2(n525), .ZN(n891) );
  NAND2_X1 U572 ( .A1(G114), .A2(n891), .ZN(n528) );
  NOR2_X2 U573 ( .A1(G2104), .A2(n526), .ZN(n889) );
  NAND2_X1 U574 ( .A1(G126), .A2(n889), .ZN(n527) );
  NAND2_X1 U575 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U576 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U577 ( .A(n531), .B(KEYINPUT92), .ZN(G164) );
  XOR2_X1 U578 ( .A(G543), .B(KEYINPUT0), .Z(n564) );
  INV_X1 U579 ( .A(G651), .ZN(n532) );
  NAND2_X1 U580 ( .A1(n788), .A2(G78), .ZN(n536) );
  NOR2_X1 U581 ( .A1(G543), .A2(n532), .ZN(n533) );
  XOR2_X1 U582 ( .A(KEYINPUT66), .B(n533), .Z(n534) );
  XNOR2_X1 U583 ( .A(KEYINPUT1), .B(n534), .ZN(n797) );
  NAND2_X1 U584 ( .A1(G65), .A2(n797), .ZN(n535) );
  NAND2_X1 U585 ( .A1(n536), .A2(n535), .ZN(n539) );
  NOR2_X1 U586 ( .A1(G651), .A2(G543), .ZN(n790) );
  NAND2_X1 U587 ( .A1(G91), .A2(n790), .ZN(n537) );
  XNOR2_X1 U588 ( .A(KEYINPUT67), .B(n537), .ZN(n538) );
  NOR2_X1 U589 ( .A1(n539), .A2(n538), .ZN(n541) );
  NAND2_X1 U590 ( .A1(n794), .A2(G53), .ZN(n540) );
  NAND2_X1 U591 ( .A1(n541), .A2(n540), .ZN(G299) );
  NAND2_X1 U592 ( .A1(n794), .A2(G52), .ZN(n543) );
  NAND2_X1 U593 ( .A1(G64), .A2(n797), .ZN(n542) );
  NAND2_X1 U594 ( .A1(n543), .A2(n542), .ZN(n548) );
  NAND2_X1 U595 ( .A1(G77), .A2(n788), .ZN(n545) );
  NAND2_X1 U596 ( .A1(G90), .A2(n790), .ZN(n544) );
  NAND2_X1 U597 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U598 ( .A(KEYINPUT9), .B(n546), .Z(n547) );
  NOR2_X1 U599 ( .A1(n548), .A2(n547), .ZN(G171) );
  NAND2_X1 U600 ( .A1(n790), .A2(G89), .ZN(n549) );
  XNOR2_X1 U601 ( .A(n549), .B(KEYINPUT4), .ZN(n551) );
  NAND2_X1 U602 ( .A1(G76), .A2(n788), .ZN(n550) );
  NAND2_X1 U603 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U604 ( .A(n552), .B(KEYINPUT5), .ZN(n557) );
  NAND2_X1 U605 ( .A1(n794), .A2(G51), .ZN(n554) );
  NAND2_X1 U606 ( .A1(G63), .A2(n797), .ZN(n553) );
  NAND2_X1 U607 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U608 ( .A(KEYINPUT6), .B(n555), .Z(n556) );
  NAND2_X1 U609 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U610 ( .A(n558), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U611 ( .A1(n794), .A2(G49), .ZN(n559) );
  XOR2_X1 U612 ( .A(KEYINPUT82), .B(n559), .Z(n560) );
  NOR2_X1 U613 ( .A1(n797), .A2(n560), .ZN(n562) );
  NAND2_X1 U614 ( .A1(G651), .A2(G74), .ZN(n561) );
  NAND2_X1 U615 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U616 ( .A(n563), .B(KEYINPUT83), .ZN(n566) );
  NAND2_X1 U617 ( .A1(G87), .A2(n564), .ZN(n565) );
  NAND2_X1 U618 ( .A1(n566), .A2(n565), .ZN(G288) );
  XOR2_X1 U619 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U620 ( .A1(G88), .A2(n790), .ZN(n567) );
  XNOR2_X1 U621 ( .A(n567), .B(KEYINPUT84), .ZN(n569) );
  NAND2_X1 U622 ( .A1(n788), .A2(G75), .ZN(n568) );
  NAND2_X1 U623 ( .A1(n569), .A2(n568), .ZN(n573) );
  NAND2_X1 U624 ( .A1(n794), .A2(G50), .ZN(n571) );
  NAND2_X1 U625 ( .A1(G62), .A2(n797), .ZN(n570) );
  NAND2_X1 U626 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U627 ( .A1(n573), .A2(n572), .ZN(G166) );
  XNOR2_X1 U628 ( .A(KEYINPUT93), .B(G166), .ZN(G303) );
  NAND2_X1 U629 ( .A1(n790), .A2(G86), .ZN(n575) );
  NAND2_X1 U630 ( .A1(G61), .A2(n797), .ZN(n574) );
  NAND2_X1 U631 ( .A1(n575), .A2(n574), .ZN(n578) );
  NAND2_X1 U632 ( .A1(n788), .A2(G73), .ZN(n576) );
  XOR2_X1 U633 ( .A(KEYINPUT2), .B(n576), .Z(n577) );
  NOR2_X1 U634 ( .A1(n578), .A2(n577), .ZN(n580) );
  NAND2_X1 U635 ( .A1(n794), .A2(G48), .ZN(n579) );
  NAND2_X1 U636 ( .A1(n580), .A2(n579), .ZN(G305) );
  AND2_X1 U637 ( .A1(G60), .A2(n797), .ZN(n584) );
  NAND2_X1 U638 ( .A1(G72), .A2(n788), .ZN(n582) );
  NAND2_X1 U639 ( .A1(G85), .A2(n790), .ZN(n581) );
  NAND2_X1 U640 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U641 ( .A1(n584), .A2(n583), .ZN(n586) );
  NAND2_X1 U642 ( .A1(n794), .A2(G47), .ZN(n585) );
  NAND2_X1 U643 ( .A1(n586), .A2(n585), .ZN(G290) );
  NAND2_X1 U644 ( .A1(G113), .A2(n891), .ZN(n588) );
  NAND2_X1 U645 ( .A1(G137), .A2(n895), .ZN(n587) );
  NAND2_X1 U646 ( .A1(n588), .A2(n587), .ZN(n596) );
  NAND2_X1 U647 ( .A1(n889), .A2(G125), .ZN(n592) );
  NAND2_X1 U648 ( .A1(n589), .A2(G101), .ZN(n590) );
  XOR2_X1 U649 ( .A(n590), .B(KEYINPUT23), .Z(n591) );
  NAND2_X1 U650 ( .A1(n592), .A2(n591), .ZN(n594) );
  XNOR2_X1 U651 ( .A(n594), .B(n593), .ZN(n595) );
  NOR2_X1 U652 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U653 ( .A(n597), .B(KEYINPUT64), .ZN(G160) );
  NAND2_X1 U654 ( .A1(G160), .A2(G40), .ZN(n699) );
  INV_X1 U655 ( .A(n699), .ZN(n598) );
  NOR2_X1 U656 ( .A1(G2084), .A2(n626), .ZN(n648) );
  NAND2_X1 U657 ( .A1(G8), .A2(n648), .ZN(n599) );
  XNOR2_X1 U658 ( .A(n599), .B(KEYINPUT98), .ZN(n658) );
  AND2_X1 U659 ( .A1(n626), .A2(G1341), .ZN(n611) );
  XOR2_X1 U660 ( .A(KEYINPUT70), .B(KEYINPUT14), .Z(n601) );
  NAND2_X1 U661 ( .A1(G56), .A2(n797), .ZN(n600) );
  XNOR2_X1 U662 ( .A(n601), .B(n600), .ZN(n608) );
  NAND2_X1 U663 ( .A1(n788), .A2(G68), .ZN(n602) );
  XNOR2_X1 U664 ( .A(KEYINPUT71), .B(n602), .ZN(n605) );
  NAND2_X1 U665 ( .A1(n790), .A2(G81), .ZN(n603) );
  XOR2_X1 U666 ( .A(KEYINPUT12), .B(n603), .Z(n604) );
  NOR2_X1 U667 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U668 ( .A(n606), .B(KEYINPUT13), .ZN(n607) );
  NOR2_X1 U669 ( .A1(n608), .A2(n607), .ZN(n610) );
  NAND2_X1 U670 ( .A1(n794), .A2(G43), .ZN(n609) );
  NAND2_X1 U671 ( .A1(n610), .A2(n609), .ZN(n986) );
  INV_X1 U672 ( .A(G1996), .ZN(n946) );
  NOR2_X1 U673 ( .A1(n626), .A2(n946), .ZN(n612) );
  XNOR2_X1 U674 ( .A(n612), .B(KEYINPUT26), .ZN(n613) );
  NAND2_X1 U675 ( .A1(G92), .A2(n790), .ZN(n621) );
  NAND2_X1 U676 ( .A1(n788), .A2(G79), .ZN(n616) );
  NAND2_X1 U677 ( .A1(G66), .A2(n797), .ZN(n615) );
  NAND2_X1 U678 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U679 ( .A1(n794), .A2(G54), .ZN(n617) );
  XOR2_X1 U680 ( .A(KEYINPUT72), .B(n617), .Z(n618) );
  NOR2_X1 U681 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U682 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U683 ( .A(n622), .B(KEYINPUT15), .ZN(n970) );
  NOR2_X1 U684 ( .A1(n625), .A2(n970), .ZN(n624) );
  NAND2_X1 U685 ( .A1(n625), .A2(n970), .ZN(n630) );
  INV_X1 U686 ( .A(n626), .ZN(n643) );
  NOR2_X1 U687 ( .A1(n643), .A2(G1348), .ZN(n628) );
  NOR2_X1 U688 ( .A1(G2067), .A2(n626), .ZN(n627) );
  NOR2_X1 U689 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U690 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U691 ( .A1(n632), .A2(n631), .ZN(n637) );
  INV_X1 U692 ( .A(G299), .ZN(n976) );
  NAND2_X1 U693 ( .A1(n643), .A2(G2072), .ZN(n633) );
  XNOR2_X1 U694 ( .A(n633), .B(KEYINPUT27), .ZN(n635) );
  INV_X1 U695 ( .A(G1956), .ZN(n996) );
  NOR2_X1 U696 ( .A1(n996), .A2(n643), .ZN(n634) );
  NOR2_X1 U697 ( .A1(n635), .A2(n634), .ZN(n638) );
  NAND2_X1 U698 ( .A1(n976), .A2(n638), .ZN(n636) );
  NAND2_X1 U699 ( .A1(n637), .A2(n636), .ZN(n641) );
  NOR2_X1 U700 ( .A1(n976), .A2(n638), .ZN(n639) );
  XOR2_X1 U701 ( .A(n639), .B(KEYINPUT28), .Z(n640) );
  NAND2_X1 U702 ( .A1(n641), .A2(n640), .ZN(n642) );
  XOR2_X1 U703 ( .A(KEYINPUT29), .B(n642), .Z(n647) );
  XNOR2_X1 U704 ( .A(G1961), .B(KEYINPUT99), .ZN(n993) );
  NAND2_X1 U705 ( .A1(n626), .A2(n993), .ZN(n645) );
  XNOR2_X1 U706 ( .A(G2078), .B(KEYINPUT25), .ZN(n945) );
  NAND2_X1 U707 ( .A1(n643), .A2(n945), .ZN(n644) );
  NAND2_X1 U708 ( .A1(n645), .A2(n644), .ZN(n652) );
  NAND2_X1 U709 ( .A1(n652), .A2(G171), .ZN(n646) );
  NAND2_X1 U710 ( .A1(n647), .A2(n646), .ZN(n657) );
  NAND2_X1 U711 ( .A1(G8), .A2(n626), .ZN(n692) );
  NOR2_X1 U712 ( .A1(G1966), .A2(n692), .ZN(n659) );
  NOR2_X1 U713 ( .A1(n659), .A2(n648), .ZN(n649) );
  NAND2_X1 U714 ( .A1(G8), .A2(n649), .ZN(n650) );
  XNOR2_X1 U715 ( .A(KEYINPUT30), .B(n650), .ZN(n651) );
  NOR2_X1 U716 ( .A1(G168), .A2(n651), .ZN(n654) );
  NOR2_X1 U717 ( .A1(G171), .A2(n652), .ZN(n653) );
  NOR2_X1 U718 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U719 ( .A(KEYINPUT31), .B(n655), .Z(n656) );
  NAND2_X1 U720 ( .A1(n657), .A2(n656), .ZN(n662) );
  NAND2_X1 U721 ( .A1(n658), .A2(n662), .ZN(n660) );
  NOR2_X1 U722 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U723 ( .A(n661), .B(KEYINPUT101), .ZN(n685) );
  NAND2_X1 U724 ( .A1(G1976), .A2(G288), .ZN(n979) );
  AND2_X1 U725 ( .A1(n685), .A2(n979), .ZN(n671) );
  NAND2_X1 U726 ( .A1(G286), .A2(n662), .ZN(n663) );
  XNOR2_X1 U727 ( .A(n663), .B(KEYINPUT102), .ZN(n668) );
  NOR2_X1 U728 ( .A1(G1971), .A2(n692), .ZN(n665) );
  NOR2_X1 U729 ( .A1(G2090), .A2(n626), .ZN(n664) );
  NOR2_X1 U730 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U731 ( .A1(n666), .A2(G303), .ZN(n667) );
  NAND2_X1 U732 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U733 ( .A1(n669), .A2(G8), .ZN(n670) );
  XNOR2_X1 U734 ( .A(n670), .B(KEYINPUT32), .ZN(n684) );
  AND2_X1 U735 ( .A1(n671), .A2(n684), .ZN(n679) );
  INV_X1 U736 ( .A(n979), .ZN(n674) );
  NOR2_X1 U737 ( .A1(G1976), .A2(G288), .ZN(n981) );
  NOR2_X1 U738 ( .A1(G1971), .A2(G303), .ZN(n672) );
  NOR2_X1 U739 ( .A1(n981), .A2(n672), .ZN(n673) );
  OR2_X1 U740 ( .A1(n674), .A2(n673), .ZN(n675) );
  OR2_X1 U741 ( .A1(n692), .A2(n675), .ZN(n677) );
  INV_X1 U742 ( .A(KEYINPUT33), .ZN(n676) );
  NAND2_X1 U743 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U744 ( .A1(n679), .A2(n678), .ZN(n682) );
  NAND2_X1 U745 ( .A1(n981), .A2(KEYINPUT33), .ZN(n680) );
  NOR2_X1 U746 ( .A1(n680), .A2(n692), .ZN(n681) );
  NOR2_X1 U747 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U748 ( .A(G1981), .B(G305), .Z(n967) );
  AND2_X1 U749 ( .A1(n683), .A2(n967), .ZN(n697) );
  NAND2_X1 U750 ( .A1(n685), .A2(n684), .ZN(n688) );
  NOR2_X1 U751 ( .A1(G2090), .A2(G303), .ZN(n686) );
  NAND2_X1 U752 ( .A1(G8), .A2(n686), .ZN(n687) );
  NAND2_X1 U753 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U754 ( .A1(n689), .A2(n692), .ZN(n695) );
  NOR2_X1 U755 ( .A1(G1981), .A2(G305), .ZN(n690) );
  XNOR2_X1 U756 ( .A(n690), .B(KEYINPUT24), .ZN(n691) );
  XNOR2_X1 U757 ( .A(n691), .B(KEYINPUT97), .ZN(n693) );
  OR2_X1 U758 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U759 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X2 U760 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U761 ( .A(n698), .B(KEYINPUT103), .ZN(n733) );
  XNOR2_X1 U762 ( .A(G1986), .B(G290), .ZN(n974) );
  NOR2_X1 U763 ( .A1(n700), .A2(n699), .ZN(n745) );
  NAND2_X1 U764 ( .A1(n974), .A2(n745), .ZN(n731) );
  NAND2_X1 U765 ( .A1(G95), .A2(n898), .ZN(n702) );
  NAND2_X1 U766 ( .A1(G131), .A2(n895), .ZN(n701) );
  NAND2_X1 U767 ( .A1(n702), .A2(n701), .ZN(n706) );
  NAND2_X1 U768 ( .A1(G107), .A2(n891), .ZN(n704) );
  NAND2_X1 U769 ( .A1(G119), .A2(n889), .ZN(n703) );
  NAND2_X1 U770 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U771 ( .A1(n706), .A2(n705), .ZN(n869) );
  INV_X1 U772 ( .A(G1991), .ZN(n734) );
  NOR2_X1 U773 ( .A1(n869), .A2(n734), .ZN(n715) );
  NAND2_X1 U774 ( .A1(G117), .A2(n891), .ZN(n708) );
  NAND2_X1 U775 ( .A1(G129), .A2(n889), .ZN(n707) );
  NAND2_X1 U776 ( .A1(n708), .A2(n707), .ZN(n711) );
  NAND2_X1 U777 ( .A1(n898), .A2(G105), .ZN(n709) );
  XOR2_X1 U778 ( .A(KEYINPUT38), .B(n709), .Z(n710) );
  NOR2_X1 U779 ( .A1(n711), .A2(n710), .ZN(n713) );
  NAND2_X1 U780 ( .A1(n895), .A2(G141), .ZN(n712) );
  NAND2_X1 U781 ( .A1(n713), .A2(n712), .ZN(n885) );
  AND2_X1 U782 ( .A1(n885), .A2(G1996), .ZN(n714) );
  NOR2_X1 U783 ( .A1(n715), .A2(n714), .ZN(n931) );
  INV_X1 U784 ( .A(n745), .ZN(n716) );
  NOR2_X1 U785 ( .A1(n931), .A2(n716), .ZN(n737) );
  INV_X1 U786 ( .A(n737), .ZN(n728) );
  XNOR2_X1 U787 ( .A(G2067), .B(KEYINPUT37), .ZN(n717) );
  XNOR2_X1 U788 ( .A(n717), .B(KEYINPUT94), .ZN(n742) );
  NAND2_X1 U789 ( .A1(G104), .A2(n898), .ZN(n719) );
  NAND2_X1 U790 ( .A1(G140), .A2(n895), .ZN(n718) );
  NAND2_X1 U791 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U792 ( .A(KEYINPUT34), .B(n720), .ZN(n725) );
  NAND2_X1 U793 ( .A1(G116), .A2(n891), .ZN(n722) );
  NAND2_X1 U794 ( .A1(G128), .A2(n889), .ZN(n721) );
  NAND2_X1 U795 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U796 ( .A(n723), .B(KEYINPUT35), .Z(n724) );
  NOR2_X1 U797 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U798 ( .A(KEYINPUT36), .B(n726), .Z(n727) );
  XNOR2_X1 U799 ( .A(KEYINPUT95), .B(n727), .ZN(n880) );
  NOR2_X1 U800 ( .A1(n742), .A2(n880), .ZN(n920) );
  NAND2_X1 U801 ( .A1(n745), .A2(n920), .ZN(n740) );
  NAND2_X1 U802 ( .A1(n728), .A2(n740), .ZN(n729) );
  XOR2_X1 U803 ( .A(n729), .B(KEYINPUT96), .Z(n730) );
  AND2_X1 U804 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U805 ( .A1(n733), .A2(n732), .ZN(n748) );
  NOR2_X1 U806 ( .A1(G1996), .A2(n885), .ZN(n933) );
  AND2_X1 U807 ( .A1(n734), .A2(n869), .ZN(n919) );
  NOR2_X1 U808 ( .A1(G1986), .A2(G290), .ZN(n735) );
  NOR2_X1 U809 ( .A1(n919), .A2(n735), .ZN(n736) );
  NOR2_X1 U810 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U811 ( .A1(n933), .A2(n738), .ZN(n739) );
  XNOR2_X1 U812 ( .A(n739), .B(KEYINPUT39), .ZN(n741) );
  NAND2_X1 U813 ( .A1(n741), .A2(n740), .ZN(n743) );
  NAND2_X1 U814 ( .A1(n742), .A2(n880), .ZN(n930) );
  NAND2_X1 U815 ( .A1(n743), .A2(n930), .ZN(n744) );
  XNOR2_X1 U816 ( .A(KEYINPUT104), .B(n744), .ZN(n746) );
  NAND2_X1 U817 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U818 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U819 ( .A(n749), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U820 ( .A(G2443), .B(G2446), .Z(n752) );
  XNOR2_X1 U821 ( .A(G2427), .B(G2451), .ZN(n751) );
  XNOR2_X1 U822 ( .A(n752), .B(n751), .ZN(n758) );
  XOR2_X1 U823 ( .A(G2430), .B(G2454), .Z(n754) );
  XNOR2_X1 U824 ( .A(G1348), .B(G1341), .ZN(n753) );
  XNOR2_X1 U825 ( .A(n754), .B(n753), .ZN(n756) );
  XOR2_X1 U826 ( .A(G2435), .B(G2438), .Z(n755) );
  XNOR2_X1 U827 ( .A(n756), .B(n755), .ZN(n757) );
  XOR2_X1 U828 ( .A(n758), .B(n757), .Z(n759) );
  AND2_X1 U829 ( .A1(G14), .A2(n759), .ZN(G401) );
  AND2_X1 U830 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U831 ( .A(G120), .ZN(G236) );
  INV_X1 U832 ( .A(G69), .ZN(G235) );
  INV_X1 U833 ( .A(G108), .ZN(G238) );
  INV_X1 U834 ( .A(G132), .ZN(G219) );
  NAND2_X1 U835 ( .A1(G7), .A2(G661), .ZN(n760) );
  XNOR2_X1 U836 ( .A(n760), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U837 ( .A(G223), .B(KEYINPUT69), .ZN(n831) );
  NAND2_X1 U838 ( .A1(n831), .A2(G567), .ZN(n761) );
  XOR2_X1 U839 ( .A(KEYINPUT11), .B(n761), .Z(G234) );
  INV_X1 U840 ( .A(G860), .ZN(n787) );
  OR2_X1 U841 ( .A1(n986), .A2(n787), .ZN(G153) );
  INV_X1 U842 ( .A(G171), .ZN(G301) );
  NAND2_X1 U843 ( .A1(G868), .A2(G301), .ZN(n763) );
  OR2_X1 U844 ( .A1(n970), .A2(G868), .ZN(n762) );
  NAND2_X1 U845 ( .A1(n763), .A2(n762), .ZN(G284) );
  INV_X1 U846 ( .A(G868), .ZN(n764) );
  NOR2_X1 U847 ( .A1(G286), .A2(n764), .ZN(n766) );
  NOR2_X1 U848 ( .A1(G868), .A2(G299), .ZN(n765) );
  NOR2_X1 U849 ( .A1(n766), .A2(n765), .ZN(n767) );
  XOR2_X1 U850 ( .A(KEYINPUT73), .B(n767), .Z(G297) );
  NAND2_X1 U851 ( .A1(n787), .A2(G559), .ZN(n768) );
  NAND2_X1 U852 ( .A1(n768), .A2(n970), .ZN(n769) );
  XNOR2_X1 U853 ( .A(n769), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U854 ( .A1(G868), .A2(n986), .ZN(n770) );
  XNOR2_X1 U855 ( .A(KEYINPUT74), .B(n770), .ZN(n773) );
  NAND2_X1 U856 ( .A1(G868), .A2(n970), .ZN(n771) );
  NOR2_X1 U857 ( .A1(G559), .A2(n771), .ZN(n772) );
  NOR2_X1 U858 ( .A1(n773), .A2(n772), .ZN(G282) );
  XOR2_X1 U859 ( .A(G2100), .B(KEYINPUT78), .Z(n785) );
  XOR2_X1 U860 ( .A(G2096), .B(KEYINPUT77), .Z(n783) );
  NAND2_X1 U861 ( .A1(G111), .A2(n891), .ZN(n774) );
  XNOR2_X1 U862 ( .A(n774), .B(KEYINPUT76), .ZN(n778) );
  XOR2_X1 U863 ( .A(KEYINPUT75), .B(KEYINPUT18), .Z(n776) );
  NAND2_X1 U864 ( .A1(G123), .A2(n889), .ZN(n775) );
  XNOR2_X1 U865 ( .A(n776), .B(n775), .ZN(n777) );
  NAND2_X1 U866 ( .A1(n778), .A2(n777), .ZN(n782) );
  NAND2_X1 U867 ( .A1(G99), .A2(n898), .ZN(n780) );
  NAND2_X1 U868 ( .A1(G135), .A2(n895), .ZN(n779) );
  NAND2_X1 U869 ( .A1(n780), .A2(n779), .ZN(n781) );
  NOR2_X1 U870 ( .A1(n782), .A2(n781), .ZN(n918) );
  XNOR2_X1 U871 ( .A(n783), .B(n918), .ZN(n784) );
  NAND2_X1 U872 ( .A1(n785), .A2(n784), .ZN(G156) );
  NAND2_X1 U873 ( .A1(G559), .A2(n970), .ZN(n786) );
  XOR2_X1 U874 ( .A(n986), .B(n786), .Z(n807) );
  NAND2_X1 U875 ( .A1(n787), .A2(n807), .ZN(n801) );
  NAND2_X1 U876 ( .A1(n788), .A2(G80), .ZN(n789) );
  XOR2_X1 U877 ( .A(KEYINPUT79), .B(n789), .Z(n792) );
  NAND2_X1 U878 ( .A1(n790), .A2(G93), .ZN(n791) );
  NAND2_X1 U879 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U880 ( .A(KEYINPUT80), .B(n793), .Z(n796) );
  NAND2_X1 U881 ( .A1(n794), .A2(G55), .ZN(n795) );
  NAND2_X1 U882 ( .A1(n796), .A2(n795), .ZN(n800) );
  NAND2_X1 U883 ( .A1(G67), .A2(n797), .ZN(n798) );
  XNOR2_X1 U884 ( .A(KEYINPUT81), .B(n798), .ZN(n799) );
  NOR2_X1 U885 ( .A1(n800), .A2(n799), .ZN(n809) );
  XOR2_X1 U886 ( .A(n801), .B(n809), .Z(G145) );
  XNOR2_X1 U887 ( .A(KEYINPUT19), .B(G299), .ZN(n802) );
  XNOR2_X1 U888 ( .A(n802), .B(G305), .ZN(n803) );
  XNOR2_X1 U889 ( .A(n809), .B(n803), .ZN(n805) );
  XNOR2_X1 U890 ( .A(G290), .B(G166), .ZN(n804) );
  XNOR2_X1 U891 ( .A(n805), .B(n804), .ZN(n806) );
  XNOR2_X1 U892 ( .A(n806), .B(G288), .ZN(n907) );
  XNOR2_X1 U893 ( .A(n807), .B(n907), .ZN(n808) );
  NAND2_X1 U894 ( .A1(n808), .A2(G868), .ZN(n811) );
  OR2_X1 U895 ( .A1(G868), .A2(n809), .ZN(n810) );
  NAND2_X1 U896 ( .A1(n811), .A2(n810), .ZN(G295) );
  XOR2_X1 U897 ( .A(KEYINPUT21), .B(KEYINPUT85), .Z(n815) );
  NAND2_X1 U898 ( .A1(G2078), .A2(G2084), .ZN(n812) );
  XOR2_X1 U899 ( .A(KEYINPUT20), .B(n812), .Z(n813) );
  NAND2_X1 U900 ( .A1(n813), .A2(G2090), .ZN(n814) );
  XNOR2_X1 U901 ( .A(n815), .B(n814), .ZN(n816) );
  NAND2_X1 U902 ( .A1(G2072), .A2(n816), .ZN(G158) );
  XNOR2_X1 U903 ( .A(KEYINPUT86), .B(G44), .ZN(n817) );
  XNOR2_X1 U904 ( .A(n817), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U905 ( .A(KEYINPUT68), .B(G82), .Z(G220) );
  NOR2_X1 U906 ( .A1(G220), .A2(G219), .ZN(n819) );
  XNOR2_X1 U907 ( .A(KEYINPUT22), .B(KEYINPUT87), .ZN(n818) );
  XNOR2_X1 U908 ( .A(n819), .B(n818), .ZN(n820) );
  NOR2_X1 U909 ( .A1(G218), .A2(n820), .ZN(n821) );
  XNOR2_X1 U910 ( .A(KEYINPUT88), .B(n821), .ZN(n822) );
  NAND2_X1 U911 ( .A1(n822), .A2(G96), .ZN(n836) );
  NAND2_X1 U912 ( .A1(n836), .A2(G2106), .ZN(n828) );
  NOR2_X1 U913 ( .A1(G235), .A2(G236), .ZN(n823) );
  XNOR2_X1 U914 ( .A(n823), .B(KEYINPUT89), .ZN(n824) );
  NOR2_X1 U915 ( .A1(G238), .A2(n824), .ZN(n825) );
  NAND2_X1 U916 ( .A1(G57), .A2(n825), .ZN(n837) );
  NAND2_X1 U917 ( .A1(G567), .A2(n837), .ZN(n826) );
  XNOR2_X1 U918 ( .A(KEYINPUT90), .B(n826), .ZN(n827) );
  NAND2_X1 U919 ( .A1(n828), .A2(n827), .ZN(n839) );
  NAND2_X1 U920 ( .A1(G483), .A2(G661), .ZN(n829) );
  NOR2_X1 U921 ( .A1(n839), .A2(n829), .ZN(n835) );
  NAND2_X1 U922 ( .A1(n835), .A2(G36), .ZN(n830) );
  XOR2_X1 U923 ( .A(KEYINPUT91), .B(n830), .Z(G176) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n831), .ZN(G217) );
  NAND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n832) );
  XNOR2_X1 U926 ( .A(KEYINPUT105), .B(n832), .ZN(n833) );
  NAND2_X1 U927 ( .A1(n833), .A2(G661), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U929 ( .A1(n835), .A2(n834), .ZN(G188) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  NOR2_X1 U932 ( .A1(n837), .A2(n836), .ZN(n838) );
  XNOR2_X1 U933 ( .A(n838), .B(KEYINPUT106), .ZN(G325) );
  INV_X1 U934 ( .A(G325), .ZN(G261) );
  INV_X1 U935 ( .A(n839), .ZN(G319) );
  XOR2_X1 U936 ( .A(KEYINPUT42), .B(G2090), .Z(n841) );
  XNOR2_X1 U937 ( .A(G2078), .B(G2072), .ZN(n840) );
  XNOR2_X1 U938 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U939 ( .A(n842), .B(G2096), .Z(n844) );
  XNOR2_X1 U940 ( .A(G2067), .B(G2084), .ZN(n843) );
  XNOR2_X1 U941 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U942 ( .A(G2100), .B(KEYINPUT43), .Z(n846) );
  XNOR2_X1 U943 ( .A(G2678), .B(KEYINPUT107), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U945 ( .A(n848), .B(n847), .Z(G227) );
  XOR2_X1 U946 ( .A(G1976), .B(G1971), .Z(n850) );
  XNOR2_X1 U947 ( .A(G1966), .B(G1956), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U949 ( .A(n851), .B(KEYINPUT41), .Z(n853) );
  XNOR2_X1 U950 ( .A(G1996), .B(G1991), .ZN(n852) );
  XNOR2_X1 U951 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U952 ( .A(G2474), .B(G1981), .Z(n855) );
  XNOR2_X1 U953 ( .A(G1986), .B(G1961), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(n856) );
  XNOR2_X1 U955 ( .A(n857), .B(n856), .ZN(G229) );
  NAND2_X1 U956 ( .A1(n895), .A2(G136), .ZN(n864) );
  NAND2_X1 U957 ( .A1(G112), .A2(n891), .ZN(n859) );
  NAND2_X1 U958 ( .A1(G100), .A2(n898), .ZN(n858) );
  NAND2_X1 U959 ( .A1(n859), .A2(n858), .ZN(n862) );
  NAND2_X1 U960 ( .A1(n889), .A2(G124), .ZN(n860) );
  XOR2_X1 U961 ( .A(KEYINPUT44), .B(n860), .Z(n861) );
  NOR2_X1 U962 ( .A1(n862), .A2(n861), .ZN(n863) );
  NAND2_X1 U963 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U964 ( .A(KEYINPUT108), .B(n865), .Z(G162) );
  XOR2_X1 U965 ( .A(KEYINPUT110), .B(KEYINPUT46), .Z(n867) );
  XNOR2_X1 U966 ( .A(KEYINPUT115), .B(KEYINPUT48), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U968 ( .A(n868), .B(KEYINPUT114), .Z(n871) );
  XNOR2_X1 U969 ( .A(n869), .B(n918), .ZN(n870) );
  XNOR2_X1 U970 ( .A(n871), .B(n870), .ZN(n884) );
  NAND2_X1 U971 ( .A1(G118), .A2(n891), .ZN(n873) );
  NAND2_X1 U972 ( .A1(G130), .A2(n889), .ZN(n872) );
  NAND2_X1 U973 ( .A1(n873), .A2(n872), .ZN(n879) );
  NAND2_X1 U974 ( .A1(G106), .A2(n898), .ZN(n875) );
  NAND2_X1 U975 ( .A1(G142), .A2(n895), .ZN(n874) );
  NAND2_X1 U976 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U977 ( .A(KEYINPUT45), .B(n876), .ZN(n877) );
  XNOR2_X1 U978 ( .A(KEYINPUT109), .B(n877), .ZN(n878) );
  NOR2_X1 U979 ( .A1(n879), .A2(n878), .ZN(n881) );
  XNOR2_X1 U980 ( .A(n881), .B(n880), .ZN(n882) );
  XNOR2_X1 U981 ( .A(n882), .B(G162), .ZN(n883) );
  XNOR2_X1 U982 ( .A(n884), .B(n883), .ZN(n887) );
  XOR2_X1 U983 ( .A(G164), .B(n885), .Z(n886) );
  XNOR2_X1 U984 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U985 ( .A(n888), .B(G160), .ZN(n903) );
  NAND2_X1 U986 ( .A1(n889), .A2(G127), .ZN(n890) );
  XNOR2_X1 U987 ( .A(n890), .B(KEYINPUT112), .ZN(n893) );
  NAND2_X1 U988 ( .A1(G115), .A2(n891), .ZN(n892) );
  NAND2_X1 U989 ( .A1(n893), .A2(n892), .ZN(n894) );
  XNOR2_X1 U990 ( .A(n894), .B(KEYINPUT47), .ZN(n897) );
  NAND2_X1 U991 ( .A1(G139), .A2(n895), .ZN(n896) );
  NAND2_X1 U992 ( .A1(n897), .A2(n896), .ZN(n901) );
  NAND2_X1 U993 ( .A1(G103), .A2(n898), .ZN(n899) );
  XNOR2_X1 U994 ( .A(KEYINPUT111), .B(n899), .ZN(n900) );
  NOR2_X1 U995 ( .A1(n901), .A2(n900), .ZN(n902) );
  XNOR2_X1 U996 ( .A(KEYINPUT113), .B(n902), .ZN(n924) );
  XNOR2_X1 U997 ( .A(n903), .B(n924), .ZN(n904) );
  NOR2_X1 U998 ( .A1(G37), .A2(n904), .ZN(G395) );
  XNOR2_X1 U999 ( .A(n986), .B(G286), .ZN(n906) );
  XNOR2_X1 U1000 ( .A(G171), .B(n970), .ZN(n905) );
  XNOR2_X1 U1001 ( .A(n906), .B(n905), .ZN(n908) );
  XNOR2_X1 U1002 ( .A(n908), .B(n907), .ZN(n909) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n909), .ZN(G397) );
  NOR2_X1 U1004 ( .A1(G227), .A2(G229), .ZN(n911) );
  XNOR2_X1 U1005 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n910) );
  XNOR2_X1 U1006 ( .A(n911), .B(n910), .ZN(n912) );
  NOR2_X1 U1007 ( .A1(G401), .A2(n912), .ZN(n913) );
  AND2_X1 U1008 ( .A1(G319), .A2(n913), .ZN(n915) );
  NOR2_X1 U1009 ( .A1(G395), .A2(G397), .ZN(n914) );
  NAND2_X1 U1010 ( .A1(n915), .A2(n914), .ZN(G225) );
  INV_X1 U1011 ( .A(G225), .ZN(G308) );
  INV_X1 U1012 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1013 ( .A(G2084), .B(KEYINPUT117), .ZN(n916) );
  XNOR2_X1 U1014 ( .A(n916), .B(G160), .ZN(n917) );
  NOR2_X1 U1015 ( .A1(n918), .A2(n917), .ZN(n922) );
  NOR2_X1 U1016 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1017 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1018 ( .A(KEYINPUT118), .B(n923), .ZN(n940) );
  XNOR2_X1 U1019 ( .A(KEYINPUT119), .B(n924), .ZN(n925) );
  XOR2_X1 U1020 ( .A(G2072), .B(n925), .Z(n927) );
  XOR2_X1 U1021 ( .A(G164), .B(G2078), .Z(n926) );
  NOR2_X1 U1022 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1023 ( .A(KEYINPUT50), .B(n928), .ZN(n929) );
  XNOR2_X1 U1024 ( .A(n929), .B(KEYINPUT120), .ZN(n938) );
  NAND2_X1 U1025 ( .A1(n931), .A2(n930), .ZN(n936) );
  XOR2_X1 U1026 ( .A(G2090), .B(G162), .Z(n932) );
  NOR2_X1 U1027 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1028 ( .A(n934), .B(KEYINPUT51), .ZN(n935) );
  NOR2_X1 U1029 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1030 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1031 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1032 ( .A(KEYINPUT52), .B(n941), .ZN(n942) );
  INV_X1 U1033 ( .A(KEYINPUT55), .ZN(n963) );
  NAND2_X1 U1034 ( .A1(n942), .A2(n963), .ZN(n943) );
  NAND2_X1 U1035 ( .A1(n943), .A2(G29), .ZN(n1026) );
  XNOR2_X1 U1036 ( .A(G2090), .B(G35), .ZN(n958) );
  XOR2_X1 U1037 ( .A(G2072), .B(G33), .Z(n944) );
  NAND2_X1 U1038 ( .A1(n944), .A2(G28), .ZN(n955) );
  XNOR2_X1 U1039 ( .A(n945), .B(G27), .ZN(n948) );
  XNOR2_X1 U1040 ( .A(n946), .B(G32), .ZN(n947) );
  NAND2_X1 U1041 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1042 ( .A(KEYINPUT121), .B(n949), .ZN(n953) );
  XNOR2_X1 U1043 ( .A(G2067), .B(G26), .ZN(n951) );
  XNOR2_X1 U1044 ( .A(G1991), .B(G25), .ZN(n950) );
  NOR2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1047 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1048 ( .A(KEYINPUT53), .B(n956), .ZN(n957) );
  NOR2_X1 U1049 ( .A1(n958), .A2(n957), .ZN(n961) );
  XOR2_X1 U1050 ( .A(G2084), .B(KEYINPUT54), .Z(n959) );
  XNOR2_X1 U1051 ( .A(G34), .B(n959), .ZN(n960) );
  NAND2_X1 U1052 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1053 ( .A(n963), .B(n962), .ZN(n965) );
  INV_X1 U1054 ( .A(G29), .ZN(n964) );
  NAND2_X1 U1055 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1056 ( .A1(G11), .A2(n966), .ZN(n1024) );
  XNOR2_X1 U1057 ( .A(G16), .B(KEYINPUT56), .ZN(n992) );
  XNOR2_X1 U1058 ( .A(G1966), .B(G168), .ZN(n968) );
  NAND2_X1 U1059 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1060 ( .A(n969), .B(KEYINPUT57), .ZN(n990) );
  XNOR2_X1 U1061 ( .A(G1348), .B(n970), .ZN(n972) );
  XNOR2_X1 U1062 ( .A(G171), .B(G1961), .ZN(n971) );
  NAND2_X1 U1063 ( .A1(n972), .A2(n971), .ZN(n973) );
  NOR2_X1 U1064 ( .A1(n974), .A2(n973), .ZN(n985) );
  XNOR2_X1 U1065 ( .A(G1971), .B(KEYINPUT122), .ZN(n975) );
  XNOR2_X1 U1066 ( .A(n975), .B(G303), .ZN(n978) );
  XNOR2_X1 U1067 ( .A(n976), .B(n996), .ZN(n977) );
  NOR2_X1 U1068 ( .A1(n978), .A2(n977), .ZN(n980) );
  NAND2_X1 U1069 ( .A1(n980), .A2(n979), .ZN(n982) );
  NOR2_X1 U1070 ( .A1(n982), .A2(n981), .ZN(n983) );
  XOR2_X1 U1071 ( .A(KEYINPUT123), .B(n983), .Z(n984) );
  NAND2_X1 U1072 ( .A1(n985), .A2(n984), .ZN(n988) );
  XNOR2_X1 U1073 ( .A(G1341), .B(n986), .ZN(n987) );
  NOR2_X1 U1074 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1075 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1076 ( .A1(n992), .A2(n991), .ZN(n1022) );
  INV_X1 U1077 ( .A(G16), .ZN(n1020) );
  XNOR2_X1 U1078 ( .A(n993), .B(G5), .ZN(n1016) );
  XOR2_X1 U1079 ( .A(G1966), .B(G21), .Z(n1006) );
  XOR2_X1 U1080 ( .A(G4), .B(KEYINPUT124), .Z(n995) );
  XNOR2_X1 U1081 ( .A(G1348), .B(KEYINPUT59), .ZN(n994) );
  XNOR2_X1 U1082 ( .A(n995), .B(n994), .ZN(n1002) );
  XNOR2_X1 U1083 ( .A(G20), .B(n996), .ZN(n1000) );
  XNOR2_X1 U1084 ( .A(G1341), .B(G19), .ZN(n998) );
  XNOR2_X1 U1085 ( .A(G1981), .B(G6), .ZN(n997) );
  NOR2_X1 U1086 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1087 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1088 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1089 ( .A(KEYINPUT125), .B(n1003), .Z(n1004) );
  XNOR2_X1 U1090 ( .A(KEYINPUT60), .B(n1004), .ZN(n1005) );
  NAND2_X1 U1091 ( .A1(n1006), .A2(n1005), .ZN(n1014) );
  XNOR2_X1 U1092 ( .A(G1986), .B(G24), .ZN(n1008) );
  XNOR2_X1 U1093 ( .A(G1971), .B(G22), .ZN(n1007) );
  NOR2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1011) );
  XOR2_X1 U1095 ( .A(G1976), .B(KEYINPUT126), .Z(n1009) );
  XNOR2_X1 U1096 ( .A(G23), .B(n1009), .ZN(n1010) );
  NAND2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1098 ( .A(KEYINPUT58), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1099 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1100 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1101 ( .A(n1017), .B(KEYINPUT61), .ZN(n1018) );
  XNOR2_X1 U1102 ( .A(KEYINPUT127), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1103 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1104 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1105 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1106 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1027), .Z(G311) );
  INV_X1 U1108 ( .A(G311), .ZN(G150) );
endmodule

