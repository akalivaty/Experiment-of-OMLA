

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U554 ( .A(n661), .ZN(n648) );
  XNOR2_X1 U555 ( .A(n601), .B(KEYINPUT30), .ZN(n602) );
  NOR2_X1 U556 ( .A1(n695), .A2(n694), .ZN(n699) );
  NOR2_X2 U557 ( .A1(n528), .A2(n527), .ZN(G160) );
  XNOR2_X2 U558 ( .A(n517), .B(KEYINPUT66), .ZN(n715) );
  INV_X1 U559 ( .A(KEYINPUT91), .ZN(n601) );
  XNOR2_X1 U560 ( .A(n603), .B(n602), .ZN(n604) );
  INV_X1 U561 ( .A(KEYINPUT92), .ZN(n605) );
  XNOR2_X1 U562 ( .A(n612), .B(KEYINPUT31), .ZN(n613) );
  XNOR2_X1 U563 ( .A(n614), .B(n613), .ZN(n677) );
  INV_X1 U564 ( .A(KEYINPUT100), .ZN(n709) );
  XNOR2_X1 U565 ( .A(n710), .B(n709), .ZN(n740) );
  INV_X1 U566 ( .A(KEYINPUT13), .ZN(n636) );
  INV_X1 U567 ( .A(KEYINPUT17), .ZN(n521) );
  NOR2_X2 U568 ( .A1(G2104), .A2(n519), .ZN(n895) );
  XOR2_X1 U569 ( .A(G543), .B(KEYINPUT0), .Z(n540) );
  NAND2_X1 U570 ( .A1(n889), .A2(G137), .ZN(n524) );
  NOR2_X1 U571 ( .A1(G651), .A2(n578), .ZN(n796) );
  NAND2_X1 U572 ( .A1(n641), .A2(n640), .ZN(n946) );
  NAND2_X1 U573 ( .A1(n526), .A2(n525), .ZN(n527) );
  NOR2_X1 U574 ( .A1(n537), .A2(n536), .ZN(G164) );
  INV_X1 U575 ( .A(G2105), .ZN(n519) );
  AND2_X1 U576 ( .A1(G2104), .A2(n519), .ZN(n517) );
  NAND2_X1 U577 ( .A1(n715), .A2(G101), .ZN(n518) );
  XNOR2_X1 U578 ( .A(KEYINPUT23), .B(n518), .ZN(n528) );
  NAND2_X1 U579 ( .A1(G125), .A2(n895), .ZN(n520) );
  XOR2_X1 U580 ( .A(KEYINPUT65), .B(n520), .Z(n526) );
  NOR2_X1 U581 ( .A1(G2104), .A2(G2105), .ZN(n522) );
  XNOR2_X2 U582 ( .A(n522), .B(n521), .ZN(n889) );
  AND2_X1 U583 ( .A1(G2104), .A2(G2105), .ZN(n898) );
  NAND2_X1 U584 ( .A1(G113), .A2(n898), .ZN(n523) );
  AND2_X1 U585 ( .A1(n524), .A2(n523), .ZN(n525) );
  NAND2_X1 U586 ( .A1(G114), .A2(n898), .ZN(n530) );
  NAND2_X1 U587 ( .A1(G126), .A2(n895), .ZN(n529) );
  NAND2_X1 U588 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U589 ( .A(n531), .B(KEYINPUT83), .ZN(n533) );
  NAND2_X1 U590 ( .A1(G102), .A2(n715), .ZN(n532) );
  NAND2_X1 U591 ( .A1(n533), .A2(n532), .ZN(n537) );
  NAND2_X1 U592 ( .A1(n889), .A2(G138), .ZN(n535) );
  INV_X1 U593 ( .A(KEYINPUT84), .ZN(n534) );
  XNOR2_X1 U594 ( .A(n535), .B(n534), .ZN(n536) );
  NOR2_X1 U595 ( .A1(G543), .A2(G651), .ZN(n538) );
  XNOR2_X1 U596 ( .A(n538), .B(KEYINPUT64), .ZN(n793) );
  NAND2_X1 U597 ( .A1(G89), .A2(n793), .ZN(n539) );
  XNOR2_X1 U598 ( .A(n539), .B(KEYINPUT4), .ZN(n543) );
  INV_X1 U599 ( .A(G651), .ZN(n545) );
  XOR2_X1 U600 ( .A(KEYINPUT67), .B(n540), .Z(n578) );
  OR2_X1 U601 ( .A1(n545), .A2(n578), .ZN(n541) );
  XOR2_X2 U602 ( .A(KEYINPUT68), .B(n541), .Z(n797) );
  NAND2_X1 U603 ( .A1(G76), .A2(n797), .ZN(n542) );
  NAND2_X1 U604 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U605 ( .A(n544), .B(KEYINPUT5), .ZN(n551) );
  NOR2_X1 U606 ( .A1(G543), .A2(n545), .ZN(n546) );
  XOR2_X1 U607 ( .A(KEYINPUT1), .B(n546), .Z(n792) );
  NAND2_X1 U608 ( .A1(G63), .A2(n792), .ZN(n548) );
  NAND2_X1 U609 ( .A1(G51), .A2(n796), .ZN(n547) );
  NAND2_X1 U610 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U611 ( .A(KEYINPUT6), .B(n549), .Z(n550) );
  NAND2_X1 U612 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U613 ( .A(n552), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U614 ( .A1(G64), .A2(n792), .ZN(n554) );
  NAND2_X1 U615 ( .A1(G52), .A2(n796), .ZN(n553) );
  NAND2_X1 U616 ( .A1(n554), .A2(n553), .ZN(n559) );
  NAND2_X1 U617 ( .A1(G90), .A2(n793), .ZN(n556) );
  NAND2_X1 U618 ( .A1(G77), .A2(n797), .ZN(n555) );
  NAND2_X1 U619 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U620 ( .A(KEYINPUT9), .B(n557), .Z(n558) );
  NOR2_X1 U621 ( .A1(n559), .A2(n558), .ZN(G171) );
  INV_X1 U622 ( .A(G171), .ZN(G301) );
  NAND2_X1 U623 ( .A1(G65), .A2(n792), .ZN(n561) );
  NAND2_X1 U624 ( .A1(G53), .A2(n796), .ZN(n560) );
  NAND2_X1 U625 ( .A1(n561), .A2(n560), .ZN(n565) );
  NAND2_X1 U626 ( .A1(G91), .A2(n793), .ZN(n563) );
  NAND2_X1 U627 ( .A1(G78), .A2(n797), .ZN(n562) );
  NAND2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n564) );
  OR2_X1 U629 ( .A1(n565), .A2(n564), .ZN(G299) );
  NAND2_X1 U630 ( .A1(G62), .A2(n792), .ZN(n567) );
  NAND2_X1 U631 ( .A1(G50), .A2(n796), .ZN(n566) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U633 ( .A(KEYINPUT82), .B(n568), .Z(n572) );
  NAND2_X1 U634 ( .A1(n793), .A2(G88), .ZN(n570) );
  NAND2_X1 U635 ( .A1(n797), .A2(G75), .ZN(n569) );
  AND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(G303) );
  INV_X1 U638 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U639 ( .A(G168), .B(KEYINPUT8), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n573), .B(KEYINPUT77), .ZN(G286) );
  NAND2_X1 U641 ( .A1(G49), .A2(n796), .ZN(n575) );
  NAND2_X1 U642 ( .A1(G74), .A2(G651), .ZN(n574) );
  NAND2_X1 U643 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U644 ( .A1(n792), .A2(n576), .ZN(n577) );
  XNOR2_X1 U645 ( .A(n577), .B(KEYINPUT80), .ZN(n580) );
  NAND2_X1 U646 ( .A1(G87), .A2(n578), .ZN(n579) );
  NAND2_X1 U647 ( .A1(n580), .A2(n579), .ZN(G288) );
  NAND2_X1 U648 ( .A1(G86), .A2(n793), .ZN(n582) );
  NAND2_X1 U649 ( .A1(n792), .A2(G61), .ZN(n581) );
  NAND2_X1 U650 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U651 ( .A(KEYINPUT81), .B(n583), .Z(n586) );
  NAND2_X1 U652 ( .A1(n797), .A2(G73), .ZN(n584) );
  XOR2_X1 U653 ( .A(KEYINPUT2), .B(n584), .Z(n585) );
  NOR2_X1 U654 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U655 ( .A1(n796), .A2(G48), .ZN(n587) );
  NAND2_X1 U656 ( .A1(n588), .A2(n587), .ZN(G305) );
  NAND2_X1 U657 ( .A1(G60), .A2(n792), .ZN(n590) );
  NAND2_X1 U658 ( .A1(G47), .A2(n796), .ZN(n589) );
  NAND2_X1 U659 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U660 ( .A(KEYINPUT70), .B(n591), .ZN(n594) );
  NAND2_X1 U661 ( .A1(G72), .A2(n797), .ZN(n592) );
  XNOR2_X1 U662 ( .A(KEYINPUT69), .B(n592), .ZN(n593) );
  NOR2_X1 U663 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X1 U664 ( .A1(G85), .A2(n793), .ZN(n595) );
  NAND2_X1 U665 ( .A1(n596), .A2(n595), .ZN(G290) );
  NOR2_X1 U666 ( .A1(G164), .A2(G1384), .ZN(n736) );
  NAND2_X1 U667 ( .A1(G160), .A2(G40), .ZN(n735) );
  INV_X1 U668 ( .A(n735), .ZN(n597) );
  NAND2_X2 U669 ( .A1(n736), .A2(n597), .ZN(n661) );
  AND2_X1 U670 ( .A1(G8), .A2(n661), .ZN(n711) );
  INV_X1 U671 ( .A(n711), .ZN(n705) );
  INV_X1 U672 ( .A(G1966), .ZN(n598) );
  AND2_X1 U673 ( .A1(n598), .A2(G8), .ZN(n599) );
  AND2_X1 U674 ( .A1(n661), .A2(n599), .ZN(n675) );
  NOR2_X1 U675 ( .A1(G2084), .A2(n661), .ZN(n674) );
  NOR2_X1 U676 ( .A1(n675), .A2(n674), .ZN(n600) );
  NAND2_X1 U677 ( .A1(G8), .A2(n600), .ZN(n603) );
  NOR2_X1 U678 ( .A1(G168), .A2(n604), .ZN(n606) );
  XNOR2_X1 U679 ( .A(n606), .B(n605), .ZN(n611) );
  XNOR2_X1 U680 ( .A(G2078), .B(KEYINPUT25), .ZN(n919) );
  NAND2_X1 U681 ( .A1(n648), .A2(n919), .ZN(n607) );
  XNOR2_X1 U682 ( .A(n607), .B(KEYINPUT89), .ZN(n609) );
  NOR2_X1 U683 ( .A1(n648), .A2(G1961), .ZN(n608) );
  NOR2_X1 U684 ( .A1(n609), .A2(n608), .ZN(n615) );
  NAND2_X1 U685 ( .A1(G301), .A2(n615), .ZN(n610) );
  NAND2_X1 U686 ( .A1(n611), .A2(n610), .ZN(n614) );
  INV_X1 U687 ( .A(KEYINPUT93), .ZN(n612) );
  NOR2_X1 U688 ( .A1(n615), .A2(G301), .ZN(n616) );
  XOR2_X1 U689 ( .A(KEYINPUT90), .B(n616), .Z(n660) );
  NAND2_X1 U690 ( .A1(G66), .A2(n792), .ZN(n618) );
  NAND2_X1 U691 ( .A1(G92), .A2(n793), .ZN(n617) );
  NAND2_X1 U692 ( .A1(n618), .A2(n617), .ZN(n623) );
  NAND2_X1 U693 ( .A1(n796), .A2(G54), .ZN(n620) );
  NAND2_X1 U694 ( .A1(G79), .A2(n797), .ZN(n619) );
  NAND2_X1 U695 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U696 ( .A(KEYINPUT76), .B(n621), .ZN(n622) );
  NOR2_X1 U697 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U698 ( .A(n624), .B(KEYINPUT15), .ZN(n775) );
  NAND2_X1 U699 ( .A1(G1348), .A2(n661), .ZN(n626) );
  NAND2_X1 U700 ( .A1(G2067), .A2(n648), .ZN(n625) );
  NAND2_X1 U701 ( .A1(n626), .A2(n625), .ZN(n645) );
  NOR2_X1 U702 ( .A1(n775), .A2(n645), .ZN(n644) );
  INV_X1 U703 ( .A(G1996), .ZN(n920) );
  NOR2_X1 U704 ( .A1(n661), .A2(n920), .ZN(n627) );
  XOR2_X1 U705 ( .A(n627), .B(KEYINPUT26), .Z(n629) );
  NAND2_X1 U706 ( .A1(n661), .A2(G1341), .ZN(n628) );
  NAND2_X1 U707 ( .A1(n629), .A2(n628), .ZN(n642) );
  NAND2_X1 U708 ( .A1(G56), .A2(n792), .ZN(n630) );
  XOR2_X1 U709 ( .A(KEYINPUT14), .B(n630), .Z(n639) );
  NAND2_X1 U710 ( .A1(G68), .A2(n797), .ZN(n635) );
  XOR2_X1 U711 ( .A(KEYINPUT12), .B(KEYINPUT74), .Z(n632) );
  NAND2_X1 U712 ( .A1(G81), .A2(n793), .ZN(n631) );
  XNOR2_X1 U713 ( .A(n632), .B(n631), .ZN(n633) );
  XNOR2_X1 U714 ( .A(KEYINPUT73), .B(n633), .ZN(n634) );
  NAND2_X1 U715 ( .A1(n635), .A2(n634), .ZN(n637) );
  XNOR2_X1 U716 ( .A(n637), .B(n636), .ZN(n638) );
  NOR2_X1 U717 ( .A1(n639), .A2(n638), .ZN(n641) );
  NAND2_X1 U718 ( .A1(n796), .A2(G43), .ZN(n640) );
  NOR2_X1 U719 ( .A1(n642), .A2(n946), .ZN(n643) );
  NOR2_X1 U720 ( .A1(n644), .A2(n643), .ZN(n647) );
  AND2_X1 U721 ( .A1(n775), .A2(n645), .ZN(n646) );
  NOR2_X1 U722 ( .A1(n647), .A2(n646), .ZN(n653) );
  NAND2_X1 U723 ( .A1(n648), .A2(G2072), .ZN(n649) );
  XOR2_X1 U724 ( .A(KEYINPUT27), .B(n649), .Z(n651) );
  NAND2_X1 U725 ( .A1(G1956), .A2(n661), .ZN(n650) );
  NAND2_X1 U726 ( .A1(n651), .A2(n650), .ZN(n654) );
  NOR2_X1 U727 ( .A1(G299), .A2(n654), .ZN(n652) );
  NOR2_X1 U728 ( .A1(n653), .A2(n652), .ZN(n657) );
  NAND2_X1 U729 ( .A1(G299), .A2(n654), .ZN(n655) );
  XOR2_X1 U730 ( .A(KEYINPUT28), .B(n655), .Z(n656) );
  NOR2_X1 U731 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U732 ( .A(KEYINPUT29), .B(n658), .ZN(n659) );
  NAND2_X1 U733 ( .A1(n660), .A2(n659), .ZN(n676) );
  NOR2_X1 U734 ( .A1(G1971), .A2(n705), .ZN(n663) );
  NOR2_X1 U735 ( .A1(G2090), .A2(n661), .ZN(n662) );
  NOR2_X1 U736 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U737 ( .A(KEYINPUT94), .B(n664), .Z(n665) );
  NOR2_X1 U738 ( .A1(G166), .A2(n665), .ZN(n666) );
  XNOR2_X1 U739 ( .A(n666), .B(KEYINPUT95), .ZN(n668) );
  AND2_X1 U740 ( .A1(n676), .A2(n668), .ZN(n667) );
  NAND2_X1 U741 ( .A1(n677), .A2(n667), .ZN(n672) );
  INV_X1 U742 ( .A(n668), .ZN(n669) );
  OR2_X1 U743 ( .A1(n669), .A2(G286), .ZN(n670) );
  AND2_X1 U744 ( .A1(n670), .A2(G8), .ZN(n671) );
  NAND2_X1 U745 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U746 ( .A(n673), .B(KEYINPUT32), .ZN(n682) );
  NAND2_X1 U747 ( .A1(G8), .A2(n674), .ZN(n680) );
  AND2_X1 U748 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U749 ( .A1(n675), .A2(n678), .ZN(n679) );
  NAND2_X1 U750 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U751 ( .A1(n682), .A2(n681), .ZN(n704) );
  NOR2_X1 U752 ( .A1(G1971), .A2(G303), .ZN(n683) );
  NOR2_X1 U753 ( .A1(G1976), .A2(G288), .ZN(n943) );
  NOR2_X1 U754 ( .A1(n683), .A2(n943), .ZN(n684) );
  NAND2_X1 U755 ( .A1(n704), .A2(n684), .ZN(n685) );
  NAND2_X1 U756 ( .A1(G1976), .A2(G288), .ZN(n950) );
  NAND2_X1 U757 ( .A1(n685), .A2(n950), .ZN(n690) );
  NOR2_X1 U758 ( .A1(n705), .A2(n690), .ZN(n686) );
  NOR2_X1 U759 ( .A1(n686), .A2(KEYINPUT33), .ZN(n687) );
  NAND2_X1 U760 ( .A1(n687), .A2(KEYINPUT96), .ZN(n688) );
  NAND2_X1 U761 ( .A1(G1981), .A2(G305), .ZN(n957) );
  NAND2_X1 U762 ( .A1(n688), .A2(n957), .ZN(n695) );
  NAND2_X1 U763 ( .A1(n943), .A2(KEYINPUT33), .ZN(n689) );
  XNOR2_X1 U764 ( .A(n689), .B(KEYINPUT97), .ZN(n692) );
  NOR2_X1 U765 ( .A1(n690), .A2(KEYINPUT96), .ZN(n691) );
  NOR2_X1 U766 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U767 ( .A1(n693), .A2(n705), .ZN(n694) );
  NOR2_X1 U768 ( .A1(G1981), .A2(G305), .ZN(n960) );
  INV_X1 U769 ( .A(KEYINPUT33), .ZN(n696) );
  NOR2_X1 U770 ( .A1(KEYINPUT96), .A2(n696), .ZN(n697) );
  NOR2_X1 U771 ( .A1(n960), .A2(n697), .ZN(n698) );
  NAND2_X1 U772 ( .A1(n699), .A2(n698), .ZN(n708) );
  NOR2_X1 U773 ( .A1(G2090), .A2(G303), .ZN(n700) );
  XNOR2_X1 U774 ( .A(KEYINPUT98), .B(n700), .ZN(n701) );
  NAND2_X1 U775 ( .A1(n701), .A2(G8), .ZN(n702) );
  XOR2_X1 U776 ( .A(KEYINPUT99), .B(n702), .Z(n703) );
  NAND2_X1 U777 ( .A1(n704), .A2(n703), .ZN(n706) );
  NAND2_X1 U778 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U779 ( .A1(n708), .A2(n707), .ZN(n710) );
  XNOR2_X1 U780 ( .A(n960), .B(KEYINPUT24), .ZN(n712) );
  NAND2_X1 U781 ( .A1(n712), .A2(n711), .ZN(n738) );
  NAND2_X1 U782 ( .A1(G117), .A2(n898), .ZN(n714) );
  NAND2_X1 U783 ( .A1(G129), .A2(n895), .ZN(n713) );
  NAND2_X1 U784 ( .A1(n714), .A2(n713), .ZN(n720) );
  NAND2_X1 U785 ( .A1(G105), .A2(n715), .ZN(n716) );
  XNOR2_X1 U786 ( .A(n716), .B(KEYINPUT38), .ZN(n718) );
  NAND2_X1 U787 ( .A1(G141), .A2(n889), .ZN(n717) );
  NAND2_X1 U788 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U789 ( .A1(n720), .A2(n719), .ZN(n871) );
  AND2_X1 U790 ( .A1(n920), .A2(n871), .ZN(n1005) );
  NAND2_X1 U791 ( .A1(G131), .A2(n889), .ZN(n722) );
  NAND2_X1 U792 ( .A1(G119), .A2(n895), .ZN(n721) );
  NAND2_X1 U793 ( .A1(n722), .A2(n721), .ZN(n726) );
  NAND2_X1 U794 ( .A1(n898), .A2(G107), .ZN(n724) );
  NAND2_X1 U795 ( .A1(G95), .A2(n715), .ZN(n723) );
  NAND2_X1 U796 ( .A1(n724), .A2(n723), .ZN(n725) );
  OR2_X1 U797 ( .A1(n726), .A2(n725), .ZN(n884) );
  NAND2_X1 U798 ( .A1(G1991), .A2(n884), .ZN(n727) );
  XOR2_X1 U799 ( .A(KEYINPUT88), .B(n727), .Z(n729) );
  NOR2_X1 U800 ( .A1(n871), .A2(n920), .ZN(n728) );
  NOR2_X1 U801 ( .A1(n729), .A2(n728), .ZN(n754) );
  INV_X1 U802 ( .A(n754), .ZN(n1012) );
  NOR2_X1 U803 ( .A1(G1986), .A2(G290), .ZN(n730) );
  NOR2_X1 U804 ( .A1(G1991), .A2(n884), .ZN(n1003) );
  NOR2_X1 U805 ( .A1(n730), .A2(n1003), .ZN(n731) );
  NOR2_X1 U806 ( .A1(n1012), .A2(n731), .ZN(n732) );
  NOR2_X1 U807 ( .A1(n1005), .A2(n732), .ZN(n733) );
  XOR2_X1 U808 ( .A(n733), .B(KEYINPUT101), .Z(n734) );
  XNOR2_X1 U809 ( .A(KEYINPUT39), .B(n734), .ZN(n737) );
  NOR2_X1 U810 ( .A1(n736), .A2(n735), .ZN(n763) );
  NAND2_X1 U811 ( .A1(n737), .A2(n763), .ZN(n753) );
  AND2_X1 U812 ( .A1(n738), .A2(n753), .ZN(n739) );
  NAND2_X1 U813 ( .A1(n740), .A2(n739), .ZN(n761) );
  NAND2_X1 U814 ( .A1(G104), .A2(n715), .ZN(n741) );
  XOR2_X1 U815 ( .A(KEYINPUT85), .B(n741), .Z(n743) );
  NAND2_X1 U816 ( .A1(n889), .A2(G140), .ZN(n742) );
  NAND2_X1 U817 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U818 ( .A(KEYINPUT34), .B(n744), .ZN(n751) );
  NAND2_X1 U819 ( .A1(n898), .A2(G116), .ZN(n745) );
  XNOR2_X1 U820 ( .A(n745), .B(KEYINPUT86), .ZN(n747) );
  NAND2_X1 U821 ( .A1(G128), .A2(n895), .ZN(n746) );
  NAND2_X1 U822 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U823 ( .A(KEYINPUT35), .B(n748), .ZN(n749) );
  XNOR2_X1 U824 ( .A(KEYINPUT87), .B(n749), .ZN(n750) );
  NOR2_X1 U825 ( .A1(n751), .A2(n750), .ZN(n752) );
  XOR2_X1 U826 ( .A(KEYINPUT36), .B(n752), .Z(n903) );
  XOR2_X1 U827 ( .A(KEYINPUT37), .B(G2067), .Z(n762) );
  AND2_X1 U828 ( .A1(n903), .A2(n762), .ZN(n1018) );
  NAND2_X1 U829 ( .A1(n1018), .A2(n763), .ZN(n759) );
  INV_X1 U830 ( .A(n753), .ZN(n757) );
  XOR2_X1 U831 ( .A(G1986), .B(G290), .Z(n944) );
  NAND2_X1 U832 ( .A1(n754), .A2(n944), .ZN(n755) );
  NAND2_X1 U833 ( .A1(n755), .A2(n763), .ZN(n756) );
  OR2_X1 U834 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U835 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U836 ( .A1(n761), .A2(n760), .ZN(n765) );
  NOR2_X1 U837 ( .A1(n903), .A2(n762), .ZN(n1022) );
  NAND2_X1 U838 ( .A1(n1022), .A2(n763), .ZN(n764) );
  NAND2_X1 U839 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U840 ( .A(n766), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U841 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U842 ( .A(G57), .ZN(G237) );
  INV_X1 U843 ( .A(G132), .ZN(G219) );
  NAND2_X1 U844 ( .A1(G7), .A2(G661), .ZN(n767) );
  XNOR2_X1 U845 ( .A(n767), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U846 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n769) );
  INV_X1 U847 ( .A(G223), .ZN(n837) );
  NAND2_X1 U848 ( .A1(G567), .A2(n837), .ZN(n768) );
  XNOR2_X1 U849 ( .A(n769), .B(n768), .ZN(G234) );
  XNOR2_X1 U850 ( .A(G860), .B(KEYINPUT75), .ZN(n774) );
  OR2_X1 U851 ( .A1(n946), .A2(n774), .ZN(G153) );
  NAND2_X1 U852 ( .A1(G868), .A2(G301), .ZN(n771) );
  INV_X1 U853 ( .A(G868), .ZN(n811) );
  NAND2_X1 U854 ( .A1(n775), .A2(n811), .ZN(n770) );
  NAND2_X1 U855 ( .A1(n771), .A2(n770), .ZN(G284) );
  NOR2_X1 U856 ( .A1(G286), .A2(n811), .ZN(n773) );
  NOR2_X1 U857 ( .A1(G868), .A2(G299), .ZN(n772) );
  NOR2_X1 U858 ( .A1(n773), .A2(n772), .ZN(G297) );
  NAND2_X1 U859 ( .A1(n774), .A2(G559), .ZN(n776) );
  INV_X1 U860 ( .A(n775), .ZN(n963) );
  NAND2_X1 U861 ( .A1(n776), .A2(n963), .ZN(n777) );
  XNOR2_X1 U862 ( .A(n777), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U863 ( .A1(n963), .A2(G868), .ZN(n778) );
  NOR2_X1 U864 ( .A1(G559), .A2(n778), .ZN(n779) );
  XNOR2_X1 U865 ( .A(n779), .B(KEYINPUT78), .ZN(n781) );
  NOR2_X1 U866 ( .A1(n946), .A2(G868), .ZN(n780) );
  NOR2_X1 U867 ( .A1(n781), .A2(n780), .ZN(G282) );
  NAND2_X1 U868 ( .A1(G123), .A2(n895), .ZN(n782) );
  XNOR2_X1 U869 ( .A(n782), .B(KEYINPUT18), .ZN(n784) );
  NAND2_X1 U870 ( .A1(n898), .A2(G111), .ZN(n783) );
  NAND2_X1 U871 ( .A1(n784), .A2(n783), .ZN(n788) );
  NAND2_X1 U872 ( .A1(n889), .A2(G135), .ZN(n786) );
  NAND2_X1 U873 ( .A1(G99), .A2(n715), .ZN(n785) );
  NAND2_X1 U874 ( .A1(n786), .A2(n785), .ZN(n787) );
  NOR2_X1 U875 ( .A1(n788), .A2(n787), .ZN(n1002) );
  XOR2_X1 U876 ( .A(G2096), .B(n1002), .Z(n789) );
  NOR2_X1 U877 ( .A1(G2100), .A2(n789), .ZN(n790) );
  XNOR2_X1 U878 ( .A(KEYINPUT79), .B(n790), .ZN(G156) );
  NAND2_X1 U879 ( .A1(n963), .A2(G559), .ZN(n809) );
  XNOR2_X1 U880 ( .A(n946), .B(n809), .ZN(n791) );
  NOR2_X1 U881 ( .A1(n791), .A2(G860), .ZN(n802) );
  NAND2_X1 U882 ( .A1(G67), .A2(n792), .ZN(n795) );
  NAND2_X1 U883 ( .A1(G93), .A2(n793), .ZN(n794) );
  NAND2_X1 U884 ( .A1(n795), .A2(n794), .ZN(n801) );
  NAND2_X1 U885 ( .A1(n796), .A2(G55), .ZN(n799) );
  NAND2_X1 U886 ( .A1(G80), .A2(n797), .ZN(n798) );
  NAND2_X1 U887 ( .A1(n799), .A2(n798), .ZN(n800) );
  OR2_X1 U888 ( .A1(n801), .A2(n800), .ZN(n812) );
  XOR2_X1 U889 ( .A(n802), .B(n812), .Z(G145) );
  XNOR2_X1 U890 ( .A(KEYINPUT19), .B(G299), .ZN(n803) );
  XNOR2_X1 U891 ( .A(n803), .B(G290), .ZN(n806) );
  XOR2_X1 U892 ( .A(n812), .B(n946), .Z(n804) );
  XNOR2_X1 U893 ( .A(n804), .B(G288), .ZN(n805) );
  XNOR2_X1 U894 ( .A(n806), .B(n805), .ZN(n808) );
  XNOR2_X1 U895 ( .A(G305), .B(G166), .ZN(n807) );
  XNOR2_X1 U896 ( .A(n808), .B(n807), .ZN(n908) );
  XOR2_X1 U897 ( .A(n908), .B(n809), .Z(n810) );
  NAND2_X1 U898 ( .A1(G868), .A2(n810), .ZN(n814) );
  NAND2_X1 U899 ( .A1(n812), .A2(n811), .ZN(n813) );
  NAND2_X1 U900 ( .A1(n814), .A2(n813), .ZN(G295) );
  NAND2_X1 U901 ( .A1(G2078), .A2(G2084), .ZN(n815) );
  XOR2_X1 U902 ( .A(KEYINPUT20), .B(n815), .Z(n816) );
  NAND2_X1 U903 ( .A1(G2090), .A2(n816), .ZN(n817) );
  XNOR2_X1 U904 ( .A(KEYINPUT21), .B(n817), .ZN(n818) );
  NAND2_X1 U905 ( .A1(n818), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U906 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U907 ( .A(KEYINPUT71), .B(G82), .ZN(G220) );
  NOR2_X1 U908 ( .A1(G219), .A2(G220), .ZN(n819) );
  XOR2_X1 U909 ( .A(KEYINPUT22), .B(n819), .Z(n820) );
  NOR2_X1 U910 ( .A1(G218), .A2(n820), .ZN(n821) );
  NAND2_X1 U911 ( .A1(G96), .A2(n821), .ZN(n842) );
  NAND2_X1 U912 ( .A1(n842), .A2(G2106), .ZN(n825) );
  NAND2_X1 U913 ( .A1(G120), .A2(G69), .ZN(n822) );
  NOR2_X1 U914 ( .A1(G237), .A2(n822), .ZN(n823) );
  NAND2_X1 U915 ( .A1(G108), .A2(n823), .ZN(n841) );
  NAND2_X1 U916 ( .A1(n841), .A2(G567), .ZN(n824) );
  NAND2_X1 U917 ( .A1(n825), .A2(n824), .ZN(n844) );
  NAND2_X1 U918 ( .A1(G483), .A2(G661), .ZN(n826) );
  NOR2_X1 U919 ( .A1(n844), .A2(n826), .ZN(n840) );
  NAND2_X1 U920 ( .A1(n840), .A2(G36), .ZN(G176) );
  XNOR2_X1 U921 ( .A(G2454), .B(G2451), .ZN(n835) );
  XNOR2_X1 U922 ( .A(G2430), .B(G2446), .ZN(n833) );
  XOR2_X1 U923 ( .A(G2435), .B(G2427), .Z(n828) );
  XNOR2_X1 U924 ( .A(KEYINPUT102), .B(G2438), .ZN(n827) );
  XNOR2_X1 U925 ( .A(n828), .B(n827), .ZN(n829) );
  XOR2_X1 U926 ( .A(n829), .B(G2443), .Z(n831) );
  XNOR2_X1 U927 ( .A(G1341), .B(G1348), .ZN(n830) );
  XNOR2_X1 U928 ( .A(n831), .B(n830), .ZN(n832) );
  XNOR2_X1 U929 ( .A(n833), .B(n832), .ZN(n834) );
  XNOR2_X1 U930 ( .A(n835), .B(n834), .ZN(n836) );
  NAND2_X1 U931 ( .A1(n836), .A2(G14), .ZN(n912) );
  XNOR2_X1 U932 ( .A(KEYINPUT103), .B(n912), .ZN(G401) );
  NAND2_X1 U933 ( .A1(G2106), .A2(n837), .ZN(G217) );
  AND2_X1 U934 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U935 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U936 ( .A1(G3), .A2(G1), .ZN(n839) );
  NAND2_X1 U937 ( .A1(n840), .A2(n839), .ZN(G188) );
  XOR2_X1 U938 ( .A(G69), .B(KEYINPUT104), .Z(G235) );
  INV_X1 U940 ( .A(G120), .ZN(G236) );
  INV_X1 U941 ( .A(G96), .ZN(G221) );
  NOR2_X1 U942 ( .A1(n842), .A2(n841), .ZN(n843) );
  XNOR2_X1 U943 ( .A(n843), .B(KEYINPUT105), .ZN(G261) );
  INV_X1 U944 ( .A(G261), .ZN(G325) );
  INV_X1 U945 ( .A(n844), .ZN(G319) );
  XNOR2_X1 U946 ( .A(G1956), .B(G2474), .ZN(n854) );
  XOR2_X1 U947 ( .A(G1986), .B(G1971), .Z(n846) );
  XNOR2_X1 U948 ( .A(G1981), .B(G1966), .ZN(n845) );
  XNOR2_X1 U949 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U950 ( .A(G1991), .B(G1976), .Z(n848) );
  XNOR2_X1 U951 ( .A(G1996), .B(G1961), .ZN(n847) );
  XNOR2_X1 U952 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U953 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U954 ( .A(KEYINPUT106), .B(KEYINPUT41), .ZN(n851) );
  XNOR2_X1 U955 ( .A(n852), .B(n851), .ZN(n853) );
  XNOR2_X1 U956 ( .A(n854), .B(n853), .ZN(G229) );
  XOR2_X1 U957 ( .A(G2100), .B(G2096), .Z(n856) );
  XNOR2_X1 U958 ( .A(KEYINPUT42), .B(G2678), .ZN(n855) );
  XNOR2_X1 U959 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U960 ( .A(KEYINPUT43), .B(G2090), .Z(n858) );
  XNOR2_X1 U961 ( .A(G2067), .B(G2072), .ZN(n857) );
  XNOR2_X1 U962 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U963 ( .A(n860), .B(n859), .Z(n862) );
  XNOR2_X1 U964 ( .A(G2078), .B(G2084), .ZN(n861) );
  XNOR2_X1 U965 ( .A(n862), .B(n861), .ZN(G227) );
  NAND2_X1 U966 ( .A1(G124), .A2(n895), .ZN(n863) );
  XNOR2_X1 U967 ( .A(n863), .B(KEYINPUT44), .ZN(n866) );
  NAND2_X1 U968 ( .A1(G136), .A2(n889), .ZN(n864) );
  XOR2_X1 U969 ( .A(KEYINPUT107), .B(n864), .Z(n865) );
  NAND2_X1 U970 ( .A1(n866), .A2(n865), .ZN(n870) );
  NAND2_X1 U971 ( .A1(n898), .A2(G112), .ZN(n868) );
  NAND2_X1 U972 ( .A1(G100), .A2(n715), .ZN(n867) );
  NAND2_X1 U973 ( .A1(n868), .A2(n867), .ZN(n869) );
  NOR2_X1 U974 ( .A1(n870), .A2(n869), .ZN(G162) );
  XOR2_X1 U975 ( .A(G162), .B(n871), .Z(n873) );
  XNOR2_X1 U976 ( .A(G164), .B(G160), .ZN(n872) );
  XNOR2_X1 U977 ( .A(n873), .B(n872), .ZN(n888) );
  XOR2_X1 U978 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n875) );
  XNOR2_X1 U979 ( .A(KEYINPUT112), .B(KEYINPUT111), .ZN(n874) );
  XNOR2_X1 U980 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U981 ( .A(n1002), .B(n876), .ZN(n886) );
  NAND2_X1 U982 ( .A1(n889), .A2(G139), .ZN(n878) );
  NAND2_X1 U983 ( .A1(G103), .A2(n715), .ZN(n877) );
  NAND2_X1 U984 ( .A1(n878), .A2(n877), .ZN(n883) );
  NAND2_X1 U985 ( .A1(G115), .A2(n898), .ZN(n880) );
  NAND2_X1 U986 ( .A1(G127), .A2(n895), .ZN(n879) );
  NAND2_X1 U987 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U988 ( .A(KEYINPUT47), .B(n881), .Z(n882) );
  NOR2_X1 U989 ( .A1(n883), .A2(n882), .ZN(n1013) );
  XNOR2_X1 U990 ( .A(n884), .B(n1013), .ZN(n885) );
  XNOR2_X1 U991 ( .A(n886), .B(n885), .ZN(n887) );
  XOR2_X1 U992 ( .A(n888), .B(n887), .Z(n905) );
  NAND2_X1 U993 ( .A1(n889), .A2(G142), .ZN(n890) );
  XNOR2_X1 U994 ( .A(KEYINPUT110), .B(n890), .ZN(n893) );
  NAND2_X1 U995 ( .A1(G106), .A2(n715), .ZN(n891) );
  XOR2_X1 U996 ( .A(KEYINPUT109), .B(n891), .Z(n892) );
  NAND2_X1 U997 ( .A1(n893), .A2(n892), .ZN(n894) );
  XNOR2_X1 U998 ( .A(n894), .B(KEYINPUT45), .ZN(n897) );
  NAND2_X1 U999 ( .A1(G130), .A2(n895), .ZN(n896) );
  NAND2_X1 U1000 ( .A1(n897), .A2(n896), .ZN(n901) );
  NAND2_X1 U1001 ( .A1(n898), .A2(G118), .ZN(n899) );
  XOR2_X1 U1002 ( .A(KEYINPUT108), .B(n899), .Z(n900) );
  NOR2_X1 U1003 ( .A1(n901), .A2(n900), .ZN(n902) );
  XNOR2_X1 U1004 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U1005 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n906), .ZN(n907) );
  XOR2_X1 U1007 ( .A(KEYINPUT113), .B(n907), .Z(G395) );
  XNOR2_X1 U1008 ( .A(G171), .B(G286), .ZN(n909) );
  XNOR2_X1 U1009 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1010 ( .A(n910), .B(n963), .ZN(n911) );
  NOR2_X1 U1011 ( .A1(G37), .A2(n911), .ZN(G397) );
  NAND2_X1 U1012 ( .A1(G319), .A2(n912), .ZN(n915) );
  NOR2_X1 U1013 ( .A1(G229), .A2(G227), .ZN(n913) );
  XNOR2_X1 U1014 ( .A(n913), .B(KEYINPUT49), .ZN(n914) );
  NOR2_X1 U1015 ( .A1(n915), .A2(n914), .ZN(n916) );
  XNOR2_X1 U1016 ( .A(KEYINPUT114), .B(n916), .ZN(n918) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1018 ( .A1(n918), .A2(n917), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1021 ( .A(KEYINPUT55), .B(KEYINPUT117), .Z(n938) );
  XNOR2_X1 U1022 ( .A(G2090), .B(G35), .ZN(n933) );
  XNOR2_X1 U1023 ( .A(G27), .B(n919), .ZN(n928) );
  XOR2_X1 U1024 ( .A(G2067), .B(G26), .Z(n922) );
  XNOR2_X1 U1025 ( .A(n920), .B(G32), .ZN(n921) );
  NAND2_X1 U1026 ( .A1(n922), .A2(n921), .ZN(n926) );
  XOR2_X1 U1027 ( .A(G1991), .B(G25), .Z(n923) );
  NAND2_X1 U1028 ( .A1(n923), .A2(G28), .ZN(n924) );
  XNOR2_X1 U1029 ( .A(KEYINPUT116), .B(n924), .ZN(n925) );
  NOR2_X1 U1030 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1031 ( .A1(n928), .A2(n927), .ZN(n930) );
  XNOR2_X1 U1032 ( .A(G33), .B(G2072), .ZN(n929) );
  NOR2_X1 U1033 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1034 ( .A(KEYINPUT53), .B(n931), .ZN(n932) );
  NOR2_X1 U1035 ( .A1(n933), .A2(n932), .ZN(n936) );
  XOR2_X1 U1036 ( .A(G2084), .B(G34), .Z(n934) );
  XNOR2_X1 U1037 ( .A(KEYINPUT54), .B(n934), .ZN(n935) );
  NAND2_X1 U1038 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1039 ( .A(n938), .B(n937), .ZN(n940) );
  XNOR2_X1 U1040 ( .A(KEYINPUT118), .B(G29), .ZN(n939) );
  NOR2_X1 U1041 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1042 ( .A(KEYINPUT119), .B(n941), .ZN(n942) );
  NAND2_X1 U1043 ( .A1(n942), .A2(G11), .ZN(n1001) );
  XNOR2_X1 U1044 ( .A(G16), .B(KEYINPUT56), .ZN(n971) );
  XNOR2_X1 U1045 ( .A(n943), .B(KEYINPUT123), .ZN(n945) );
  NAND2_X1 U1046 ( .A1(n945), .A2(n944), .ZN(n948) );
  XNOR2_X1 U1047 ( .A(G1341), .B(n946), .ZN(n947) );
  NOR2_X1 U1048 ( .A1(n948), .A2(n947), .ZN(n969) );
  XNOR2_X1 U1049 ( .A(G166), .B(G1971), .ZN(n956) );
  XOR2_X1 U1050 ( .A(G1956), .B(KEYINPUT122), .Z(n949) );
  XNOR2_X1 U1051 ( .A(G299), .B(n949), .ZN(n951) );
  NAND2_X1 U1052 ( .A1(n951), .A2(n950), .ZN(n954) );
  XOR2_X1 U1053 ( .A(G1961), .B(G301), .Z(n952) );
  XNOR2_X1 U1054 ( .A(KEYINPUT121), .B(n952), .ZN(n953) );
  NOR2_X1 U1055 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1056 ( .A1(n956), .A2(n955), .ZN(n967) );
  XNOR2_X1 U1057 ( .A(G1966), .B(G168), .ZN(n958) );
  NAND2_X1 U1058 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1059 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1060 ( .A(KEYINPUT120), .B(n961), .Z(n962) );
  XNOR2_X1 U1061 ( .A(KEYINPUT57), .B(n962), .ZN(n965) );
  XNOR2_X1 U1062 ( .A(n963), .B(G1348), .ZN(n964) );
  NAND2_X1 U1063 ( .A1(n965), .A2(n964), .ZN(n966) );
  NOR2_X1 U1064 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1065 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n999) );
  INV_X1 U1067 ( .A(G16), .ZN(n997) );
  XOR2_X1 U1068 ( .A(KEYINPUT125), .B(G4), .Z(n973) );
  XNOR2_X1 U1069 ( .A(G1348), .B(KEYINPUT59), .ZN(n972) );
  XNOR2_X1 U1070 ( .A(n973), .B(n972), .ZN(n977) );
  XNOR2_X1 U1071 ( .A(G1981), .B(G6), .ZN(n975) );
  XNOR2_X1 U1072 ( .A(G1956), .B(G20), .ZN(n974) );
  NOR2_X1 U1073 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1074 ( .A1(n977), .A2(n976), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(KEYINPUT124), .B(G1341), .ZN(n978) );
  XNOR2_X1 U1076 ( .A(G19), .B(n978), .ZN(n979) );
  NOR2_X1 U1077 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1078 ( .A(KEYINPUT126), .B(n981), .ZN(n982) );
  XNOR2_X1 U1079 ( .A(n982), .B(KEYINPUT60), .ZN(n986) );
  XNOR2_X1 U1080 ( .A(G1966), .B(G21), .ZN(n984) );
  XNOR2_X1 U1081 ( .A(G1961), .B(G5), .ZN(n983) );
  NOR2_X1 U1082 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1083 ( .A1(n986), .A2(n985), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(G1971), .B(G22), .ZN(n988) );
  XNOR2_X1 U1085 ( .A(G23), .B(G1976), .ZN(n987) );
  NOR2_X1 U1086 ( .A1(n988), .A2(n987), .ZN(n990) );
  XOR2_X1 U1087 ( .A(G1986), .B(G24), .Z(n989) );
  NAND2_X1 U1088 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1089 ( .A(KEYINPUT58), .B(n991), .ZN(n992) );
  NOR2_X1 U1090 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1091 ( .A(n994), .B(KEYINPUT127), .Z(n995) );
  XNOR2_X1 U1092 ( .A(KEYINPUT61), .B(n995), .ZN(n996) );
  NAND2_X1 U1093 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1094 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NOR2_X1 U1095 ( .A1(n1001), .A2(n1000), .ZN(n1029) );
  NOR2_X1 U1096 ( .A1(n1003), .A2(n1002), .ZN(n1010) );
  XOR2_X1 U1097 ( .A(G160), .B(G2084), .Z(n1008) );
  XOR2_X1 U1098 ( .A(G2090), .B(G162), .Z(n1004) );
  NOR2_X1 U1099 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1100 ( .A(KEYINPUT51), .B(n1006), .ZN(n1007) );
  NOR2_X1 U1101 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1102 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1103 ( .A1(n1012), .A2(n1011), .ZN(n1020) );
  XOR2_X1 U1104 ( .A(G2072), .B(n1013), .Z(n1015) );
  XOR2_X1 U1105 ( .A(G164), .B(G2078), .Z(n1014) );
  NOR2_X1 U1106 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1107 ( .A(KEYINPUT50), .B(n1016), .Z(n1017) );
  NOR2_X1 U1108 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1109 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1111 ( .A(KEYINPUT52), .B(n1023), .Z(n1024) );
  NOR2_X1 U1112 ( .A1(KEYINPUT55), .A2(n1024), .ZN(n1026) );
  INV_X1 U1113 ( .A(G29), .ZN(n1025) );
  NOR2_X1 U1114 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1115 ( .A(n1027), .B(KEYINPUT115), .ZN(n1028) );
  NAND2_X1 U1116 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1117 ( .A(KEYINPUT62), .B(n1030), .Z(G311) );
  INV_X1 U1118 ( .A(G311), .ZN(G150) );
endmodule

