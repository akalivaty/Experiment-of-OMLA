//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 0 0 0 1 0 1 1 1 1 0 0 1 0 1 0 0 0 1 1 0 0 0 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 0 0 1 1 0 0 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n557,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n611,
    new_n612, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1138, new_n1139;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT66), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  AND2_X1   g017(.A1(G2072), .A2(G2078), .ZN(new_n443));
  NAND3_X1  g018(.A1(new_n443), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI211_X1 g039(.A(G137), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n466), .B1(new_n468), .B2(G101), .ZN(new_n469));
  AND4_X1   g044(.A1(new_n466), .A2(new_n462), .A3(G101), .A4(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n465), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g046(.A(G125), .B1(new_n463), .B2(new_n464), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n462), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n471), .A2(new_n474), .ZN(G160));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(new_n467), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n479), .A2(new_n462), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  MUX2_X1   g060(.A(G100), .B(G112), .S(G2105), .Z(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2104), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n482), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  INV_X1    g064(.A(G126), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n490), .B1(new_n477), .B2(new_n478), .ZN(new_n491));
  AND2_X1   g066(.A1(G114), .A2(G2104), .ZN(new_n492));
  OAI21_X1  g067(.A(G2105), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(KEYINPUT4), .A2(G138), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n494), .B1(new_n477), .B2(new_n478), .ZN(new_n495));
  NAND2_X1  g070(.A1(G102), .A2(G2104), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n462), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  OAI211_X1 g073(.A(G138), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n493), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT68), .ZN(new_n503));
  AND2_X1   g078(.A1(KEYINPUT4), .A2(G138), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n504), .B1(new_n463), .B2(new_n464), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(new_n496), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(new_n462), .B1(new_n500), .B2(new_n499), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT68), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n507), .A2(new_n508), .A3(new_n493), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(G164));
  XNOR2_X1  g086(.A(KEYINPUT5), .B(G543), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT6), .B(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G50), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n514), .A2(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n518), .A2(new_n521), .ZN(G166));
  XNOR2_X1  g097(.A(KEYINPUT69), .B(G89), .ZN(new_n523));
  INV_X1    g098(.A(G51), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n514), .A2(new_n523), .B1(new_n516), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n525), .A2(new_n529), .ZN(G168));
  INV_X1    g105(.A(new_n514), .ZN(new_n531));
  INV_X1    g106(.A(new_n516), .ZN(new_n532));
  AOI22_X1  g107(.A1(G90), .A2(new_n531), .B1(new_n532), .B2(G52), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT71), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n533), .B(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(new_n512), .ZN(new_n537));
  INV_X1    g112(.A(G64), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT70), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n520), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n541), .B1(new_n540), .B2(new_n539), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n535), .A2(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  INV_X1    g120(.A(G43), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n514), .A2(new_n545), .B1(new_n516), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT73), .ZN(new_n548));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G56), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n537), .B2(new_n550), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n520), .B1(new_n551), .B2(KEYINPUT72), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n552), .B1(KEYINPUT72), .B2(new_n551), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(G188));
  NAND3_X1  g136(.A1(new_n513), .A2(G53), .A3(G543), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT9), .ZN(new_n563));
  OR2_X1    g138(.A1(new_n563), .A2(KEYINPUT74), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(KEYINPUT74), .ZN(new_n565));
  INV_X1    g140(.A(G91), .ZN(new_n566));
  OR3_X1    g141(.A1(new_n514), .A2(KEYINPUT75), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT75), .B1(new_n514), .B2(new_n566), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n537), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n567), .A2(new_n568), .B1(G651), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n564), .A2(new_n565), .A3(new_n572), .ZN(G299));
  INV_X1    g148(.A(G168), .ZN(G286));
  INV_X1    g149(.A(G166), .ZN(G303));
  NAND2_X1  g150(.A1(new_n531), .A2(G87), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n532), .A2(G49), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(G288));
  NAND3_X1  g154(.A1(new_n513), .A2(G48), .A3(G543), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT77), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n513), .A2(KEYINPUT77), .A3(G48), .A4(G543), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n512), .A2(new_n513), .A3(G86), .ZN(new_n584));
  AND3_X1   g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n512), .A2(G61), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n520), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n588), .A2(KEYINPUT76), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT76), .ZN(new_n590));
  AOI211_X1 g165(.A(new_n590), .B(new_n520), .C1(new_n586), .C2(new_n587), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n585), .B1(new_n589), .B2(new_n591), .ZN(G305));
  INV_X1    g167(.A(G85), .ZN(new_n593));
  INV_X1    g168(.A(G47), .ZN(new_n594));
  OAI22_X1  g169(.A1(new_n514), .A2(new_n593), .B1(new_n516), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n596), .A2(new_n520), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(new_n531), .A2(G92), .ZN(new_n600));
  XOR2_X1   g175(.A(new_n600), .B(KEYINPUT10), .Z(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n537), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n604), .A2(G651), .B1(new_n532), .B2(G54), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  MUX2_X1   g181(.A(new_n606), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g182(.A(new_n606), .B(G301), .S(G868), .Z(G321));
  MUX2_X1   g183(.A(G299), .B(G286), .S(G868), .Z(G297));
  XNOR2_X1  g184(.A(G297), .B(KEYINPUT78), .ZN(G280));
  INV_X1    g185(.A(new_n606), .ZN(new_n611));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(G860), .ZN(G148));
  NAND2_X1  g188(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  MUX2_X1   g189(.A(new_n554), .B(new_n614), .S(G868), .Z(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g191(.A1(new_n483), .A2(new_n467), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT12), .ZN(new_n618));
  XNOR2_X1  g193(.A(KEYINPUT79), .B(KEYINPUT13), .ZN(new_n619));
  AND2_X1   g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n618), .A2(new_n619), .ZN(new_n621));
  OAI22_X1  g196(.A1(new_n620), .A2(new_n621), .B1(KEYINPUT80), .B2(G2100), .ZN(new_n622));
  NAND2_X1  g197(.A1(KEYINPUT80), .A2(G2100), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  MUX2_X1   g200(.A(G99), .B(G111), .S(G2105), .Z(new_n626));
  AOI22_X1  g201(.A1(new_n481), .A2(G123), .B1(G2104), .B2(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(G135), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(new_n483), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(G2096), .Z(new_n630));
  NAND3_X1  g205(.A1(new_n624), .A2(new_n625), .A3(new_n630), .ZN(G156));
  XNOR2_X1  g206(.A(G2443), .B(G2446), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT82), .ZN(new_n633));
  XOR2_X1   g208(.A(G2451), .B(G2454), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(KEYINPUT14), .ZN(new_n640));
  XOR2_X1   g215(.A(KEYINPUT15), .B(G2435), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2427), .ZN(new_n643));
  INV_X1    g218(.A(G2430), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n640), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(new_n644), .B2(new_n643), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n639), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n639), .A2(new_n646), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(G14), .A3(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(G401));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT83), .Z(new_n652));
  NOR2_X1   g227(.A1(G2072), .A2(G2078), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n443), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n654), .B(KEYINPUT17), .ZN(new_n658));
  OAI211_X1 g233(.A(new_n655), .B(new_n657), .C1(new_n652), .C2(new_n658), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n652), .A2(new_n658), .A3(new_n656), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n656), .B(new_n651), .C1(new_n443), .C2(new_n653), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT18), .Z(new_n662));
  NAND3_X1  g237(.A1(new_n659), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT84), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2096), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2100), .ZN(G227));
  XOR2_X1   g241(.A(G1971), .B(G1976), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1956), .B(G2474), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1961), .B(G1966), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AND2_X1   g246(.A1(new_n669), .A2(new_n670), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n668), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n668), .A2(new_n671), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT20), .Z(new_n675));
  AOI211_X1 g250(.A(new_n673), .B(new_n675), .C1(new_n668), .C2(new_n672), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1991), .B(G1996), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1981), .B(G1986), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n678), .B(new_n681), .ZN(G229));
  INV_X1    g257(.A(KEYINPUT36), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(KEYINPUT86), .ZN(new_n684));
  MUX2_X1   g259(.A(G95), .B(G107), .S(G2105), .Z(new_n685));
  AOI22_X1  g260(.A1(new_n481), .A2(G119), .B1(G2104), .B2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(G131), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n686), .B1(new_n687), .B2(new_n483), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n688), .A2(KEYINPUT85), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(KEYINPUT85), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  MUX2_X1   g266(.A(G25), .B(new_n691), .S(G29), .Z(new_n692));
  XOR2_X1   g267(.A(KEYINPUT35), .B(G1991), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(G16), .A2(G24), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(new_n598), .B2(G16), .ZN(new_n696));
  INV_X1    g271(.A(G1986), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  MUX2_X1   g273(.A(G6), .B(G305), .S(G16), .Z(new_n699));
  XOR2_X1   g274(.A(KEYINPUT32), .B(G1981), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G23), .ZN(new_n703));
  INV_X1    g278(.A(G288), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n703), .B1(new_n704), .B2(new_n702), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT33), .B(G1976), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(G16), .A2(G22), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G166), .B2(G16), .ZN(new_n709));
  INV_X1    g284(.A(G1971), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n701), .A2(new_n707), .A3(new_n711), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n694), .B(new_n698), .C1(new_n712), .C2(KEYINPUT34), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n712), .A2(KEYINPUT34), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n684), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n683), .A2(KEYINPUT86), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(G29), .A2(G33), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT87), .ZN(new_n719));
  AOI21_X1  g294(.A(KEYINPUT25), .B1(new_n468), .B2(G103), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n468), .A2(KEYINPUT25), .A3(G103), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n484), .A2(G139), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n479), .A2(G127), .ZN(new_n725));
  NAND2_X1  g300(.A1(G115), .A2(G2104), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n462), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G29), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n719), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G2072), .ZN(new_n732));
  INV_X1    g307(.A(G2084), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT24), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n730), .B1(new_n734), .B2(G34), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT88), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n735), .A2(new_n736), .B1(new_n734), .B2(G34), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n736), .B2(new_n735), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT89), .ZN(new_n739));
  INV_X1    g314(.A(G160), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n739), .B1(new_n730), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n730), .A2(G32), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n468), .A2(G105), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n484), .A2(G141), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n481), .A2(G129), .ZN(new_n745));
  NAND3_X1  g320(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT26), .Z(new_n747));
  AND4_X1   g322(.A1(new_n743), .A2(new_n744), .A3(new_n745), .A4(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n742), .B1(new_n748), .B2(new_n730), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT27), .B(G1996), .Z(new_n750));
  OAI221_X1 g325(.A(new_n732), .B1(new_n733), .B2(new_n741), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT90), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n730), .A2(G27), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G164), .B2(new_n730), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT94), .B(G2078), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(G299), .A2(G16), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n702), .A2(G20), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT23), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT96), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G1956), .ZN(new_n763));
  NOR2_X1   g338(.A1(G29), .A2(G35), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G162), .B2(G29), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT29), .Z(new_n766));
  INV_X1    g341(.A(G2090), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT95), .ZN(new_n769));
  NOR2_X1   g344(.A1(G16), .A2(G19), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n555), .B2(G16), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G1341), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(G171), .A2(new_n702), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G5), .B2(new_n702), .ZN(new_n775));
  INV_X1    g350(.A(G1961), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT31), .B(G11), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT92), .B(G28), .ZN(new_n779));
  AOI21_X1  g354(.A(G29), .B1(new_n779), .B2(KEYINPUT30), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n780), .A2(KEYINPUT93), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(KEYINPUT93), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(KEYINPUT30), .B2(new_n779), .ZN(new_n783));
  OAI221_X1 g358(.A(new_n778), .B1(new_n781), .B2(new_n783), .C1(new_n629), .C2(new_n730), .ZN(new_n784));
  NOR2_X1   g359(.A1(G168), .A2(new_n702), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n702), .B2(G21), .ZN(new_n786));
  INV_X1    g361(.A(G1966), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n784), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n749), .A2(new_n750), .B1(new_n741), .B2(new_n733), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n777), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n611), .A2(G16), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G4), .B2(G16), .ZN(new_n792));
  INV_X1    g367(.A(G1348), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n792), .A2(new_n793), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n730), .A2(G26), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT28), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n481), .A2(G128), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n484), .A2(G140), .ZN(new_n799));
  MUX2_X1   g374(.A(G104), .B(G116), .S(G2105), .Z(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(G2104), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n798), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n797), .B1(new_n803), .B2(new_n730), .ZN(new_n804));
  INV_X1    g379(.A(G2067), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n794), .A2(new_n795), .A3(new_n806), .ZN(new_n807));
  OAI22_X1  g382(.A1(new_n775), .A2(new_n776), .B1(new_n766), .B2(new_n767), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n786), .A2(new_n787), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT91), .Z(new_n810));
  NOR4_X1   g385(.A1(new_n790), .A2(new_n807), .A3(new_n808), .A4(new_n810), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n757), .A2(new_n763), .A3(new_n773), .A4(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n717), .A2(new_n812), .ZN(G311));
  INV_X1    g388(.A(G311), .ZN(G150));
  INV_X1    g389(.A(G93), .ZN(new_n815));
  INV_X1    g390(.A(G55), .ZN(new_n816));
  OAI22_X1  g391(.A1(new_n514), .A2(new_n815), .B1(new_n516), .B2(new_n816), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n818), .A2(new_n520), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n554), .B(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n606), .A2(new_n612), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n826), .A2(KEYINPUT39), .ZN(new_n827));
  INV_X1    g402(.A(G860), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(KEYINPUT39), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n820), .A2(new_n828), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT37), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n832), .ZN(G145));
  XNOR2_X1  g408(.A(new_n691), .B(new_n618), .ZN(new_n834));
  MUX2_X1   g409(.A(G106), .B(G118), .S(G2105), .Z(new_n835));
  AOI22_X1  g410(.A1(new_n481), .A2(G130), .B1(G2104), .B2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(G142), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n836), .B1(new_n837), .B2(new_n483), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n834), .B(new_n838), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n802), .B(new_n502), .Z(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n748), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(new_n728), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n629), .B(new_n488), .ZN(new_n846));
  XOR2_X1   g421(.A(G160), .B(KEYINPUT98), .Z(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n841), .A2(new_n844), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n845), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(KEYINPUT99), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT99), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n845), .A2(new_n852), .A3(new_n848), .A4(new_n849), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n848), .B1(new_n845), .B2(new_n849), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n855), .A2(G37), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g433(.A1(new_n821), .A2(G868), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n614), .B(KEYINPUT100), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n822), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n606), .B(G299), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n862), .A2(KEYINPUT41), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(KEYINPUT41), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT101), .ZN(new_n867));
  OAI22_X1  g442(.A1(new_n866), .A2(new_n867), .B1(new_n861), .B2(new_n862), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n868), .B1(new_n867), .B2(new_n866), .ZN(new_n869));
  XNOR2_X1  g444(.A(G305), .B(G303), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n598), .B(G288), .Z(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT102), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(new_n871), .B2(new_n870), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT42), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n874), .B(KEYINPUT103), .Z(new_n877));
  OAI21_X1  g452(.A(new_n876), .B1(new_n877), .B2(new_n875), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n869), .B(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n859), .B1(new_n879), .B2(G868), .ZN(G295));
  AOI21_X1  g455(.A(new_n859), .B1(new_n879), .B2(G868), .ZN(G331));
  INV_X1    g456(.A(KEYINPUT44), .ZN(new_n882));
  OR2_X1    g457(.A1(G168), .A2(KEYINPUT104), .ZN(new_n883));
  NAND2_X1  g458(.A1(G168), .A2(KEYINPUT104), .ZN(new_n884));
  NAND3_X1  g459(.A1(G301), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n885), .B1(G301), .B2(new_n884), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n886), .A2(new_n822), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n822), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n889), .A2(new_n862), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n888), .A2(KEYINPUT105), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(KEYINPUT105), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n891), .A2(new_n887), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n890), .B1(new_n865), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(G37), .B1(new_n877), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n893), .ZN(new_n897));
  INV_X1    g472(.A(new_n862), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT106), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n863), .A2(new_n899), .A3(new_n864), .ZN(new_n900));
  OAI211_X1 g475(.A(new_n889), .B(new_n900), .C1(new_n899), .C2(new_n864), .ZN(new_n901));
  AOI22_X1  g476(.A1(new_n897), .A2(new_n898), .B1(new_n901), .B2(KEYINPUT107), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n901), .A2(KEYINPUT107), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n877), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n896), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n905), .A2(KEYINPUT43), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n877), .A2(new_n894), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n895), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT43), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n882), .B1(new_n906), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n905), .A2(new_n909), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n908), .A2(KEYINPUT43), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT44), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n911), .A2(new_n914), .ZN(G397));
  INV_X1    g490(.A(KEYINPUT125), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT46), .ZN(new_n917));
  INV_X1    g492(.A(G1384), .ZN(new_n918));
  AOI21_X1  g493(.A(KEYINPUT45), .B1(new_n502), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(G40), .ZN(new_n920));
  NOR3_X1   g495(.A1(new_n471), .A2(new_n474), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n922), .A2(G1996), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n916), .A2(KEYINPUT46), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n917), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n922), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n802), .B(new_n805), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n927), .B1(new_n929), .B2(new_n842), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n926), .B(new_n930), .C1(new_n924), .C2(new_n917), .ZN(new_n931));
  XOR2_X1   g506(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n932));
  XNOR2_X1  g507(.A(new_n931), .B(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n691), .B(new_n693), .ZN(new_n934));
  OR2_X1    g509(.A1(new_n934), .A2(KEYINPUT110), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(KEYINPUT110), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n935), .A2(new_n927), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n923), .A2(new_n748), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(KEYINPUT109), .ZN(new_n939));
  INV_X1    g514(.A(G1996), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n928), .B1(new_n940), .B2(new_n748), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n939), .B1(new_n927), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n937), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n598), .A2(new_n697), .ZN(new_n944));
  XOR2_X1   g519(.A(new_n944), .B(KEYINPUT108), .Z(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n927), .ZN(new_n946));
  XOR2_X1   g521(.A(new_n946), .B(KEYINPUT48), .Z(new_n947));
  OAI21_X1  g522(.A(new_n933), .B1(new_n943), .B2(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n942), .A2(new_n690), .A3(new_n689), .A4(new_n693), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n803), .A2(new_n805), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n922), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(G1384), .B1(new_n507), .B2(new_n493), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n953), .A2(KEYINPUT50), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n508), .B1(new_n507), .B2(new_n493), .ZN(new_n956));
  AND4_X1   g531(.A1(new_n508), .A2(new_n493), .A3(new_n498), .A4(new_n501), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n918), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT50), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n955), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n960), .A2(new_n733), .A3(new_n921), .ZN(new_n961));
  INV_X1    g536(.A(new_n921), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT116), .B1(new_n919), .B2(new_n962), .ZN(new_n963));
  OAI211_X1 g538(.A(KEYINPUT45), .B(new_n918), .C1(new_n956), .C2(new_n957), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT116), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n965), .B(new_n921), .C1(new_n953), .C2(KEYINPUT45), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n963), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n967), .A2(KEYINPUT117), .A3(new_n787), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n961), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT117), .B1(new_n967), .B2(new_n787), .ZN(new_n970));
  OAI21_X1  g545(.A(G8), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G8), .ZN(new_n972));
  NOR2_X1   g547(.A1(G168), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT122), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT51), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n971), .A2(new_n974), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n967), .A2(new_n787), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT117), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n981), .A2(new_n968), .A3(new_n961), .ZN(new_n982));
  OAI211_X1 g557(.A(G8), .B(new_n976), .C1(new_n982), .C2(G286), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n982), .A2(G8), .A3(G286), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n978), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT62), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT112), .ZN(new_n987));
  OAI211_X1 g562(.A(G303), .B(G8), .C1(new_n987), .C2(KEYINPUT55), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(KEYINPUT55), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n988), .B(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT45), .B1(new_n510), .B2(new_n918), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT111), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n962), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(G1384), .B1(new_n503), .B2(new_n509), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n502), .A2(new_n918), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT45), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI22_X1  g572(.A1(new_n994), .A2(KEYINPUT45), .B1(new_n997), .B2(KEYINPUT111), .ZN(new_n998));
  AOI21_X1  g573(.A(G1971), .B1(new_n993), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n954), .B1(new_n994), .B2(KEYINPUT50), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n1000), .A2(G2090), .A3(new_n962), .ZN(new_n1001));
  OAI211_X1 g576(.A(G8), .B(new_n990), .C1(new_n999), .C2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n502), .A2(G160), .A3(G40), .A4(new_n918), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(G8), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT113), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1004), .A2(KEYINPUT113), .A3(G8), .ZN(new_n1008));
  AOI22_X1  g583(.A1(new_n1007), .A2(new_n1008), .B1(G1976), .B2(new_n704), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1003), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n704), .A2(G1976), .ZN(new_n1012));
  AOI211_X1 g587(.A(new_n1006), .B(new_n972), .C1(new_n953), .C2(new_n921), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT113), .B1(new_n1004), .B2(G8), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1012), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OR2_X1    g590(.A1(new_n704), .A2(G1976), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n1010), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1011), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT114), .B1(new_n1015), .B2(KEYINPUT52), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT49), .ZN(new_n1021));
  INV_X1    g596(.A(G1981), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n585), .B(new_n1022), .C1(new_n589), .C2(new_n591), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n1024));
  OAI21_X1  g599(.A(G1981), .B1(new_n1024), .B2(new_n588), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT115), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  AOI22_X1  g601(.A1(new_n1021), .A2(new_n1026), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1027));
  OR2_X1    g602(.A1(new_n1026), .A2(new_n1021), .ZN(new_n1028));
  AOI22_X1  g603(.A1(new_n1019), .A2(new_n1020), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1002), .A2(new_n1018), .A3(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n958), .A2(new_n992), .A3(new_n996), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n998), .A2(new_n921), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n710), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n995), .A2(new_n959), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1034), .B1(new_n958), .B2(new_n959), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1035), .A2(new_n962), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n767), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1033), .A2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n990), .B1(new_n1038), .B2(G8), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1030), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT62), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n978), .A2(new_n983), .A3(new_n1041), .A4(new_n984), .ZN(new_n1042));
  INV_X1    g617(.A(G2078), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n998), .A2(new_n1031), .A3(new_n1043), .A4(new_n921), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n960), .A2(new_n921), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n1044), .A2(new_n1045), .B1(new_n1046), .B2(new_n776), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1043), .A2(KEYINPUT53), .ZN(new_n1048));
  OR2_X1    g623(.A1(new_n967), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(G301), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n986), .A2(new_n1040), .A3(new_n1042), .A4(new_n1050), .ZN(new_n1051));
  AOI211_X1 g626(.A(G1976), .B(G288), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1023), .ZN(new_n1053));
  OAI22_X1  g628(.A1(new_n1052), .A2(new_n1053), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1009), .A2(new_n1003), .A3(new_n1010), .A4(new_n1016), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1054), .B1(new_n1060), .B2(new_n1002), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT63), .ZN(new_n1062));
  INV_X1    g637(.A(new_n990), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n710), .A2(new_n1032), .B1(new_n1036), .B2(new_n767), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1063), .B1(new_n1064), .B2(new_n972), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1059), .A2(new_n1065), .A3(new_n1002), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n982), .A2(G8), .A3(G168), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1062), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1067), .ZN(new_n1069));
  OAI21_X1  g644(.A(G8), .B1(new_n999), .B2(new_n1001), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1062), .B1(new_n1070), .B2(new_n1063), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1069), .A2(new_n1071), .A3(new_n1002), .A4(new_n1059), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1061), .B1(new_n1068), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1046), .A2(new_n776), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1074), .A2(new_n1075), .A3(new_n1049), .ZN(new_n1076));
  XNOR2_X1  g651(.A(G301), .B(KEYINPUT54), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NOR4_X1   g653(.A1(new_n997), .A2(new_n919), .A3(new_n962), .A4(new_n1048), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n1047), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1078), .A2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n985), .A2(new_n1040), .A3(KEYINPUT123), .A4(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n572), .A2(new_n563), .ZN(new_n1085));
  XOR2_X1   g660(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n1086));
  OAI22_X1  g661(.A1(G299), .A2(new_n1084), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  OR2_X1    g662(.A1(new_n1087), .A2(KEYINPUT119), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(KEYINPUT119), .ZN(new_n1089));
  XNOR2_X1  g664(.A(KEYINPUT56), .B(G2072), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n998), .A2(new_n1031), .A3(new_n921), .A4(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(G1956), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1092), .B1(new_n1035), .B2(new_n962), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1088), .A2(new_n1089), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1091), .A2(new_n1093), .A3(new_n1087), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n793), .B1(new_n1000), .B2(new_n962), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n953), .A2(new_n805), .A3(new_n921), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n606), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1094), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1096), .A2(new_n606), .A3(new_n1097), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(KEYINPUT60), .B1(new_n1101), .B2(new_n1098), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n606), .A2(KEYINPUT60), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1096), .A2(new_n1097), .A3(new_n1103), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1091), .A2(new_n1093), .A3(new_n1087), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1087), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1102), .B(new_n1104), .C1(new_n1107), .C2(KEYINPUT61), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n1109));
  XOR2_X1   g684(.A(KEYINPUT120), .B(G1996), .Z(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n993), .A2(new_n998), .A3(new_n1111), .ZN(new_n1112));
  XOR2_X1   g687(.A(KEYINPUT58), .B(G1341), .Z(new_n1113));
  NAND2_X1  g688(.A1(new_n1004), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1109), .B1(new_n1115), .B2(new_n555), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1109), .ZN(new_n1117));
  AOI211_X1 g692(.A(new_n554), .B(new_n1117), .C1(new_n1112), .C2(new_n1114), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1095), .A2(KEYINPUT61), .ZN(new_n1119));
  OAI22_X1  g694(.A1(new_n1116), .A2(new_n1118), .B1(new_n1094), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1099), .B1(new_n1108), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1083), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1078), .A2(new_n1081), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1066), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT123), .B1(new_n1124), .B2(new_n985), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1051), .B(new_n1073), .C1(new_n1122), .C2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n945), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(new_n697), .B2(new_n598), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n943), .B1(new_n927), .B2(new_n1128), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1126), .A2(KEYINPUT124), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(KEYINPUT124), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n952), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT127), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  OAI211_X1 g709(.A(KEYINPUT127), .B(new_n952), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g711(.A1(new_n906), .A2(new_n910), .ZN(new_n1138));
  NOR4_X1   g712(.A1(G229), .A2(G227), .A3(new_n460), .A4(G401), .ZN(new_n1139));
  AND3_X1   g713(.A1(new_n1138), .A2(new_n857), .A3(new_n1139), .ZN(G308));
  NAND3_X1  g714(.A1(new_n1138), .A2(new_n857), .A3(new_n1139), .ZN(G225));
endmodule


