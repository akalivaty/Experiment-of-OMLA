

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584;

  XNOR2_X1 U323 ( .A(KEYINPUT54), .B(KEYINPUT117), .ZN(n540) );
  XNOR2_X1 U324 ( .A(n360), .B(KEYINPUT95), .ZN(n361) );
  XOR2_X1 U325 ( .A(n395), .B(n394), .Z(n542) );
  XNOR2_X1 U326 ( .A(n344), .B(KEYINPUT24), .ZN(n345) );
  XNOR2_X1 U327 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U328 ( .A(n391), .B(n345), .ZN(n346) );
  XNOR2_X1 U329 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U330 ( .A(n541), .B(n540), .ZN(n543) );
  XNOR2_X1 U331 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U332 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U333 ( .A(n362), .B(n361), .ZN(n563) );
  XNOR2_X1 U334 ( .A(n354), .B(n353), .ZN(n359) );
  XNOR2_X1 U335 ( .A(n444), .B(n443), .ZN(n445) );
  NOR2_X1 U336 ( .A1(n548), .A2(n547), .ZN(n559) );
  INV_X1 U337 ( .A(G43GAT), .ZN(n448) );
  XNOR2_X1 U338 ( .A(n448), .B(KEYINPUT40), .ZN(n449) );
  XNOR2_X1 U339 ( .A(n450), .B(n449), .ZN(G1330GAT) );
  XOR2_X1 U340 ( .A(G78GAT), .B(G71GAT), .Z(n292) );
  XNOR2_X1 U341 ( .A(G22GAT), .B(G183GAT), .ZN(n291) );
  XNOR2_X1 U342 ( .A(n292), .B(n291), .ZN(n296) );
  XOR2_X1 U343 ( .A(KEYINPUT14), .B(KEYINPUT80), .Z(n294) );
  XNOR2_X1 U344 ( .A(G64GAT), .B(KEYINPUT81), .ZN(n293) );
  XNOR2_X1 U345 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U346 ( .A(n296), .B(n295), .Z(n301) );
  XOR2_X1 U347 ( .A(G15GAT), .B(G127GAT), .Z(n334) );
  XOR2_X1 U348 ( .A(KEYINPUT84), .B(KEYINPUT12), .Z(n298) );
  NAND2_X1 U349 ( .A1(G231GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U350 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U351 ( .A(n334), .B(n299), .ZN(n300) );
  XNOR2_X1 U352 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U353 ( .A(G8GAT), .B(KEYINPUT78), .Z(n368) );
  XOR2_X1 U354 ( .A(KEYINPUT13), .B(G57GAT), .Z(n442) );
  XOR2_X1 U355 ( .A(n368), .B(n442), .Z(n303) );
  XNOR2_X1 U356 ( .A(G211GAT), .B(G155GAT), .ZN(n302) );
  XNOR2_X1 U357 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U358 ( .A(n305), .B(n304), .Z(n310) );
  XOR2_X1 U359 ( .A(KEYINPUT72), .B(G1GAT), .Z(n422) );
  XOR2_X1 U360 ( .A(KEYINPUT15), .B(KEYINPUT83), .Z(n307) );
  XNOR2_X1 U361 ( .A(KEYINPUT82), .B(KEYINPUT79), .ZN(n306) );
  XNOR2_X1 U362 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U363 ( .A(n422), .B(n308), .ZN(n309) );
  XNOR2_X1 U364 ( .A(n310), .B(n309), .ZN(n578) );
  XOR2_X1 U365 ( .A(G36GAT), .B(G190GAT), .Z(n364) );
  XOR2_X1 U366 ( .A(KEYINPUT9), .B(KEYINPUT66), .Z(n312) );
  XNOR2_X1 U367 ( .A(G92GAT), .B(KEYINPUT11), .ZN(n311) );
  XNOR2_X1 U368 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U369 ( .A(n364), .B(n313), .Z(n317) );
  XOR2_X1 U370 ( .A(G29GAT), .B(G43GAT), .Z(n315) );
  XNOR2_X1 U371 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n314) );
  XNOR2_X1 U372 ( .A(n315), .B(n314), .ZN(n425) );
  XOR2_X1 U373 ( .A(G50GAT), .B(G162GAT), .Z(n348) );
  XNOR2_X1 U374 ( .A(n425), .B(n348), .ZN(n316) );
  XNOR2_X1 U375 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U376 ( .A(n318), .B(KEYINPUT77), .Z(n320) );
  XOR2_X1 U377 ( .A(G99GAT), .B(G85GAT), .Z(n432) );
  XNOR2_X1 U378 ( .A(G218GAT), .B(n432), .ZN(n319) );
  XNOR2_X1 U379 ( .A(n320), .B(n319), .ZN(n325) );
  XOR2_X1 U380 ( .A(G106GAT), .B(KEYINPUT10), .Z(n322) );
  NAND2_X1 U381 ( .A1(G232GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U382 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U383 ( .A(G134GAT), .B(n323), .Z(n324) );
  XNOR2_X1 U384 ( .A(n325), .B(n324), .ZN(n558) );
  INV_X1 U385 ( .A(n558), .ZN(n536) );
  XNOR2_X1 U386 ( .A(n536), .B(KEYINPUT36), .ZN(n580) );
  XNOR2_X1 U387 ( .A(KEYINPUT19), .B(KEYINPUT85), .ZN(n326) );
  XNOR2_X1 U388 ( .A(n326), .B(KEYINPUT18), .ZN(n327) );
  XOR2_X1 U389 ( .A(n327), .B(KEYINPUT17), .Z(n329) );
  XNOR2_X1 U390 ( .A(G169GAT), .B(G183GAT), .ZN(n328) );
  XNOR2_X1 U391 ( .A(n329), .B(n328), .ZN(n372) );
  XOR2_X1 U392 ( .A(KEYINPUT20), .B(KEYINPUT65), .Z(n331) );
  XNOR2_X1 U393 ( .A(G99GAT), .B(G176GAT), .ZN(n330) );
  XNOR2_X1 U394 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U395 ( .A(n372), .B(n332), .ZN(n341) );
  XNOR2_X1 U396 ( .A(G113GAT), .B(G134GAT), .ZN(n333) );
  XNOR2_X1 U397 ( .A(n333), .B(KEYINPUT0), .ZN(n384) );
  XOR2_X1 U398 ( .A(n334), .B(n384), .Z(n336) );
  NAND2_X1 U399 ( .A1(G227GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U400 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U401 ( .A(G120GAT), .B(G71GAT), .Z(n436) );
  XOR2_X1 U402 ( .A(n337), .B(n436), .Z(n339) );
  XNOR2_X1 U403 ( .A(G43GAT), .B(G190GAT), .ZN(n338) );
  XNOR2_X1 U404 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X2 U405 ( .A(n341), .B(n340), .ZN(n548) );
  XOR2_X1 U406 ( .A(G141GAT), .B(G22GAT), .Z(n424) );
  XOR2_X1 U407 ( .A(G155GAT), .B(KEYINPUT2), .Z(n343) );
  XNOR2_X1 U408 ( .A(KEYINPUT3), .B(KEYINPUT88), .ZN(n342) );
  XNOR2_X1 U409 ( .A(n343), .B(n342), .ZN(n391) );
  AND2_X1 U410 ( .A1(G228GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U411 ( .A(n424), .B(n346), .ZN(n354) );
  XNOR2_X1 U412 ( .A(G106GAT), .B(G78GAT), .ZN(n347) );
  XNOR2_X1 U413 ( .A(n347), .B(G148GAT), .ZN(n434) );
  XOR2_X1 U414 ( .A(n434), .B(n348), .Z(n352) );
  XOR2_X1 U415 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n350) );
  XNOR2_X1 U416 ( .A(KEYINPUT89), .B(KEYINPUT86), .ZN(n349) );
  XNOR2_X1 U417 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U418 ( .A(KEYINPUT87), .B(G204GAT), .Z(n356) );
  XNOR2_X1 U419 ( .A(G197GAT), .B(G211GAT), .ZN(n355) );
  XNOR2_X1 U420 ( .A(n356), .B(n355), .ZN(n358) );
  XOR2_X1 U421 ( .A(G218GAT), .B(KEYINPUT21), .Z(n357) );
  XNOR2_X1 U422 ( .A(n358), .B(n357), .ZN(n373) );
  XNOR2_X1 U423 ( .A(n359), .B(n373), .ZN(n544) );
  AND2_X1 U424 ( .A1(n548), .A2(n544), .ZN(n362) );
  XNOR2_X1 U425 ( .A(KEYINPUT96), .B(KEYINPUT26), .ZN(n360) );
  XNOR2_X1 U426 ( .A(G176GAT), .B(G92GAT), .ZN(n363) );
  XNOR2_X1 U427 ( .A(n363), .B(G64GAT), .ZN(n433) );
  XOR2_X1 U428 ( .A(n364), .B(n433), .Z(n366) );
  NAND2_X1 U429 ( .A1(G226GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U430 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U431 ( .A(n367), .B(KEYINPUT93), .Z(n370) );
  XNOR2_X1 U432 ( .A(n368), .B(KEYINPUT94), .ZN(n369) );
  XNOR2_X1 U433 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U434 ( .A(n372), .B(n371), .ZN(n374) );
  XNOR2_X1 U435 ( .A(n374), .B(n373), .ZN(n538) );
  XOR2_X1 U436 ( .A(KEYINPUT27), .B(n538), .Z(n510) );
  NOR2_X1 U437 ( .A1(n563), .A2(n510), .ZN(n375) );
  XNOR2_X1 U438 ( .A(n375), .B(KEYINPUT97), .ZN(n396) );
  XOR2_X1 U439 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n377) );
  XNOR2_X1 U440 ( .A(KEYINPUT5), .B(KEYINPUT91), .ZN(n376) );
  XNOR2_X1 U441 ( .A(n377), .B(n376), .ZN(n395) );
  XOR2_X1 U442 ( .A(G85GAT), .B(G148GAT), .Z(n379) );
  XNOR2_X1 U443 ( .A(G141GAT), .B(G127GAT), .ZN(n378) );
  XNOR2_X1 U444 ( .A(n379), .B(n378), .ZN(n383) );
  XOR2_X1 U445 ( .A(KEYINPUT92), .B(G57GAT), .Z(n381) );
  XNOR2_X1 U446 ( .A(G1GAT), .B(G120GAT), .ZN(n380) );
  XNOR2_X1 U447 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U448 ( .A(n383), .B(n382), .Z(n389) );
  XOR2_X1 U449 ( .A(G162GAT), .B(n384), .Z(n386) );
  NAND2_X1 U450 ( .A1(G225GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U451 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U452 ( .A(G29GAT), .B(n387), .ZN(n388) );
  XNOR2_X1 U453 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U454 ( .A(n390), .B(KEYINPUT90), .Z(n393) );
  XNOR2_X1 U455 ( .A(n391), .B(KEYINPUT6), .ZN(n392) );
  XNOR2_X1 U456 ( .A(n393), .B(n392), .ZN(n394) );
  NAND2_X1 U457 ( .A1(n396), .A2(n542), .ZN(n400) );
  INV_X1 U458 ( .A(n538), .ZN(n489) );
  NOR2_X1 U459 ( .A1(n548), .A2(n489), .ZN(n397) );
  NOR2_X1 U460 ( .A1(n544), .A2(n397), .ZN(n398) );
  XOR2_X1 U461 ( .A(KEYINPUT25), .B(n398), .Z(n399) );
  NOR2_X1 U462 ( .A1(n400), .A2(n399), .ZN(n404) );
  XOR2_X1 U463 ( .A(KEYINPUT28), .B(n544), .Z(n513) );
  NAND2_X1 U464 ( .A1(n548), .A2(n513), .ZN(n401) );
  NOR2_X1 U465 ( .A1(n401), .A2(n510), .ZN(n402) );
  NOR2_X1 U466 ( .A1(n542), .A2(n402), .ZN(n403) );
  NOR2_X1 U467 ( .A1(n404), .A2(n403), .ZN(n405) );
  XOR2_X1 U468 ( .A(KEYINPUT98), .B(n405), .Z(n453) );
  NOR2_X1 U469 ( .A1(n580), .A2(n453), .ZN(n406) );
  NAND2_X1 U470 ( .A1(n578), .A2(n406), .ZN(n407) );
  XNOR2_X1 U471 ( .A(KEYINPUT104), .B(n407), .ZN(n408) );
  XNOR2_X1 U472 ( .A(n408), .B(KEYINPUT37), .ZN(n485) );
  XOR2_X1 U473 ( .A(KEYINPUT71), .B(KEYINPUT68), .Z(n410) );
  XNOR2_X1 U474 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n409) );
  XNOR2_X1 U475 ( .A(n410), .B(n409), .ZN(n429) );
  XOR2_X1 U476 ( .A(G113GAT), .B(G197GAT), .Z(n412) );
  XNOR2_X1 U477 ( .A(G36GAT), .B(G50GAT), .ZN(n411) );
  XNOR2_X1 U478 ( .A(n412), .B(n411), .ZN(n416) );
  XOR2_X1 U479 ( .A(KEYINPUT73), .B(KEYINPUT70), .Z(n414) );
  XNOR2_X1 U480 ( .A(G169GAT), .B(G15GAT), .ZN(n413) );
  XNOR2_X1 U481 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U482 ( .A(n416), .B(n415), .Z(n421) );
  XOR2_X1 U483 ( .A(KEYINPUT67), .B(G8GAT), .Z(n418) );
  NAND2_X1 U484 ( .A1(G229GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U485 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U486 ( .A(KEYINPUT69), .B(n419), .ZN(n420) );
  XNOR2_X1 U487 ( .A(n421), .B(n420), .ZN(n423) );
  XOR2_X1 U488 ( .A(n423), .B(n422), .Z(n427) );
  XNOR2_X1 U489 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U490 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U491 ( .A(n429), .B(n428), .ZN(n549) );
  INV_X1 U492 ( .A(n549), .ZN(n567) );
  XOR2_X1 U493 ( .A(KEYINPUT76), .B(KEYINPUT74), .Z(n431) );
  XNOR2_X1 U494 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n430) );
  XNOR2_X1 U495 ( .A(n431), .B(n430), .ZN(n446) );
  XOR2_X1 U496 ( .A(n433), .B(n432), .Z(n440) );
  XOR2_X1 U497 ( .A(n434), .B(KEYINPUT75), .Z(n438) );
  NAND2_X1 U498 ( .A1(G230GAT), .A2(G233GAT), .ZN(n435) );
  XOR2_X1 U499 ( .A(n440), .B(n439), .Z(n444) );
  XNOR2_X1 U500 ( .A(G204GAT), .B(KEYINPUT33), .ZN(n441) );
  XOR2_X1 U501 ( .A(n446), .B(n445), .Z(n575) );
  INV_X1 U502 ( .A(n575), .ZN(n504) );
  NOR2_X1 U503 ( .A1(n567), .A2(n504), .ZN(n454) );
  NAND2_X1 U504 ( .A1(n485), .A2(n454), .ZN(n447) );
  XNOR2_X1 U505 ( .A(n447), .B(KEYINPUT38), .ZN(n473) );
  NOR2_X1 U506 ( .A1(n473), .A2(n548), .ZN(n450) );
  NOR2_X1 U507 ( .A1(n578), .A2(n558), .ZN(n451) );
  XOR2_X1 U508 ( .A(KEYINPUT16), .B(n451), .Z(n452) );
  NOR2_X1 U509 ( .A1(n453), .A2(n452), .ZN(n476) );
  NAND2_X1 U510 ( .A1(n454), .A2(n476), .ZN(n462) );
  NOR2_X1 U511 ( .A1(n542), .A2(n462), .ZN(n456) );
  XNOR2_X1 U512 ( .A(KEYINPUT34), .B(KEYINPUT99), .ZN(n455) );
  XNOR2_X1 U513 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U514 ( .A(G1GAT), .B(n457), .ZN(G1324GAT) );
  NOR2_X1 U515 ( .A1(n489), .A2(n462), .ZN(n458) );
  XOR2_X1 U516 ( .A(G8GAT), .B(n458), .Z(G1325GAT) );
  NOR2_X1 U517 ( .A1(n548), .A2(n462), .ZN(n460) );
  XNOR2_X1 U518 ( .A(KEYINPUT100), .B(KEYINPUT35), .ZN(n459) );
  XNOR2_X1 U519 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U520 ( .A(G15GAT), .B(n461), .ZN(G1326GAT) );
  NOR2_X1 U521 ( .A1(n513), .A2(n462), .ZN(n464) );
  XNOR2_X1 U522 ( .A(KEYINPUT101), .B(KEYINPUT102), .ZN(n463) );
  XNOR2_X1 U523 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U524 ( .A(G22GAT), .B(n465), .ZN(G1327GAT) );
  XOR2_X1 U525 ( .A(KEYINPUT105), .B(KEYINPUT39), .Z(n467) );
  XNOR2_X1 U526 ( .A(G29GAT), .B(KEYINPUT103), .ZN(n466) );
  XNOR2_X1 U527 ( .A(n467), .B(n466), .ZN(n469) );
  NOR2_X1 U528 ( .A1(n542), .A2(n473), .ZN(n468) );
  XOR2_X1 U529 ( .A(n469), .B(n468), .Z(G1328GAT) );
  INV_X1 U530 ( .A(KEYINPUT106), .ZN(n471) );
  NOR2_X1 U531 ( .A1(n489), .A2(n473), .ZN(n470) );
  XNOR2_X1 U532 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U533 ( .A(G36GAT), .B(n472), .ZN(G1329GAT) );
  NOR2_X1 U534 ( .A1(n473), .A2(n513), .ZN(n474) );
  XOR2_X1 U535 ( .A(G50GAT), .B(n474), .Z(G1331GAT) );
  XNOR2_X1 U536 ( .A(n575), .B(KEYINPUT41), .ZN(n497) );
  INV_X1 U537 ( .A(n497), .ZN(n528) );
  NAND2_X1 U538 ( .A1(n497), .A2(n567), .ZN(n475) );
  XNOR2_X1 U539 ( .A(n475), .B(KEYINPUT107), .ZN(n486) );
  NAND2_X1 U540 ( .A1(n476), .A2(n486), .ZN(n477) );
  XNOR2_X1 U541 ( .A(n477), .B(KEYINPUT108), .ZN(n482) );
  NOR2_X1 U542 ( .A1(n542), .A2(n482), .ZN(n478) );
  XOR2_X1 U543 ( .A(KEYINPUT42), .B(n478), .Z(n479) );
  XNOR2_X1 U544 ( .A(G57GAT), .B(n479), .ZN(G1332GAT) );
  NOR2_X1 U545 ( .A1(n489), .A2(n482), .ZN(n480) );
  XOR2_X1 U546 ( .A(G64GAT), .B(n480), .Z(G1333GAT) );
  NOR2_X1 U547 ( .A1(n548), .A2(n482), .ZN(n481) );
  XOR2_X1 U548 ( .A(G71GAT), .B(n481), .Z(G1334GAT) );
  NOR2_X1 U549 ( .A1(n482), .A2(n513), .ZN(n484) );
  XNOR2_X1 U550 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n483) );
  XNOR2_X1 U551 ( .A(n484), .B(n483), .ZN(G1335GAT) );
  NAND2_X1 U552 ( .A1(n486), .A2(n485), .ZN(n493) );
  NOR2_X1 U553 ( .A1(n542), .A2(n493), .ZN(n488) );
  XNOR2_X1 U554 ( .A(G85GAT), .B(KEYINPUT109), .ZN(n487) );
  XNOR2_X1 U555 ( .A(n488), .B(n487), .ZN(G1336GAT) );
  NOR2_X1 U556 ( .A1(n489), .A2(n493), .ZN(n490) );
  XOR2_X1 U557 ( .A(KEYINPUT110), .B(n490), .Z(n491) );
  XNOR2_X1 U558 ( .A(G92GAT), .B(n491), .ZN(G1337GAT) );
  NOR2_X1 U559 ( .A1(n548), .A2(n493), .ZN(n492) );
  XOR2_X1 U560 ( .A(G99GAT), .B(n492), .Z(G1338GAT) );
  NOR2_X1 U561 ( .A1(n513), .A2(n493), .ZN(n495) );
  XNOR2_X1 U562 ( .A(KEYINPUT44), .B(KEYINPUT111), .ZN(n494) );
  XNOR2_X1 U563 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U564 ( .A(G106GAT), .B(n496), .ZN(G1339GAT) );
  AND2_X1 U565 ( .A1(n549), .A2(n497), .ZN(n498) );
  XNOR2_X1 U566 ( .A(n498), .B(KEYINPUT46), .ZN(n500) );
  NAND2_X1 U567 ( .A1(n578), .A2(n536), .ZN(n499) );
  NOR2_X1 U568 ( .A1(n500), .A2(n499), .ZN(n501) );
  XNOR2_X1 U569 ( .A(n501), .B(KEYINPUT47), .ZN(n507) );
  NOR2_X1 U570 ( .A1(n578), .A2(n580), .ZN(n502) );
  XOR2_X1 U571 ( .A(KEYINPUT45), .B(n502), .Z(n503) );
  NOR2_X1 U572 ( .A1(n504), .A2(n503), .ZN(n505) );
  NAND2_X1 U573 ( .A1(n505), .A2(n567), .ZN(n506) );
  NAND2_X1 U574 ( .A1(n507), .A2(n506), .ZN(n509) );
  XNOR2_X1 U575 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n509), .B(n508), .ZN(n539) );
  NOR2_X1 U577 ( .A1(n542), .A2(n510), .ZN(n511) );
  NAND2_X1 U578 ( .A1(n539), .A2(n511), .ZN(n512) );
  XOR2_X1 U579 ( .A(KEYINPUT112), .B(n512), .Z(n525) );
  NAND2_X1 U580 ( .A1(n513), .A2(n525), .ZN(n514) );
  NOR2_X1 U581 ( .A1(n548), .A2(n514), .ZN(n522) );
  NAND2_X1 U582 ( .A1(n549), .A2(n522), .ZN(n515) );
  XNOR2_X1 U583 ( .A(n515), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT113), .B(KEYINPUT49), .Z(n517) );
  NAND2_X1 U585 ( .A1(n522), .A2(n497), .ZN(n516) );
  XNOR2_X1 U586 ( .A(n517), .B(n516), .ZN(n518) );
  XOR2_X1 U587 ( .A(G120GAT), .B(n518), .Z(G1341GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n520) );
  INV_X1 U589 ( .A(n578), .ZN(n556) );
  NAND2_X1 U590 ( .A1(n522), .A2(n556), .ZN(n519) );
  XNOR2_X1 U591 ( .A(n520), .B(n519), .ZN(n521) );
  XOR2_X1 U592 ( .A(G127GAT), .B(n521), .Z(G1342GAT) );
  XOR2_X1 U593 ( .A(G134GAT), .B(KEYINPUT51), .Z(n524) );
  NAND2_X1 U594 ( .A1(n522), .A2(n558), .ZN(n523) );
  XNOR2_X1 U595 ( .A(n524), .B(n523), .ZN(G1343GAT) );
  INV_X1 U596 ( .A(n563), .ZN(n526) );
  NAND2_X1 U597 ( .A1(n526), .A2(n525), .ZN(n535) );
  NOR2_X1 U598 ( .A1(n567), .A2(n535), .ZN(n527) );
  XOR2_X1 U599 ( .A(G141GAT), .B(n527), .Z(G1344GAT) );
  NOR2_X1 U600 ( .A1(n535), .A2(n528), .ZN(n532) );
  XOR2_X1 U601 ( .A(KEYINPUT115), .B(KEYINPUT52), .Z(n530) );
  XNOR2_X1 U602 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n529) );
  XNOR2_X1 U603 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U604 ( .A(n532), .B(n531), .ZN(G1345GAT) );
  NOR2_X1 U605 ( .A1(n578), .A2(n535), .ZN(n533) );
  XOR2_X1 U606 ( .A(KEYINPUT116), .B(n533), .Z(n534) );
  XNOR2_X1 U607 ( .A(G155GAT), .B(n534), .ZN(G1346GAT) );
  NOR2_X1 U608 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U609 ( .A(G162GAT), .B(n537), .Z(G1347GAT) );
  NAND2_X1 U610 ( .A1(n539), .A2(n538), .ZN(n541) );
  NAND2_X1 U611 ( .A1(n543), .A2(n542), .ZN(n564) );
  NOR2_X1 U612 ( .A1(n544), .A2(n564), .ZN(n546) );
  XNOR2_X1 U613 ( .A(KEYINPUT55), .B(KEYINPUT118), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(n547) );
  NAND2_X1 U615 ( .A1(n559), .A2(n549), .ZN(n550) );
  XNOR2_X1 U616 ( .A(G169GAT), .B(n550), .ZN(G1348GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT57), .B(KEYINPUT120), .Z(n552) );
  XNOR2_X1 U618 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U620 ( .A(KEYINPUT119), .B(n553), .Z(n555) );
  NAND2_X1 U621 ( .A1(n559), .A2(n497), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(G1349GAT) );
  NAND2_X1 U623 ( .A1(n556), .A2(n559), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n557), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT58), .B(KEYINPUT121), .Z(n561) );
  NAND2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(G190GAT), .B(n562), .ZN(G1351GAT) );
  INV_X1 U629 ( .A(KEYINPUT122), .ZN(n566) );
  NOR2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(n581) );
  NOR2_X1 U632 ( .A1(n581), .A2(n567), .ZN(n571) );
  XOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n569) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n573) );
  XNOR2_X1 U638 ( .A(G204GAT), .B(KEYINPUT125), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(KEYINPUT124), .B(n574), .ZN(n577) );
  NOR2_X1 U641 ( .A1(n575), .A2(n581), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NOR2_X1 U643 ( .A1(n578), .A2(n581), .ZN(n579) );
  XOR2_X1 U644 ( .A(G211GAT), .B(n579), .Z(G1354GAT) );
  NOR2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n583) );
  XNOR2_X1 U646 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

