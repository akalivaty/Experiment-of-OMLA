

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585;

  XNOR2_X1 U323 ( .A(n456), .B(n455), .ZN(n460) );
  XNOR2_X1 U324 ( .A(n398), .B(n352), .ZN(n358) );
  XNOR2_X1 U325 ( .A(n447), .B(n446), .ZN(n524) );
  XNOR2_X1 U326 ( .A(n347), .B(n432), .ZN(n513) );
  XNOR2_X1 U327 ( .A(KEYINPUT95), .B(KEYINPUT25), .ZN(n455) );
  XNOR2_X1 U328 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n384) );
  XNOR2_X1 U329 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U330 ( .A(n385), .B(n384), .ZN(n406) );
  XOR2_X1 U331 ( .A(G176GAT), .B(G64GAT), .Z(n351) );
  INV_X1 U332 ( .A(KEYINPUT93), .ZN(n336) );
  NOR2_X1 U333 ( .A1(n412), .A2(n411), .ZN(n413) );
  XNOR2_X1 U334 ( .A(n337), .B(n336), .ZN(n338) );
  NOR2_X1 U335 ( .A1(n509), .A2(n416), .ZN(n567) );
  XNOR2_X1 U336 ( .A(n339), .B(n338), .ZN(n342) );
  XOR2_X1 U337 ( .A(n369), .B(n428), .Z(n573) );
  XOR2_X1 U338 ( .A(KEYINPUT28), .B(n464), .Z(n527) );
  XNOR2_X1 U339 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U340 ( .A(n452), .B(n451), .ZN(G1351GAT) );
  XOR2_X1 U341 ( .A(KEYINPUT72), .B(G92GAT), .Z(n292) );
  XNOR2_X1 U342 ( .A(G99GAT), .B(G85GAT), .ZN(n291) );
  XNOR2_X1 U343 ( .A(n292), .B(n291), .ZN(n366) );
  XOR2_X1 U344 ( .A(G190GAT), .B(KEYINPUT76), .Z(n329) );
  XOR2_X1 U345 ( .A(n366), .B(n329), .Z(n294) );
  NAND2_X1 U346 ( .A1(G232GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U347 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U348 ( .A(KEYINPUT10), .B(G162GAT), .Z(n296) );
  XNOR2_X1 U349 ( .A(G134GAT), .B(G106GAT), .ZN(n295) );
  XNOR2_X1 U350 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U351 ( .A(n298), .B(n297), .Z(n308) );
  XOR2_X1 U352 ( .A(G29GAT), .B(KEYINPUT8), .Z(n300) );
  XNOR2_X1 U353 ( .A(G43GAT), .B(G36GAT), .ZN(n299) );
  XNOR2_X1 U354 ( .A(n300), .B(n299), .ZN(n302) );
  XOR2_X1 U355 ( .A(G50GAT), .B(KEYINPUT7), .Z(n301) );
  XNOR2_X1 U356 ( .A(n302), .B(n301), .ZN(n382) );
  INV_X1 U357 ( .A(n382), .ZN(n306) );
  XOR2_X1 U358 ( .A(KEYINPUT75), .B(KEYINPUT9), .Z(n304) );
  XNOR2_X1 U359 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n303) );
  XNOR2_X1 U360 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U361 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U362 ( .A(n308), .B(n307), .ZN(n535) );
  INV_X1 U363 ( .A(n535), .ZN(n548) );
  XOR2_X1 U364 ( .A(KEYINPUT91), .B(KEYINPUT5), .Z(n310) );
  XNOR2_X1 U365 ( .A(KEYINPUT89), .B(KEYINPUT90), .ZN(n309) );
  XNOR2_X1 U366 ( .A(n310), .B(n309), .ZN(n328) );
  XOR2_X1 U367 ( .A(G85GAT), .B(G148GAT), .Z(n312) );
  XNOR2_X1 U368 ( .A(G29GAT), .B(G141GAT), .ZN(n311) );
  XNOR2_X1 U369 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U370 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n314) );
  XNOR2_X1 U371 ( .A(G1GAT), .B(G57GAT), .ZN(n313) );
  XNOR2_X1 U372 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U373 ( .A(n316), .B(n315), .Z(n326) );
  XOR2_X1 U374 ( .A(G127GAT), .B(G134GAT), .Z(n318) );
  XNOR2_X1 U375 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n317) );
  XNOR2_X1 U376 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U377 ( .A(G113GAT), .B(n319), .Z(n439) );
  XOR2_X1 U378 ( .A(G155GAT), .B(KEYINPUT3), .Z(n321) );
  XNOR2_X1 U379 ( .A(G162GAT), .B(KEYINPUT2), .ZN(n320) );
  XNOR2_X1 U380 ( .A(n321), .B(n320), .ZN(n427) );
  XOR2_X1 U381 ( .A(n427), .B(KEYINPUT1), .Z(n323) );
  NAND2_X1 U382 ( .A1(G225GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U383 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U384 ( .A(n439), .B(n324), .ZN(n325) );
  XNOR2_X1 U385 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U386 ( .A(n328), .B(n327), .ZN(n509) );
  XOR2_X1 U387 ( .A(n329), .B(n351), .Z(n331) );
  NAND2_X1 U388 ( .A1(G226GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U389 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U390 ( .A(n332), .B(G92GAT), .Z(n339) );
  XOR2_X1 U391 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n334) );
  XNOR2_X1 U392 ( .A(KEYINPUT18), .B(KEYINPUT82), .ZN(n333) );
  XNOR2_X1 U393 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U394 ( .A(G169GAT), .B(n335), .Z(n438) );
  XNOR2_X1 U395 ( .A(G36GAT), .B(n438), .ZN(n337) );
  XNOR2_X1 U396 ( .A(G8GAT), .B(G183GAT), .ZN(n340) );
  XNOR2_X1 U397 ( .A(n340), .B(G211GAT), .ZN(n399) );
  XNOR2_X1 U398 ( .A(KEYINPUT92), .B(n399), .ZN(n341) );
  XNOR2_X1 U399 ( .A(n342), .B(n341), .ZN(n347) );
  XOR2_X1 U400 ( .A(KEYINPUT84), .B(KEYINPUT21), .Z(n344) );
  XNOR2_X1 U401 ( .A(G197GAT), .B(G204GAT), .ZN(n343) );
  XNOR2_X1 U402 ( .A(n344), .B(n343), .ZN(n346) );
  XOR2_X1 U403 ( .A(G218GAT), .B(KEYINPUT85), .Z(n345) );
  XOR2_X1 U404 ( .A(n346), .B(n345), .Z(n432) );
  INV_X1 U405 ( .A(n513), .ZN(n414) );
  XNOR2_X1 U406 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n370) );
  XOR2_X1 U407 ( .A(KEYINPUT69), .B(KEYINPUT13), .Z(n349) );
  XNOR2_X1 U408 ( .A(G71GAT), .B(G57GAT), .ZN(n348) );
  XNOR2_X1 U409 ( .A(n349), .B(n348), .ZN(n398) );
  XOR2_X1 U410 ( .A(G120GAT), .B(G204GAT), .Z(n350) );
  INV_X1 U411 ( .A(n358), .ZN(n356) );
  XOR2_X1 U412 ( .A(KEYINPUT73), .B(KEYINPUT31), .Z(n354) );
  NAND2_X1 U413 ( .A1(G230GAT), .A2(G233GAT), .ZN(n353) );
  XOR2_X1 U414 ( .A(n354), .B(n353), .Z(n357) );
  INV_X1 U415 ( .A(n357), .ZN(n355) );
  NAND2_X1 U416 ( .A1(n356), .A2(n355), .ZN(n360) );
  NAND2_X1 U417 ( .A1(n358), .A2(n357), .ZN(n359) );
  NAND2_X1 U418 ( .A1(n360), .A2(n359), .ZN(n365) );
  XOR2_X1 U419 ( .A(KEYINPUT33), .B(KEYINPUT74), .Z(n362) );
  XNOR2_X1 U420 ( .A(KEYINPUT32), .B(KEYINPUT70), .ZN(n361) );
  XNOR2_X1 U421 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U422 ( .A(n363), .B(KEYINPUT71), .ZN(n364) );
  XNOR2_X1 U423 ( .A(n365), .B(n364), .ZN(n367) );
  XNOR2_X1 U424 ( .A(n367), .B(n366), .ZN(n369) );
  XOR2_X1 U425 ( .A(G106GAT), .B(G78GAT), .Z(n368) );
  XOR2_X1 U426 ( .A(G148GAT), .B(n368), .Z(n428) );
  XNOR2_X1 U427 ( .A(n370), .B(n573), .ZN(n529) );
  XOR2_X1 U428 ( .A(G15GAT), .B(G1GAT), .Z(n389) );
  XOR2_X1 U429 ( .A(n389), .B(KEYINPUT30), .Z(n372) );
  NAND2_X1 U430 ( .A1(G229GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U431 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U432 ( .A(G141GAT), .B(G22GAT), .Z(n420) );
  XOR2_X1 U433 ( .A(n373), .B(n420), .Z(n381) );
  XOR2_X1 U434 ( .A(G8GAT), .B(G197GAT), .Z(n375) );
  XNOR2_X1 U435 ( .A(G169GAT), .B(G113GAT), .ZN(n374) );
  XNOR2_X1 U436 ( .A(n375), .B(n374), .ZN(n379) );
  XOR2_X1 U437 ( .A(KEYINPUT65), .B(KEYINPUT67), .Z(n377) );
  XNOR2_X1 U438 ( .A(KEYINPUT29), .B(KEYINPUT66), .ZN(n376) );
  XNOR2_X1 U439 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U440 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U441 ( .A(n381), .B(n380), .ZN(n383) );
  XOR2_X1 U442 ( .A(n383), .B(n382), .Z(n495) );
  NAND2_X1 U443 ( .A1(n529), .A2(n495), .ZN(n385) );
  XOR2_X1 U444 ( .A(G155GAT), .B(G78GAT), .Z(n387) );
  XNOR2_X1 U445 ( .A(G22GAT), .B(G127GAT), .ZN(n386) );
  XNOR2_X1 U446 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U447 ( .A(n389), .B(n388), .Z(n391) );
  NAND2_X1 U448 ( .A1(G231GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U449 ( .A(n391), .B(n390), .ZN(n403) );
  XOR2_X1 U450 ( .A(KEYINPUT80), .B(KEYINPUT78), .Z(n393) );
  XNOR2_X1 U451 ( .A(KEYINPUT15), .B(KEYINPUT12), .ZN(n392) );
  XNOR2_X1 U452 ( .A(n393), .B(n392), .ZN(n397) );
  XOR2_X1 U453 ( .A(KEYINPUT79), .B(KEYINPUT14), .Z(n395) );
  XNOR2_X1 U454 ( .A(G64GAT), .B(KEYINPUT77), .ZN(n394) );
  XNOR2_X1 U455 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U456 ( .A(n397), .B(n396), .Z(n401) );
  XNOR2_X1 U457 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U458 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U459 ( .A(n403), .B(n402), .ZN(n577) );
  XOR2_X1 U460 ( .A(n577), .B(KEYINPUT111), .Z(n562) );
  INV_X1 U461 ( .A(n562), .ZN(n404) );
  NOR2_X1 U462 ( .A1(n535), .A2(n404), .ZN(n405) );
  NAND2_X1 U463 ( .A1(n406), .A2(n405), .ZN(n407) );
  XNOR2_X1 U464 ( .A(n407), .B(KEYINPUT47), .ZN(n412) );
  XOR2_X1 U465 ( .A(KEYINPUT36), .B(n535), .Z(n580) );
  NOR2_X1 U466 ( .A1(n580), .A2(n577), .ZN(n408) );
  XNOR2_X1 U467 ( .A(n408), .B(KEYINPUT45), .ZN(n409) );
  NAND2_X1 U468 ( .A1(n409), .A2(n573), .ZN(n410) );
  INV_X1 U469 ( .A(n495), .ZN(n569) );
  XOR2_X1 U470 ( .A(n569), .B(KEYINPUT68), .Z(n550) );
  NOR2_X1 U471 ( .A1(n410), .A2(n550), .ZN(n411) );
  XNOR2_X1 U472 ( .A(KEYINPUT48), .B(n413), .ZN(n523) );
  NOR2_X1 U473 ( .A1(n414), .A2(n523), .ZN(n415) );
  XOR2_X1 U474 ( .A(KEYINPUT54), .B(n415), .Z(n416) );
  XOR2_X1 U475 ( .A(KEYINPUT87), .B(KEYINPUT24), .Z(n418) );
  XNOR2_X1 U476 ( .A(G50GAT), .B(KEYINPUT23), .ZN(n417) );
  XNOR2_X1 U477 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U478 ( .A(n420), .B(n419), .Z(n422) );
  NAND2_X1 U479 ( .A1(G228GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U480 ( .A(n422), .B(n421), .ZN(n426) );
  XOR2_X1 U481 ( .A(G211GAT), .B(KEYINPUT88), .Z(n424) );
  XNOR2_X1 U482 ( .A(KEYINPUT22), .B(KEYINPUT86), .ZN(n423) );
  XNOR2_X1 U483 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U484 ( .A(n426), .B(n425), .Z(n430) );
  XNOR2_X1 U485 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U486 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U487 ( .A(n432), .B(n431), .ZN(n464) );
  NAND2_X1 U488 ( .A1(n567), .A2(n464), .ZN(n433) );
  XNOR2_X1 U489 ( .A(KEYINPUT55), .B(n433), .ZN(n448) );
  XOR2_X1 U490 ( .A(G71GAT), .B(G176GAT), .Z(n435) );
  XNOR2_X1 U491 ( .A(G15GAT), .B(G99GAT), .ZN(n434) );
  XNOR2_X1 U492 ( .A(n435), .B(n434), .ZN(n437) );
  XOR2_X1 U493 ( .A(G43GAT), .B(G190GAT), .Z(n436) );
  XNOR2_X1 U494 ( .A(n437), .B(n436), .ZN(n445) );
  XNOR2_X1 U495 ( .A(n439), .B(n438), .ZN(n443) );
  XOR2_X1 U496 ( .A(G183GAT), .B(KEYINPUT20), .Z(n441) );
  XNOR2_X1 U497 ( .A(KEYINPUT81), .B(KEYINPUT83), .ZN(n440) );
  XNOR2_X1 U498 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U499 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U500 ( .A(n445), .B(n444), .ZN(n447) );
  NAND2_X1 U501 ( .A1(G227GAT), .A2(G233GAT), .ZN(n446) );
  NAND2_X1 U502 ( .A1(n448), .A2(n524), .ZN(n561) );
  NOR2_X1 U503 ( .A1(n548), .A2(n561), .ZN(n452) );
  XNOR2_X1 U504 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n450) );
  INV_X1 U505 ( .A(G190GAT), .ZN(n449) );
  NAND2_X1 U506 ( .A1(n550), .A2(n573), .ZN(n481) );
  NOR2_X1 U507 ( .A1(n535), .A2(n577), .ZN(n453) );
  XNOR2_X1 U508 ( .A(n453), .B(KEYINPUT16), .ZN(n469) );
  NAND2_X1 U509 ( .A1(n513), .A2(n524), .ZN(n454) );
  NAND2_X1 U510 ( .A1(n454), .A2(n464), .ZN(n456) );
  XNOR2_X1 U511 ( .A(n513), .B(KEYINPUT27), .ZN(n463) );
  NOR2_X1 U512 ( .A1(n524), .A2(n464), .ZN(n458) );
  XNOR2_X1 U513 ( .A(KEYINPUT94), .B(KEYINPUT26), .ZN(n457) );
  XNOR2_X1 U514 ( .A(n458), .B(n457), .ZN(n566) );
  NAND2_X1 U515 ( .A1(n463), .A2(n566), .ZN(n459) );
  NAND2_X1 U516 ( .A1(n460), .A2(n459), .ZN(n461) );
  XOR2_X1 U517 ( .A(KEYINPUT96), .B(n461), .Z(n462) );
  NOR2_X1 U518 ( .A1(n509), .A2(n462), .ZN(n467) );
  NAND2_X1 U519 ( .A1(n509), .A2(n463), .ZN(n522) );
  OR2_X1 U520 ( .A1(n522), .A2(n527), .ZN(n465) );
  NOR2_X1 U521 ( .A1(n524), .A2(n465), .ZN(n466) );
  NOR2_X1 U522 ( .A1(n467), .A2(n466), .ZN(n478) );
  INV_X1 U523 ( .A(n478), .ZN(n468) );
  NAND2_X1 U524 ( .A1(n469), .A2(n468), .ZN(n497) );
  NOR2_X1 U525 ( .A1(n481), .A2(n497), .ZN(n476) );
  NAND2_X1 U526 ( .A1(n509), .A2(n476), .ZN(n472) );
  XOR2_X1 U527 ( .A(G1GAT), .B(KEYINPUT34), .Z(n470) );
  XNOR2_X1 U528 ( .A(KEYINPUT97), .B(n470), .ZN(n471) );
  XNOR2_X1 U529 ( .A(n472), .B(n471), .ZN(G1324GAT) );
  NAND2_X1 U530 ( .A1(n513), .A2(n476), .ZN(n473) );
  XNOR2_X1 U531 ( .A(n473), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U532 ( .A(G15GAT), .B(KEYINPUT35), .Z(n475) );
  NAND2_X1 U533 ( .A1(n476), .A2(n524), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n475), .B(n474), .ZN(G1326GAT) );
  NAND2_X1 U535 ( .A1(n527), .A2(n476), .ZN(n477) );
  XNOR2_X1 U536 ( .A(n477), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U537 ( .A(KEYINPUT98), .B(KEYINPUT39), .Z(n484) );
  NOR2_X1 U538 ( .A1(n580), .A2(n478), .ZN(n479) );
  NAND2_X1 U539 ( .A1(n479), .A2(n577), .ZN(n480) );
  XOR2_X1 U540 ( .A(KEYINPUT37), .B(n480), .Z(n508) );
  NOR2_X1 U541 ( .A1(n508), .A2(n481), .ZN(n482) );
  XNOR2_X1 U542 ( .A(KEYINPUT38), .B(n482), .ZN(n492) );
  NAND2_X1 U543 ( .A1(n492), .A2(n509), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U545 ( .A(G29GAT), .B(n485), .ZN(G1328GAT) );
  XOR2_X1 U546 ( .A(G36GAT), .B(KEYINPUT99), .Z(n487) );
  NAND2_X1 U547 ( .A1(n492), .A2(n513), .ZN(n486) );
  XNOR2_X1 U548 ( .A(n487), .B(n486), .ZN(G1329GAT) );
  XNOR2_X1 U549 ( .A(G43GAT), .B(KEYINPUT101), .ZN(n491) );
  NAND2_X1 U550 ( .A1(n492), .A2(n524), .ZN(n489) );
  XOR2_X1 U551 ( .A(KEYINPUT40), .B(KEYINPUT100), .Z(n488) );
  XNOR2_X1 U552 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n491), .B(n490), .ZN(G1330GAT) );
  XNOR2_X1 U554 ( .A(G50GAT), .B(KEYINPUT102), .ZN(n494) );
  NAND2_X1 U555 ( .A1(n527), .A2(n492), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n494), .B(n493), .ZN(G1331GAT) );
  XNOR2_X1 U557 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n499) );
  INV_X1 U558 ( .A(n529), .ZN(n553) );
  NOR2_X1 U559 ( .A1(n495), .A2(n553), .ZN(n496) );
  XNOR2_X1 U560 ( .A(n496), .B(KEYINPUT103), .ZN(n507) );
  NOR2_X1 U561 ( .A1(n507), .A2(n497), .ZN(n504) );
  NAND2_X1 U562 ( .A1(n504), .A2(n509), .ZN(n498) );
  XNOR2_X1 U563 ( .A(n499), .B(n498), .ZN(G1332GAT) );
  NAND2_X1 U564 ( .A1(n513), .A2(n504), .ZN(n500) );
  XNOR2_X1 U565 ( .A(n500), .B(KEYINPUT104), .ZN(n501) );
  XNOR2_X1 U566 ( .A(G64GAT), .B(n501), .ZN(G1333GAT) );
  XOR2_X1 U567 ( .A(G71GAT), .B(KEYINPUT105), .Z(n503) );
  NAND2_X1 U568 ( .A1(n504), .A2(n524), .ZN(n502) );
  XNOR2_X1 U569 ( .A(n503), .B(n502), .ZN(G1334GAT) );
  XOR2_X1 U570 ( .A(G78GAT), .B(KEYINPUT43), .Z(n506) );
  NAND2_X1 U571 ( .A1(n504), .A2(n527), .ZN(n505) );
  XNOR2_X1 U572 ( .A(n506), .B(n505), .ZN(G1335GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n511) );
  NOR2_X1 U574 ( .A1(n508), .A2(n507), .ZN(n519) );
  NAND2_X1 U575 ( .A1(n519), .A2(n509), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U577 ( .A(G85GAT), .B(n512), .ZN(G1336GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n515) );
  NAND2_X1 U579 ( .A1(n519), .A2(n513), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U581 ( .A(G92GAT), .B(n516), .ZN(G1337GAT) );
  NAND2_X1 U582 ( .A1(n519), .A2(n524), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n517), .B(KEYINPUT110), .ZN(n518) );
  XNOR2_X1 U584 ( .A(G99GAT), .B(n518), .ZN(G1338GAT) );
  NAND2_X1 U585 ( .A1(n527), .A2(n519), .ZN(n520) );
  XNOR2_X1 U586 ( .A(n520), .B(KEYINPUT44), .ZN(n521) );
  XNOR2_X1 U587 ( .A(G106GAT), .B(n521), .ZN(G1339GAT) );
  NOR2_X1 U588 ( .A1(n523), .A2(n522), .ZN(n539) );
  NAND2_X1 U589 ( .A1(n524), .A2(n539), .ZN(n525) );
  XOR2_X1 U590 ( .A(KEYINPUT113), .B(n525), .Z(n526) );
  NOR2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n536) );
  NAND2_X1 U592 ( .A1(n536), .A2(n550), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n528), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U594 ( .A(G120GAT), .B(KEYINPUT49), .Z(n531) );
  NAND2_X1 U595 ( .A1(n536), .A2(n529), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(G1341GAT) );
  INV_X1 U597 ( .A(n536), .ZN(n532) );
  NOR2_X1 U598 ( .A1(n562), .A2(n532), .ZN(n533) );
  XOR2_X1 U599 ( .A(KEYINPUT50), .B(n533), .Z(n534) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(n534), .ZN(G1342GAT) );
  XOR2_X1 U601 ( .A(G134GAT), .B(KEYINPUT51), .Z(n538) );
  NAND2_X1 U602 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n538), .B(n537), .ZN(G1343GAT) );
  NAND2_X1 U604 ( .A1(n566), .A2(n539), .ZN(n547) );
  NOR2_X1 U605 ( .A1(n569), .A2(n547), .ZN(n540) );
  XOR2_X1 U606 ( .A(G141GAT), .B(n540), .Z(G1344GAT) );
  NOR2_X1 U607 ( .A1(n553), .A2(n547), .ZN(n545) );
  XOR2_X1 U608 ( .A(KEYINPUT53), .B(KEYINPUT115), .Z(n542) );
  XNOR2_X1 U609 ( .A(G148GAT), .B(KEYINPUT114), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U611 ( .A(KEYINPUT52), .B(n543), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(G1345GAT) );
  NOR2_X1 U613 ( .A1(n577), .A2(n547), .ZN(n546) );
  XOR2_X1 U614 ( .A(G155GAT), .B(n546), .Z(G1346GAT) );
  NOR2_X1 U615 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U616 ( .A(G162GAT), .B(n549), .Z(G1347GAT) );
  INV_X1 U617 ( .A(n550), .ZN(n551) );
  NOR2_X1 U618 ( .A1(n551), .A2(n561), .ZN(n552) );
  XOR2_X1 U619 ( .A(G169GAT), .B(n552), .Z(G1348GAT) );
  NOR2_X1 U620 ( .A1(n561), .A2(n553), .ZN(n560) );
  XOR2_X1 U621 ( .A(KEYINPUT56), .B(KEYINPUT118), .Z(n555) );
  XNOR2_X1 U622 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U624 ( .A(n556), .B(KEYINPUT119), .Z(n558) );
  XNOR2_X1 U625 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1349GAT) );
  NOR2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n564) );
  XNOR2_X1 U629 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U633 ( .A(KEYINPUT123), .B(n568), .Z(n579) );
  NOR2_X1 U634 ( .A1(n569), .A2(n579), .ZN(n571) );
  XNOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(n572), .ZN(G1352GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n579), .ZN(n575) );
  XNOR2_X1 U639 ( .A(KEYINPUT124), .B(KEYINPUT61), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(G204GAT), .B(n576), .ZN(G1353GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n579), .ZN(n578) );
  XOR2_X1 U643 ( .A(G211GAT), .B(n578), .Z(G1354GAT) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n585) );
  XOR2_X1 U645 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(KEYINPUT125), .B(n583), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(G1355GAT) );
endmodule

