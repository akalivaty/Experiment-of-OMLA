//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 1 1 0 0 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1 1 1 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 1 1 1 1 0 0 1 1 0 1 0 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055;
  XNOR2_X1  g000(.A(G113), .B(G122), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n187), .B(new_n188), .ZN(new_n189));
  NOR2_X1   g003(.A1(G237), .A2(G953), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G214), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(G143), .A3(G214), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT18), .A2(G131), .ZN(new_n195));
  AND3_X1   g009(.A1(new_n193), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n195), .B1(new_n193), .B2(new_n194), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G140), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(KEYINPUT75), .A3(G125), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(G125), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G140), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  OAI211_X1 g018(.A(G146), .B(new_n200), .C1(new_n204), .C2(KEYINPUT75), .ZN(new_n205));
  AND2_X1   g019(.A1(new_n201), .A2(new_n203), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  AND3_X1   g022(.A1(new_n205), .A2(KEYINPUT84), .A3(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(KEYINPUT84), .B1(new_n205), .B2(new_n208), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n198), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT85), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT85), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n213), .B(new_n198), .C1(new_n209), .C2(new_n210), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  OAI211_X1 g029(.A(KEYINPUT16), .B(new_n200), .C1(new_n204), .C2(KEYINPUT75), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT16), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n201), .A2(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n207), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G131), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n221), .B1(new_n193), .B2(new_n194), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n193), .A2(new_n221), .A3(new_n194), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n206), .A2(KEYINPUT19), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n200), .B1(new_n204), .B2(KEYINPUT75), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n224), .B1(new_n225), .B2(KEYINPUT19), .ZN(new_n226));
  OAI221_X1 g040(.A(new_n220), .B1(new_n222), .B2(new_n223), .C1(new_n226), .C2(G146), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n189), .B1(new_n215), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT86), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n216), .A2(new_n207), .A3(new_n218), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT76), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT76), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n216), .A2(new_n233), .A3(new_n207), .A4(new_n218), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n232), .A2(new_n220), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT17), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n236), .B1(new_n223), .B2(new_n222), .ZN(new_n237));
  OR2_X1    g051(.A1(new_n222), .A2(new_n236), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AOI22_X1  g053(.A1(new_n214), .A2(new_n212), .B1(new_n235), .B2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n230), .B1(new_n240), .B2(new_n189), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n219), .B1(KEYINPUT76), .B2(new_n231), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(new_n239), .A3(new_n234), .ZN(new_n243));
  AND4_X1   g057(.A1(new_n230), .A2(new_n215), .A3(new_n189), .A4(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n229), .B1(new_n241), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT20), .ZN(new_n246));
  NOR2_X1   g060(.A1(G475), .A2(G902), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n205), .A2(new_n208), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT84), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n205), .A2(KEYINPUT84), .A3(new_n208), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n213), .B1(new_n253), .B2(new_n198), .ZN(new_n254));
  INV_X1    g068(.A(new_n214), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n189), .B(new_n243), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(KEYINPUT86), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n215), .A2(new_n230), .A3(new_n189), .A4(new_n243), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n228), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n247), .ZN(new_n260));
  OAI21_X1  g074(.A(KEYINPUT20), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n248), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G128), .ZN(new_n263));
  AOI21_X1  g077(.A(KEYINPUT13), .B1(new_n263), .B2(G143), .ZN(new_n264));
  INV_X1    g078(.A(G134), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(G128), .B(G143), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n266), .B(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G122), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n269), .A2(KEYINPUT87), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(KEYINPUT87), .ZN(new_n271));
  OAI21_X1  g085(.A(G116), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G107), .ZN(new_n273));
  INV_X1    g087(.A(G116), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G122), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n272), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n273), .B1(new_n272), .B2(new_n275), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n268), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n272), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n275), .B(KEYINPUT14), .ZN(new_n281));
  OAI21_X1  g095(.A(G107), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n267), .B(new_n265), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(new_n276), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n279), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g099(.A(KEYINPUT9), .B(G234), .ZN(new_n286));
  INV_X1    g100(.A(G217), .ZN(new_n287));
  NOR3_X1   g101(.A1(new_n286), .A2(new_n287), .A3(G953), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n285), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n279), .A2(new_n284), .A3(new_n288), .ZN(new_n291));
  AOI21_X1  g105(.A(G902), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G478), .ZN(new_n293));
  NOR2_X1   g107(.A1(KEYINPUT88), .A2(KEYINPUT15), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(KEYINPUT88), .A2(KEYINPUT15), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n293), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  OR2_X1    g112(.A1(new_n292), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n292), .A2(new_n298), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n240), .A2(new_n189), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n303), .B1(new_n258), .B2(new_n257), .ZN(new_n304));
  OAI21_X1  g118(.A(G475), .B1(new_n304), .B2(G902), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n262), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT11), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n307), .B1(new_n265), .B2(G137), .ZN(new_n308));
  INV_X1    g122(.A(G137), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(KEYINPUT11), .A3(G134), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n265), .A2(G137), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n308), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G131), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n308), .A2(new_n310), .A3(new_n221), .A4(new_n311), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n207), .A2(G143), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n192), .A2(G146), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n207), .A2(G143), .ZN(new_n319));
  AOI22_X1  g133(.A1(new_n318), .A2(new_n263), .B1(KEYINPUT1), .B2(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(G143), .B(G146), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT80), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n263), .A2(KEYINPUT1), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(new_n316), .A3(new_n317), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT80), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n320), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT3), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n328), .B1(new_n188), .B2(G107), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n273), .A2(KEYINPUT3), .A3(G104), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G101), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n188), .A2(G107), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT79), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n188), .A2(KEYINPUT79), .A3(G107), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n331), .A2(new_n332), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n333), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n188), .A2(G107), .ZN(new_n339));
  OAI21_X1  g153(.A(G101), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n327), .A2(new_n337), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n319), .A2(KEYINPUT1), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n325), .B(new_n342), .C1(G128), .C2(new_n321), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n343), .B1(new_n337), .B2(new_n340), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n341), .B1(new_n344), .B2(KEYINPUT81), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n337), .A2(new_n340), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n342), .B1(new_n321), .B2(G128), .ZN(new_n347));
  INV_X1    g161(.A(new_n325), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT81), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n315), .B1(new_n345), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT12), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n331), .A2(new_n335), .A3(new_n336), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(G101), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(KEYINPUT4), .A3(new_n337), .ZN(new_n357));
  NAND2_X1  g171(.A1(KEYINPUT0), .A2(G128), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n316), .A2(new_n317), .A3(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n358), .ZN(new_n360));
  NOR2_X1   g174(.A1(KEYINPUT0), .A2(G128), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n359), .B1(new_n362), .B2(new_n321), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT66), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT66), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n359), .B(new_n365), .C1(new_n362), .C2(new_n321), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT4), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n355), .A2(new_n367), .A3(G101), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n357), .A2(new_n364), .A3(new_n366), .A4(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n341), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n315), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n349), .A2(new_n370), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n337), .A2(new_n340), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n369), .A2(new_n371), .A3(new_n372), .A4(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(G110), .B(G140), .ZN(new_n377));
  INV_X1    g191(.A(G953), .ZN(new_n378));
  AND2_X1   g192(.A1(new_n378), .A2(G227), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n377), .B(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT12), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n382), .B(new_n315), .C1(new_n345), .C2(new_n352), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n354), .A2(new_n376), .A3(new_n381), .A4(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n376), .ZN(new_n385));
  AOI22_X1  g199(.A1(new_n341), .A2(new_n370), .B1(new_n373), .B2(new_n374), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n372), .B1(new_n386), .B2(new_n369), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n380), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n384), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G469), .ZN(new_n390));
  INV_X1    g204(.A(G902), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n390), .A2(new_n391), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  AOI22_X1  g208(.A1(new_n350), .A2(new_n351), .B1(new_n374), .B2(new_n327), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n344), .A2(KEYINPUT81), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n372), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n376), .B1(new_n397), .B2(new_n382), .ZN(new_n398));
  INV_X1    g212(.A(new_n383), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n380), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n371), .A2(new_n375), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n335), .A2(new_n336), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n332), .B1(new_n402), .B2(new_n331), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n337), .A2(KEYINPUT4), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n368), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n364), .A2(new_n366), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n315), .B1(new_n401), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(new_n376), .A3(new_n381), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n400), .A2(G469), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n392), .A2(new_n394), .A3(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G221), .ZN(new_n412));
  INV_X1    g226(.A(new_n286), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n412), .B1(new_n413), .B2(new_n391), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(G214), .B1(G237), .B2(G902), .ZN(new_n417));
  NAND2_X1  g231(.A1(G234), .A2(G237), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(G952), .A3(new_n378), .ZN(new_n419));
  XNOR2_X1  g233(.A(KEYINPUT21), .B(G898), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n418), .A2(G902), .A3(G953), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n419), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(G110), .B(G122), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  XOR2_X1   g239(.A(KEYINPUT2), .B(G113), .Z(new_n426));
  XNOR2_X1  g240(.A(G116), .B(G119), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(KEYINPUT2), .B(G113), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n274), .A2(G119), .ZN(new_n430));
  INV_X1    g244(.A(G119), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n431), .A2(G116), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n429), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n428), .A2(new_n433), .A3(KEYINPUT65), .ZN(new_n434));
  OR3_X1    g248(.A1(new_n426), .A2(KEYINPUT65), .A3(new_n427), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n405), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n427), .A2(KEYINPUT5), .ZN(new_n438));
  INV_X1    g252(.A(G113), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT5), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n439), .B1(new_n430), .B2(new_n440), .ZN(new_n441));
  AOI22_X1  g255(.A1(new_n438), .A2(new_n441), .B1(new_n426), .B2(new_n427), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n442), .A2(new_n337), .A3(new_n340), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT82), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n374), .A2(KEYINPUT82), .A3(new_n442), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n425), .B1(new_n437), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n436), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(new_n368), .A3(new_n357), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n450), .A2(new_n424), .A3(new_n445), .A4(new_n446), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n448), .A2(KEYINPUT6), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n363), .A2(G125), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n453), .B1(new_n349), .B2(G125), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n378), .A2(G224), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(KEYINPUT83), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n454), .B(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n458), .B(new_n425), .C1(new_n437), .C2(new_n447), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n452), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(G210), .B1(G237), .B2(G902), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n455), .A2(KEYINPUT7), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n454), .B(new_n462), .ZN(new_n463));
  XOR2_X1   g277(.A(new_n424), .B(KEYINPUT8), .Z(new_n464));
  OR2_X1    g278(.A1(new_n374), .A2(new_n442), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n464), .B1(new_n465), .B2(new_n443), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(G902), .B1(new_n467), .B2(new_n451), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n460), .A2(new_n461), .A3(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n461), .B1(new_n460), .B2(new_n468), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n417), .B(new_n423), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  NOR3_X1   g286(.A1(new_n306), .A2(new_n416), .A3(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT22), .B(G137), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n378), .A2(G221), .A3(G234), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n474), .B(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n263), .A2(G119), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n431), .A2(G128), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  XOR2_X1   g294(.A(KEYINPUT24), .B(G110), .Z(new_n481));
  NAND3_X1  g295(.A1(new_n480), .A2(new_n481), .A3(KEYINPUT74), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT74), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT24), .B(G110), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n483), .B1(new_n479), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n263), .A2(KEYINPUT23), .A3(G119), .ZN(new_n487));
  INV_X1    g301(.A(new_n477), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n487), .B(new_n478), .C1(new_n488), .C2(KEYINPUT23), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(G110), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n491), .B1(new_n242), .B2(new_n234), .ZN(new_n492));
  OAI22_X1  g306(.A1(new_n489), .A2(G110), .B1(new_n480), .B2(new_n481), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n220), .A2(new_n208), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n476), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n232), .A2(new_n220), .A3(new_n234), .ZN(new_n497));
  INV_X1    g311(.A(new_n491), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n476), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n494), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n496), .A2(new_n391), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(KEYINPUT25), .B1(new_n502), .B2(KEYINPUT77), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT77), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n496), .A2(new_n504), .A3(new_n501), .A4(new_n391), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n503), .A2(KEYINPUT78), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n287), .B1(G234), .B2(new_n391), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n502), .A2(KEYINPUT77), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT25), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n511), .A3(new_n505), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT78), .ZN(new_n513));
  OR2_X1    g327(.A1(new_n502), .A2(new_n511), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n496), .A2(new_n501), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n507), .A2(G902), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n509), .A2(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT73), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n265), .A2(G137), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n309), .A2(G134), .ZN(new_n522));
  OAI21_X1  g336(.A(G131), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AND2_X1   g337(.A1(new_n314), .A2(new_n523), .ZN(new_n524));
  AOI22_X1  g338(.A1(new_n315), .A2(new_n363), .B1(new_n524), .B2(new_n343), .ZN(new_n525));
  OAI21_X1  g339(.A(KEYINPUT64), .B1(new_n525), .B2(KEYINPUT30), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n315), .A2(new_n363), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n524), .A2(new_n343), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT64), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT30), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n526), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n314), .A2(new_n523), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT67), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n314), .A2(new_n523), .A3(KEYINPUT67), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(new_n537), .A3(new_n343), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT68), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI22_X1  g354(.A1(new_n534), .A2(new_n535), .B1(new_n320), .B2(new_n325), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n541), .A2(KEYINPUT68), .A3(new_n537), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n364), .A2(new_n315), .A3(new_n366), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n540), .A2(KEYINPUT30), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n533), .A2(new_n449), .A3(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(KEYINPUT26), .B(G101), .ZN(new_n546));
  XNOR2_X1  g360(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n546), .B(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n190), .A2(G210), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n549), .B(KEYINPUT70), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n548), .B(new_n550), .ZN(new_n551));
  AND4_X1   g365(.A1(KEYINPUT68), .A2(new_n536), .A3(new_n537), .A4(new_n343), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT68), .B1(new_n541), .B2(new_n537), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n543), .A2(new_n436), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n551), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT31), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n545), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(KEYINPUT71), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT71), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n545), .A2(new_n557), .A3(new_n561), .A4(new_n558), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n551), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n553), .A2(new_n552), .A3(new_n555), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n525), .A2(new_n436), .ZN(new_n566));
  OAI21_X1  g380(.A(KEYINPUT28), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n538), .A2(new_n543), .A3(new_n436), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT28), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n568), .A2(KEYINPUT72), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(KEYINPUT72), .B1(new_n568), .B2(new_n569), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n564), .B1(new_n567), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n558), .B1(new_n545), .B2(new_n557), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n563), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(G472), .A2(G902), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n520), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n577), .ZN(new_n579));
  AOI211_X1 g393(.A(KEYINPUT73), .B(new_n579), .C1(new_n563), .C2(new_n575), .ZN(new_n580));
  NOR3_X1   g394(.A1(new_n578), .A2(new_n580), .A3(KEYINPUT32), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT29), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n556), .A2(new_n540), .A3(new_n542), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n545), .A2(new_n582), .A3(new_n551), .A4(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n567), .A2(new_n572), .A3(new_n582), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n564), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n449), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n583), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(KEYINPUT28), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n582), .B1(new_n590), .B2(new_n572), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n391), .B(new_n584), .C1(new_n586), .C2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(G472), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n576), .A2(KEYINPUT32), .A3(new_n577), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n473), .B(new_n519), .C1(new_n581), .C2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(G101), .ZN(G3));
  NAND2_X1  g411(.A1(new_n576), .A2(new_n391), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n598), .A2(KEYINPUT89), .A3(G472), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT89), .ZN(new_n600));
  AOI21_X1  g414(.A(G902), .B1(new_n563), .B2(new_n575), .ZN(new_n601));
  INV_X1    g415(.A(G472), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n578), .A2(new_n580), .ZN(new_n605));
  AOI21_X1  g419(.A(G902), .B1(new_n384), .B2(new_n388), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n393), .B1(new_n606), .B2(new_n390), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n414), .B1(new_n607), .B2(new_n410), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n604), .A2(new_n605), .A3(new_n519), .A4(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n246), .B1(new_n245), .B2(new_n247), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n259), .A2(KEYINPUT20), .A3(new_n260), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n305), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n460), .A2(new_n468), .ZN(new_n614));
  INV_X1    g428(.A(new_n461), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n616), .A2(KEYINPUT90), .A3(new_n469), .ZN(new_n617));
  INV_X1    g431(.A(new_n417), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT90), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n618), .B1(new_n471), .B2(new_n619), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n290), .A2(new_n291), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT91), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n290), .B(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT92), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n623), .B1(new_n291), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n628), .B1(new_n627), .B2(new_n291), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n624), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n293), .A2(G902), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  OAI22_X1  g446(.A1(new_n630), .A2(new_n632), .B1(G478), .B2(new_n292), .ZN(new_n633));
  AND4_X1   g447(.A1(new_n613), .A2(new_n621), .A3(new_n423), .A4(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n610), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT34), .B(G104), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G6));
  AND2_X1   g451(.A1(new_n621), .A2(new_n423), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n257), .A2(new_n258), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n391), .B1(new_n639), .B2(new_n303), .ZN(new_n640));
  AOI22_X1  g454(.A1(new_n248), .A2(new_n261), .B1(new_n640), .B2(G475), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n301), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n610), .A2(new_n638), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT35), .B(G107), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G9));
  NAND3_X1  g460(.A1(new_n604), .A2(new_n605), .A3(new_n608), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n499), .A2(new_n494), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n476), .A2(KEYINPUT36), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(new_n650));
  AND3_X1   g464(.A1(new_n650), .A2(KEYINPUT93), .A3(new_n518), .ZN(new_n651));
  AOI21_X1  g465(.A(KEYINPUT93), .B1(new_n650), .B2(new_n518), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n513), .B1(new_n502), .B2(new_n511), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n654), .B1(new_n505), .B2(new_n503), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n653), .B1(new_n508), .B2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT94), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n306), .ZN(new_n659));
  INV_X1    g473(.A(new_n472), .ZN(new_n660));
  OAI211_X1 g474(.A(KEYINPUT94), .B(new_n653), .C1(new_n508), .C2(new_n655), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n658), .A2(new_n659), .A3(new_n660), .A4(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n647), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT95), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT37), .B(G110), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G12));
  NAND3_X1  g480(.A1(new_n515), .A2(new_n506), .A3(new_n507), .ZN(new_n667));
  AOI21_X1  g481(.A(KEYINPUT94), .B1(new_n667), .B2(new_n653), .ZN(new_n668));
  INV_X1    g482(.A(new_n661), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n576), .A2(new_n577), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(KEYINPUT73), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT32), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n576), .A2(new_n520), .A3(new_n577), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n593), .A2(new_n594), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n670), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n617), .A2(new_n620), .A3(new_n411), .A4(new_n415), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n419), .B1(new_n422), .B2(G900), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n680), .B(KEYINPUT96), .Z(new_n681));
  NOR3_X1   g495(.A1(new_n642), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G128), .ZN(G30));
  INV_X1    g498(.A(KEYINPUT40), .ZN(new_n685));
  XOR2_X1   g499(.A(new_n681), .B(KEYINPUT39), .Z(new_n686));
  NAND3_X1  g500(.A1(new_n608), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n689), .B1(new_n470), .B2(new_n471), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n616), .A2(new_n469), .A3(new_n688), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n618), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n302), .B1(new_n262), .B2(new_n305), .ZN(new_n693));
  AND3_X1   g507(.A1(new_n687), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n391), .B1(new_n589), .B2(new_n564), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n551), .B1(new_n545), .B2(new_n583), .ZN(new_n696));
  OAI21_X1  g510(.A(G472), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n594), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n675), .A2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n656), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n608), .A2(new_n686), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(KEYINPUT40), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n694), .A2(new_n699), .A3(new_n700), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G143), .ZN(G45));
  INV_X1    g518(.A(new_n681), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n613), .A2(new_n633), .A3(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n706), .A2(new_n679), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n678), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G146), .ZN(G48));
  NAND2_X1  g523(.A1(new_n389), .A2(new_n391), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(G469), .ZN(new_n711));
  AOI21_X1  g525(.A(KEYINPUT98), .B1(new_n606), .B2(new_n390), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n710), .A2(KEYINPUT98), .A3(G469), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(KEYINPUT99), .B1(new_n715), .B2(new_n415), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT99), .ZN(new_n717));
  AOI211_X1 g531(.A(new_n717), .B(new_n414), .C1(new_n713), .C2(new_n714), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n517), .A2(new_n518), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n667), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n721), .B1(new_n675), .B2(new_n676), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n719), .A2(new_n722), .A3(new_n634), .ZN(new_n723));
  XNOR2_X1  g537(.A(KEYINPUT41), .B(G113), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G15));
  AND4_X1   g539(.A1(new_n722), .A2(new_n719), .A3(new_n638), .A4(new_n643), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(new_n274), .ZN(G18));
  NAND2_X1  g541(.A1(new_n719), .A2(new_n638), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n670), .A2(new_n677), .A3(new_n659), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(new_n431), .ZN(G21));
  AND2_X1   g545(.A1(new_n560), .A2(new_n562), .ZN(new_n732));
  INV_X1    g546(.A(new_n572), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n569), .B1(new_n588), .B2(new_n583), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n551), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n574), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n577), .B1(new_n732), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT100), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n598), .A2(G472), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT100), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n742), .B(new_n577), .C1(new_n732), .C2(new_n737), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n741), .A2(new_n519), .A3(new_n693), .A4(new_n743), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n728), .A2(new_n744), .ZN(new_n745));
  XOR2_X1   g559(.A(KEYINPUT101), .B(G122), .Z(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(G24));
  NAND4_X1  g561(.A1(new_n739), .A2(new_n740), .A3(new_n656), .A4(new_n743), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n748), .A2(new_n706), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(new_n719), .A3(new_n621), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G125), .ZN(G27));
  AOI21_X1  g565(.A(KEYINPUT32), .B1(new_n576), .B2(new_n577), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n519), .B1(new_n595), .B2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n616), .A2(new_n469), .A3(new_n417), .ZN(new_n755));
  OR2_X1    g569(.A1(new_n755), .A2(new_n414), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n400), .A2(KEYINPUT102), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT102), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n758), .B(new_n380), .C1(new_n398), .C2(new_n399), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n757), .A2(G469), .A3(new_n409), .A4(new_n759), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n607), .B1(new_n760), .B2(KEYINPUT103), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT103), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n759), .A2(new_n409), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n354), .A2(new_n376), .A3(new_n383), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n758), .B1(new_n764), .B2(new_n380), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n762), .B1(new_n766), .B2(G469), .ZN(new_n767));
  OAI21_X1  g581(.A(KEYINPUT104), .B1(new_n761), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n766), .A2(new_n762), .A3(G469), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n760), .A2(KEYINPUT103), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT104), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n769), .A2(new_n770), .A3(new_n771), .A4(new_n607), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n756), .B1(new_n768), .B2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n706), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n754), .A2(KEYINPUT42), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n722), .A2(new_n773), .A3(new_n774), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT42), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n776), .A2(KEYINPUT105), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT105), .B1(new_n776), .B2(new_n777), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n775), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G131), .ZN(G33));
  NOR2_X1   g595(.A1(new_n642), .A2(new_n681), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n722), .A2(new_n773), .A3(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G134), .ZN(G36));
  AOI21_X1  g598(.A(new_n700), .B1(new_n604), .B2(new_n605), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT43), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n786), .B1(new_n641), .B2(new_n633), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n305), .B(new_n633), .C1(new_n611), .C2(new_n612), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(KEYINPUT43), .ZN(new_n789));
  OAI21_X1  g603(.A(KEYINPUT107), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n641), .A2(new_n786), .A3(new_n633), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n788), .A2(KEYINPUT43), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT107), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n785), .A2(new_n790), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT44), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n755), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n400), .A2(new_n409), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT45), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n390), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n757), .A2(KEYINPUT45), .A3(new_n409), .A4(new_n759), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n393), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n392), .B1(new_n802), .B2(KEYINPUT46), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT46), .ZN(new_n804));
  AOI211_X1 g618(.A(new_n804), .B(new_n393), .C1(new_n800), .C2(new_n801), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n415), .B(new_n686), .C1(new_n803), .C2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT106), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n763), .A2(new_n765), .A3(new_n799), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n385), .A2(new_n387), .A3(new_n380), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n810), .B1(new_n380), .B2(new_n764), .ZN(new_n811));
  OAI21_X1  g625(.A(G469), .B1(new_n811), .B2(KEYINPUT45), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n394), .B1(new_n809), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(new_n804), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n802), .A2(KEYINPUT46), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n814), .A2(new_n392), .A3(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n816), .A2(KEYINPUT106), .A3(new_n415), .A4(new_n686), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n808), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n785), .A2(new_n790), .A3(KEYINPUT44), .A4(new_n794), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n797), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G137), .ZN(G39));
  AOI21_X1  g635(.A(new_n755), .B1(new_n667), .B2(new_n720), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n774), .A2(new_n675), .A3(new_n676), .A4(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n415), .B1(new_n803), .B2(new_n805), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT47), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n816), .A2(KEYINPUT47), .A3(new_n415), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n823), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(new_n199), .ZN(G42));
  OAI211_X1 g643(.A(new_n670), .B(new_n677), .C1(new_n682), .C2(new_n707), .ZN(new_n830));
  AND4_X1   g644(.A1(new_n415), .A2(new_n621), .A3(new_n693), .A4(new_n705), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n768), .A2(new_n772), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n831), .A2(new_n699), .A3(new_n832), .A4(new_n700), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n750), .A2(new_n830), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT52), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n750), .A2(new_n830), .A3(new_n833), .A4(KEYINPUT52), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n836), .A2(KEYINPUT109), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT109), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n834), .A2(new_n839), .A3(new_n835), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n723), .B1(new_n728), .B2(new_n744), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n842), .A2(new_n730), .A3(new_n726), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n780), .A2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n596), .B1(new_n647), .B2(new_n662), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n613), .A2(new_n633), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n299), .A2(KEYINPUT108), .A3(new_n300), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT108), .B1(new_n299), .B2(new_n300), .ZN(new_n849));
  OR2_X1    g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n847), .B1(new_n850), .B2(new_n613), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(new_n660), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n852), .A2(new_n609), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n846), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n749), .A2(new_n773), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n705), .B1(new_n848), .B2(new_n849), .ZN(new_n856));
  NOR4_X1   g670(.A1(new_n613), .A2(new_n416), .A3(new_n755), .A4(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n670), .A2(new_n677), .A3(new_n857), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n783), .A2(new_n855), .A3(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT110), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n854), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  OAI221_X1 g675(.A(new_n596), .B1(new_n647), .B2(new_n662), .C1(new_n609), .C2(new_n852), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n783), .A2(new_n855), .A3(new_n858), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT110), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n861), .A2(new_n864), .A3(KEYINPUT53), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n841), .A2(new_n845), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n836), .A2(new_n837), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n862), .A2(new_n863), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n867), .A2(new_n780), .A3(new_n843), .A4(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT53), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XOR2_X1   g685(.A(KEYINPUT111), .B(KEYINPUT54), .Z(new_n872));
  NAND3_X1  g686(.A1(new_n866), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  AND4_X1   g687(.A1(new_n870), .A2(new_n780), .A3(new_n843), .A4(new_n868), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n841), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n869), .A2(KEYINPUT53), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n873), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n378), .A2(G952), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n787), .A2(new_n789), .ZN(new_n881));
  INV_X1    g695(.A(new_n419), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n741), .A2(new_n519), .A3(new_n743), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n719), .A2(new_n621), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n880), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n699), .A2(new_n721), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n716), .A2(new_n718), .A3(new_n755), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n888), .A2(new_n889), .A3(new_n882), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n887), .B1(new_n847), .B2(new_n890), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n889), .A2(new_n882), .A3(new_n881), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n892), .A2(new_n754), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n893), .A2(KEYINPUT114), .A3(KEYINPUT48), .ZN(new_n894));
  XOR2_X1   g708(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n895));
  AOI211_X1 g709(.A(new_n891), .B(new_n894), .C1(new_n893), .C2(new_n895), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n690), .A2(new_n691), .A3(new_n618), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n885), .A2(new_n719), .A3(new_n897), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n898), .B(KEYINPUT50), .Z(new_n899));
  NOR3_X1   g713(.A1(new_n890), .A2(new_n613), .A3(new_n633), .ZN(new_n900));
  INV_X1    g714(.A(new_n748), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n900), .B1(new_n901), .B2(new_n892), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT51), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n883), .A2(new_n884), .A3(new_n755), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n715), .A2(new_n414), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n826), .A2(new_n827), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n903), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n899), .A2(new_n902), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n826), .A2(new_n827), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT112), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n905), .B(KEYINPUT113), .Z(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n909), .A2(KEYINPUT112), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n904), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n899), .A2(new_n914), .A3(new_n902), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n896), .B(new_n908), .C1(KEYINPUT51), .C2(new_n915), .ZN(new_n916));
  OAI22_X1  g730(.A1(new_n879), .A2(new_n916), .B1(G952), .B2(G953), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n690), .A2(new_n691), .A3(new_n415), .A4(new_n417), .ZN(new_n918));
  INV_X1    g732(.A(new_n715), .ZN(new_n919));
  AOI211_X1 g733(.A(new_n788), .B(new_n918), .C1(KEYINPUT49), .C2(new_n919), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n888), .B(new_n920), .C1(KEYINPUT49), .C2(new_n919), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n917), .A2(new_n921), .ZN(G75));
  NOR2_X1   g736(.A1(new_n378), .A2(G952), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(G210), .A2(G902), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n925), .B1(new_n866), .B2(new_n871), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n452), .A2(new_n459), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(new_n457), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT55), .Z(new_n929));
  OR2_X1    g743(.A1(new_n929), .A2(KEYINPUT56), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n924), .B1(new_n926), .B2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT56), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n932), .B1(new_n926), .B2(KEYINPUT115), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n861), .A2(new_n864), .A3(KEYINPUT53), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n934), .A2(new_n844), .ZN(new_n935));
  AOI22_X1  g749(.A1(new_n935), .A2(new_n841), .B1(new_n870), .B2(new_n869), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT115), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n936), .A2(new_n937), .A3(new_n925), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n929), .B1(new_n933), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(KEYINPUT116), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT116), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n941), .B(new_n929), .C1(new_n933), .C2(new_n938), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n931), .B1(new_n940), .B2(new_n942), .ZN(G51));
  XNOR2_X1  g757(.A(new_n393), .B(KEYINPUT57), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n866), .A2(new_n871), .A3(new_n872), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n872), .B1(new_n866), .B2(new_n871), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n389), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n936), .A2(new_n391), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n949), .A2(new_n801), .A3(new_n800), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n923), .B1(new_n948), .B2(new_n950), .ZN(G54));
  NAND3_X1  g765(.A1(new_n949), .A2(KEYINPUT58), .A3(G475), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n952), .A2(new_n259), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n952), .A2(new_n259), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n953), .A2(new_n954), .A3(new_n923), .ZN(G60));
  NAND2_X1  g769(.A1(G478), .A2(G902), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT59), .Z(new_n957));
  NOR2_X1   g771(.A1(new_n630), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n958), .B1(new_n945), .B2(new_n946), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n924), .ZN(new_n960));
  INV_X1    g774(.A(new_n630), .ZN(new_n961));
  INV_X1    g775(.A(new_n957), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n961), .B1(new_n879), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(KEYINPUT117), .B1(new_n960), .B2(new_n963), .ZN(new_n964));
  AOI22_X1  g778(.A1(new_n874), .A2(new_n841), .B1(new_n869), .B2(KEYINPUT53), .ZN(new_n965));
  AOI22_X1  g779(.A1(new_n936), .A2(new_n872), .B1(new_n965), .B2(KEYINPUT54), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n630), .B1(new_n966), .B2(new_n957), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT117), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n967), .A2(new_n968), .A3(new_n924), .A4(new_n959), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n964), .A2(new_n969), .ZN(G63));
  NAND2_X1  g784(.A1(G217), .A2(G902), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT60), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n936), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n650), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n516), .B1(new_n936), .B2(new_n972), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n974), .A2(new_n924), .A3(new_n975), .ZN(new_n976));
  XNOR2_X1  g790(.A(KEYINPUT118), .B(KEYINPUT61), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n976), .B(new_n978), .ZN(G66));
  NAND2_X1  g793(.A1(new_n843), .A2(new_n854), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n378), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n378), .B1(new_n421), .B2(G224), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT119), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT120), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n927), .B1(G898), .B2(new_n378), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n985), .B(new_n986), .ZN(G69));
  INV_X1    g801(.A(new_n823), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT121), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n519), .B1(new_n581), .B2(new_n595), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n701), .A2(new_n755), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n851), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n989), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n722), .A2(KEYINPUT121), .A3(new_n851), .A4(new_n991), .ZN(new_n994));
  AOI22_X1  g808(.A1(new_n909), .A2(new_n988), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n750), .A2(new_n830), .A3(new_n703), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(KEYINPUT62), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT62), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n750), .A2(new_n830), .A3(new_n703), .A4(new_n998), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n820), .A2(new_n995), .A3(new_n997), .A4(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(new_n378), .ZN(new_n1001));
  AND2_X1   g815(.A1(new_n533), .A2(new_n544), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(new_n226), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  OR2_X1    g818(.A1(new_n378), .A2(G900), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(KEYINPUT123), .Z(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n750), .A2(new_n830), .ZN(new_n1008));
  INV_X1    g822(.A(new_n783), .ZN(new_n1009));
  NOR3_X1   g823(.A1(new_n1008), .A2(new_n828), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n621), .A2(new_n693), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n753), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n808), .A2(new_n817), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT124), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n808), .A2(new_n817), .A3(new_n1012), .A4(KEYINPUT124), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n780), .A2(new_n1010), .A3(new_n1017), .A4(new_n820), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1007), .B1(new_n1018), .B2(new_n378), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1004), .B1(new_n1019), .B2(new_n1003), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n378), .B1(G227), .B2(G900), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g836(.A(KEYINPUT125), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1021), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1024), .B1(new_n1019), .B2(new_n1003), .ZN(new_n1025));
  INV_X1    g839(.A(new_n1025), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1004), .A2(KEYINPUT122), .ZN(new_n1027));
  INV_X1    g841(.A(KEYINPUT122), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1001), .A2(new_n1028), .A3(new_n1003), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n1023), .B1(new_n1026), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1028), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1032));
  INV_X1    g846(.A(new_n1003), .ZN(new_n1033));
  AOI211_X1 g847(.A(KEYINPUT122), .B(new_n1033), .C1(new_n1000), .C2(new_n378), .ZN(new_n1034));
  NOR2_X1   g848(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  NOR3_X1   g849(.A1(new_n1035), .A2(new_n1025), .A3(KEYINPUT125), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1022), .B1(new_n1031), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g851(.A(KEYINPUT126), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  OAI211_X1 g853(.A(KEYINPUT126), .B(new_n1022), .C1(new_n1031), .C2(new_n1036), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1039), .A2(new_n1040), .ZN(G72));
  NAND2_X1  g855(.A1(G472), .A2(G902), .ZN(new_n1042));
  XOR2_X1   g856(.A(new_n1042), .B(KEYINPUT63), .Z(new_n1043));
  OAI21_X1  g857(.A(new_n1043), .B1(new_n1000), .B2(new_n980), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n923), .B1(new_n1044), .B2(new_n696), .ZN(new_n1045));
  OAI21_X1  g859(.A(new_n1043), .B1(new_n1018), .B2(new_n980), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n545), .A2(new_n583), .ZN(new_n1047));
  NOR2_X1   g861(.A1(new_n1047), .A2(new_n564), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n1045), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g864(.A(new_n1048), .ZN(new_n1051));
  INV_X1    g865(.A(new_n696), .ZN(new_n1052));
  NAND4_X1  g866(.A1(new_n965), .A2(new_n1051), .A3(new_n1052), .A4(new_n1043), .ZN(new_n1053));
  OR2_X1    g867(.A1(new_n1053), .A2(KEYINPUT127), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n1053), .A2(KEYINPUT127), .ZN(new_n1055));
  AOI21_X1  g869(.A(new_n1050), .B1(new_n1054), .B2(new_n1055), .ZN(G57));
endmodule


