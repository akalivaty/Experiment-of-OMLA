//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 1 0 1 0 1 1 1 1 0 0 0 0 0 0 1 1 1 0 1 1 0 1 1 1 1 0 1 1 1 0 1 1 1 1 1 0 1 1 0 0 0 0 1 0 1 1 0 0 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1335,
    new_n1336;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  XOR2_X1   g0013(.A(KEYINPUT67), .B(G238), .Z(new_n214));
  AND2_X1   g0014(.A1(KEYINPUT66), .A2(G68), .ZN(new_n215));
  NOR2_X1   g0015(.A1(KEYINPUT66), .A2(G68), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G107), .A2(G264), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n210), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G20), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n201), .B(KEYINPUT65), .Z(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n213), .B1(KEYINPUT1), .B2(new_n224), .C1(new_n227), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XOR2_X1   g0040(.A(G50), .B(G58), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  AND2_X1   g0046(.A1(KEYINPUT3), .A2(G33), .ZN(new_n247));
  NOR2_X1   g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g0049(.A(KEYINPUT7), .B1(new_n249), .B2(new_n208), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT7), .ZN(new_n251));
  NOR4_X1   g0051(.A1(new_n247), .A2(new_n248), .A3(new_n251), .A4(G20), .ZN(new_n252));
  OAI21_X1  g0052(.A(G68), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT80), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT80), .ZN(new_n255));
  OAI211_X1 g0055(.A(new_n255), .B(G68), .C1(new_n250), .C2(new_n252), .ZN(new_n256));
  INV_X1    g0056(.A(new_n201), .ZN(new_n257));
  INV_X1    g0057(.A(G58), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n257), .B1(new_n217), .B2(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n259), .A2(G20), .B1(G159), .B2(new_n260), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n254), .A2(KEYINPUT16), .A3(new_n256), .A4(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT81), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AND2_X1   g0064(.A1(new_n256), .A2(new_n261), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n265), .A2(KEYINPUT81), .A3(KEYINPUT16), .A4(new_n254), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT83), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT16), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT82), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT66), .B(G68), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n270), .B(new_n271), .C1(new_n250), .C2(new_n252), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n261), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT3), .B(G33), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n251), .B1(new_n274), .B2(G20), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n249), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n270), .B1(new_n277), .B2(new_n271), .ZN(new_n278));
  OAI211_X1 g0078(.A(new_n268), .B(new_n269), .C1(new_n273), .C2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  AND2_X1   g0080(.A1(new_n280), .A2(new_n225), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n269), .B1(new_n273), .B2(new_n278), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n281), .B1(new_n282), .B2(KEYINPUT83), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n267), .A2(new_n279), .A3(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G33), .ZN(new_n285));
  INV_X1    g0085(.A(G41), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n226), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT85), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(new_n291), .A3(G232), .ZN(new_n292));
  INV_X1    g0092(.A(G232), .ZN(new_n293));
  OAI21_X1  g0093(.A(KEYINPUT85), .B1(new_n289), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G274), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n292), .B(new_n294), .C1(new_n295), .C2(new_n288), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n274), .A2(G1698), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  AOI22_X1  g0098(.A1(new_n298), .A2(G226), .B1(G33), .B2(G87), .ZN(new_n299));
  INV_X1    g0099(.A(G1698), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n274), .A2(G223), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n287), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n296), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G190), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n305), .B1(G200), .B2(new_n303), .ZN(new_n306));
  XNOR2_X1  g0106(.A(KEYINPUT8), .B(G58), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT69), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OR3_X1    g0109(.A1(new_n308), .A2(new_n258), .A3(KEYINPUT8), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n207), .A2(G20), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n280), .A2(new_n225), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AND3_X1   g0117(.A1(new_n312), .A2(new_n313), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n318), .B1(new_n315), .B2(new_n311), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n284), .A2(new_n306), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT17), .ZN(new_n321));
  XNOR2_X1  g0121(.A(new_n320), .B(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n284), .A2(new_n319), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT84), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT84), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n284), .A2(new_n325), .A3(new_n319), .ZN(new_n326));
  INV_X1    g0126(.A(G179), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n303), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n328), .B1(G169), .B2(new_n303), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n324), .A2(new_n326), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT18), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n324), .A2(KEYINPUT18), .A3(new_n326), .A4(new_n330), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n322), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n317), .A2(G50), .A3(new_n313), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n336), .B1(G50), .B2(new_n314), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n260), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n208), .A2(G33), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n338), .B1(new_n311), .B2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n337), .B1(new_n340), .B2(new_n316), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT9), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n341), .B(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n288), .A2(new_n295), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n344), .B1(new_n290), .B2(G226), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n274), .A2(G222), .A3(new_n300), .ZN(new_n346));
  INV_X1    g0146(.A(G77), .ZN(new_n347));
  INV_X1    g0147(.A(G223), .ZN(new_n348));
  OAI221_X1 g0148(.A(new_n346), .B1(new_n347), .B2(new_n274), .C1(new_n297), .C2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT68), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n225), .B1(G33), .B2(G41), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n349), .B2(new_n350), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n345), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G200), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n343), .B(new_n355), .C1(new_n304), .C2(new_n354), .ZN(new_n356));
  XNOR2_X1  g0156(.A(new_n356), .B(KEYINPUT10), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n354), .A2(new_n327), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n358), .B1(G169), .B2(new_n354), .ZN(new_n359));
  OR2_X1    g0159(.A1(new_n359), .A2(new_n341), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  OAI22_X1  g0162(.A1(new_n271), .A2(new_n208), .B1(new_n347), .B2(new_n339), .ZN(new_n363));
  AND2_X1   g0163(.A1(new_n363), .A2(KEYINPUT77), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n260), .A2(G50), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(new_n363), .B2(KEYINPUT77), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n316), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  OR2_X1    g0167(.A1(new_n367), .A2(KEYINPUT78), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(KEYINPUT78), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT11), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n281), .A2(KEYINPUT75), .A3(new_n314), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT75), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n315), .B2(new_n316), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n373), .A2(new_n375), .A3(new_n313), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT12), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n377), .B1(new_n217), .B2(new_n315), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(G68), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n378), .B1(new_n377), .B2(new_n315), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT79), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT79), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n380), .A2(new_n385), .A3(new_n382), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n368), .A2(KEYINPUT11), .A3(new_n369), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n372), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(G238), .ZN(new_n390));
  OAI22_X1  g0190(.A1(new_n289), .A2(new_n390), .B1(new_n344), .B2(KEYINPUT76), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n391), .B1(KEYINPUT76), .B2(new_n344), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n274), .A2(G226), .A3(new_n300), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n274), .A2(G232), .A3(G1698), .ZN(new_n394));
  NAND2_X1  g0194(.A1(G33), .A2(G97), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n352), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n392), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT13), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT13), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n392), .A2(new_n400), .A3(new_n397), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n399), .A2(G179), .A3(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(G169), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n403), .B1(new_n399), .B2(new_n401), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT14), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n402), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n401), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n400), .B1(new_n392), .B2(new_n397), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n405), .B(G169), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n389), .B1(new_n406), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(G200), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(new_n407), .B2(new_n408), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n399), .A2(new_n304), .A3(new_n401), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n415), .A2(new_n387), .A3(new_n388), .A4(new_n372), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n411), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT72), .ZN(new_n418));
  XNOR2_X1  g0218(.A(new_n307), .B(new_n418), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n419), .A2(new_n260), .B1(G20), .B2(G77), .ZN(new_n420));
  OR2_X1    g0220(.A1(new_n420), .A2(KEYINPUT73), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT74), .ZN(new_n422));
  INV_X1    g0222(.A(G87), .ZN(new_n423));
  AND2_X1   g0223(.A1(new_n423), .A2(KEYINPUT15), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n423), .A2(KEYINPUT15), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n422), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  XNOR2_X1  g0226(.A(KEYINPUT15), .B(G87), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT74), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n429), .A2(new_n339), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n430), .B1(new_n420), .B2(KEYINPUT73), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n281), .B1(new_n421), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n315), .A2(new_n347), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n376), .B2(new_n347), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n274), .A2(G232), .A3(new_n300), .ZN(new_n436));
  AND2_X1   g0236(.A1(KEYINPUT70), .A2(G107), .ZN(new_n437));
  NOR2_X1   g0237(.A1(KEYINPUT70), .A2(G107), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OAI221_X1 g0239(.A(new_n436), .B1(new_n439), .B2(new_n274), .C1(new_n297), .C2(new_n214), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n352), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n344), .B1(new_n290), .B2(G244), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n441), .A2(G190), .A3(new_n442), .ZN(new_n443));
  OR2_X1    g0243(.A1(new_n443), .A2(KEYINPUT71), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n441), .A2(new_n442), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n443), .A2(KEYINPUT71), .B1(new_n445), .B2(G200), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n435), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n445), .A2(new_n327), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n449), .B1(G169), .B2(new_n445), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n435), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n335), .A2(new_n362), .A3(new_n417), .A4(new_n452), .ZN(new_n453));
  OAI211_X1 g0253(.A(G244), .B(G1698), .C1(new_n247), .C2(new_n248), .ZN(new_n454));
  OAI211_X1 g0254(.A(G238), .B(new_n300), .C1(new_n247), .C2(new_n248), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G33), .A2(G116), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT88), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n454), .A2(new_n455), .A3(KEYINPUT88), .A4(new_n456), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n459), .A2(new_n352), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n207), .A2(G45), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G250), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n463), .B1(new_n295), .B2(new_n462), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n287), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n412), .B1(new_n461), .B2(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n314), .B1(new_n426), .B2(new_n428), .ZN(new_n467));
  OR2_X1    g0267(.A1(KEYINPUT70), .A2(G107), .ZN(new_n468));
  INV_X1    g0268(.A(G97), .ZN(new_n469));
  NAND2_X1  g0269(.A1(KEYINPUT70), .A2(G107), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n468), .A2(new_n423), .A3(new_n469), .A4(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT19), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n208), .B1(new_n395), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n274), .A2(new_n208), .A3(G68), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n208), .A2(G33), .A3(G97), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n472), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n474), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n467), .B1(new_n478), .B2(new_n316), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n207), .A2(G33), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n281), .A2(new_n314), .A3(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n481), .A2(new_n423), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(KEYINPUT90), .B1(new_n466), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT90), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n471), .A2(new_n473), .B1(new_n472), .B2(new_n476), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n281), .B1(new_n487), .B2(new_n475), .ZN(new_n488));
  NOR3_X1   g0288(.A1(new_n488), .A2(new_n467), .A3(new_n482), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n460), .A2(new_n352), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n490), .A2(new_n459), .B1(new_n287), .B2(new_n464), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n486), .B(new_n489), .C1(new_n491), .C2(new_n412), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n461), .A2(G190), .A3(new_n465), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT91), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n491), .A2(KEYINPUT91), .A3(G190), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n485), .A2(new_n492), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n479), .B1(new_n429), .B2(new_n481), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT89), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT89), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n479), .B(new_n500), .C1(new_n429), .C2(new_n481), .ZN(new_n501));
  AND2_X1   g0301(.A1(new_n457), .A2(new_n458), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n460), .A2(new_n352), .ZN(new_n503));
  OAI211_X1 g0303(.A(G179), .B(new_n465), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n403), .B1(new_n461), .B2(new_n465), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n499), .B(new_n501), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n497), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(KEYINPUT86), .A2(KEYINPUT6), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(G107), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G97), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n469), .A2(G107), .ZN(new_n513));
  NAND2_X1  g0313(.A1(KEYINPUT86), .A2(KEYINPUT6), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n510), .A2(new_n512), .A3(new_n513), .A4(new_n514), .ZN(new_n515));
  AND2_X1   g0315(.A1(KEYINPUT86), .A2(KEYINPUT6), .ZN(new_n516));
  OAI211_X1 g0316(.A(G97), .B(new_n511), .C1(new_n516), .C2(new_n509), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n518), .A2(G20), .B1(G77), .B2(new_n260), .ZN(new_n519));
  INV_X1    g0319(.A(new_n439), .ZN(new_n520));
  OAI211_X1 g0320(.A(KEYINPUT87), .B(new_n520), .C1(new_n250), .C2(new_n252), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(KEYINPUT87), .B1(new_n277), .B2(new_n520), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n316), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n481), .A2(G97), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(G97), .B2(new_n315), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(G244), .B1(new_n247), .B2(new_n248), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT4), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G283), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n529), .A2(G1698), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n532), .B(G244), .C1(new_n248), .C2(new_n247), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  OAI21_X1  g0334(.A(G250), .B1(new_n247), .B2(new_n248), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n300), .B1(new_n535), .B2(KEYINPUT4), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n352), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  OR2_X1    g0337(.A1(KEYINPUT5), .A2(G41), .ZN(new_n538));
  NAND2_X1  g0338(.A1(KEYINPUT5), .A2(G41), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n462), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n540), .A2(new_n352), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n541), .A2(G257), .B1(G274), .B2(new_n540), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n537), .A2(new_n542), .A3(G179), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n540), .A2(G274), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n538), .A2(new_n539), .ZN(new_n545));
  INV_X1    g0345(.A(new_n462), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n287), .ZN(new_n548));
  INV_X1    g0348(.A(G257), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n544), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n528), .A2(new_n529), .B1(G33), .B2(G283), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n529), .B1(new_n274), .B2(G250), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n551), .B(new_n533), .C1(new_n300), .C2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n550), .B1(new_n553), .B2(new_n352), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n543), .B1(new_n554), .B2(new_n403), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n527), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(G257), .B(G1698), .C1(new_n247), .C2(new_n248), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G33), .A2(G294), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n557), .B(new_n558), .C1(new_n535), .C2(G1698), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n352), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n541), .A2(G264), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n560), .A2(new_n544), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n412), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n560), .A2(new_n304), .A3(new_n544), .A4(new_n561), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(KEYINPUT23), .B1(new_n437), .B2(new_n438), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT23), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n567), .A2(new_n511), .A3(G20), .ZN(new_n568));
  AOI21_X1  g0368(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n566), .B(new_n568), .C1(G20), .C2(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n208), .B(G87), .C1(new_n247), .C2(new_n248), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT22), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT22), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n274), .A2(new_n573), .A3(new_n208), .A4(G87), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n570), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n281), .B1(new_n575), .B2(KEYINPUT24), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n572), .A2(new_n574), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n568), .B1(G20), .B2(new_n569), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n578), .B1(new_n520), .B2(KEYINPUT23), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT24), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n576), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(KEYINPUT25), .B1(new_n315), .B2(new_n511), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT93), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(new_n511), .B2(new_n481), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n315), .A2(KEYINPUT25), .A3(new_n511), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(KEYINPUT93), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n589), .A2(new_n584), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n565), .A2(new_n583), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n316), .B1(new_n580), .B2(new_n581), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n575), .A2(KEYINPUT24), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n591), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n562), .A2(G169), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n560), .A2(G179), .A3(new_n544), .A4(new_n561), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n537), .A2(new_n542), .A3(new_n304), .ZN(new_n600));
  AOI21_X1  g0400(.A(G200), .B1(new_n537), .B2(new_n542), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n524), .B(new_n526), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n556), .A2(new_n592), .A3(new_n599), .A4(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n274), .A2(G264), .A3(G1698), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n274), .A2(G257), .A3(new_n300), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n249), .A2(G303), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n352), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n541), .A2(G270), .B1(G274), .B2(new_n540), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n373), .A2(new_n375), .A3(G116), .A4(new_n480), .ZN(new_n612));
  INV_X1    g0412(.A(G116), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n315), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n531), .B1(new_n469), .B2(G33), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n208), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n208), .A2(new_n613), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(KEYINPUT20), .B1(new_n619), .B2(new_n316), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n617), .B1(new_n615), .B2(new_n208), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT20), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n621), .A2(new_n622), .A3(new_n281), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n612), .B(new_n614), .C1(new_n620), .C2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n611), .A2(new_n624), .A3(G179), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n403), .B1(new_n609), .B2(new_n610), .ZN(new_n626));
  AOI21_X1  g0426(.A(KEYINPUT92), .B1(new_n626), .B2(new_n624), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT21), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n625), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n609), .A2(new_n610), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n630), .A2(G190), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n630), .A2(new_n412), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n624), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AOI211_X1 g0434(.A(KEYINPUT92), .B(KEYINPUT21), .C1(new_n626), .C2(new_n624), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n629), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n508), .A2(new_n604), .A3(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n453), .A2(new_n637), .ZN(G372));
  NAND2_X1  g0438(.A1(new_n416), .A2(new_n451), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n322), .B1(new_n411), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n323), .A2(new_n330), .ZN(new_n641));
  XOR2_X1   g0441(.A(KEYINPUT96), .B(KEYINPUT18), .Z(new_n642));
  XNOR2_X1  g0442(.A(new_n641), .B(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n357), .B1(new_n640), .B2(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n645), .A2(new_n360), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n537), .A2(new_n542), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(G169), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n543), .A2(new_n648), .B1(new_n524), .B2(new_n526), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n497), .A2(new_n507), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(KEYINPUT26), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n465), .B1(new_n502), .B2(new_n503), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(G200), .ZN(new_n653));
  AOI21_X1  g0453(.A(KEYINPUT94), .B1(new_n479), .B2(new_n483), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT94), .ZN(new_n655));
  NOR4_X1   g0455(.A1(new_n488), .A2(new_n655), .A3(new_n467), .A4(new_n482), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n653), .B(new_n493), .C1(new_n654), .C2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT26), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n498), .B1(new_n505), .B2(new_n506), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n649), .A2(new_n657), .A3(new_n658), .A4(new_n659), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n660), .A2(new_n659), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n651), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT95), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n651), .A2(new_n661), .A3(KEYINPUT95), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n556), .A2(new_n592), .A3(new_n602), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n657), .A2(new_n659), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n626), .A2(new_n624), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT92), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(KEYINPUT21), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n627), .A2(new_n628), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(new_n673), .A3(new_n625), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n595), .A2(new_n598), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n667), .B(new_n668), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n666), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n646), .B1(new_n453), .B2(new_n678), .ZN(G369));
  INV_X1    g0479(.A(new_n624), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G213), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(G343), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n680), .A2(new_n687), .ZN(new_n688));
  MUX2_X1   g0488(.A(new_n636), .B(new_n674), .S(new_n688), .Z(new_n689));
  XNOR2_X1  g0489(.A(KEYINPUT97), .B(G330), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n595), .A2(new_n686), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n675), .B1(new_n592), .B2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n599), .A2(new_n686), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(new_n674), .A3(new_n687), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n599), .B2(new_n686), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n698), .A2(new_n701), .ZN(G399));
  INV_X1    g0502(.A(new_n211), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(G41), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n471), .A2(G116), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(G1), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(new_n229), .B2(new_n705), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT28), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n686), .B1(new_n666), .B2(new_n676), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n508), .A2(new_n658), .A3(new_n649), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n668), .A2(new_n649), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(KEYINPUT26), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n711), .A2(new_n676), .A3(new_n713), .A4(new_n659), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n687), .ZN(new_n715));
  MUX2_X1   g0515(.A(new_n710), .B(new_n715), .S(KEYINPUT29), .Z(new_n716));
  INV_X1    g0516(.A(KEYINPUT99), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n637), .A2(KEYINPUT31), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT30), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n560), .A2(new_n561), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n554), .A2(new_n611), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n719), .B1(new_n722), .B2(new_n504), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n647), .A2(new_n630), .A3(new_n720), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n724), .A2(KEYINPUT30), .A3(new_n505), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n611), .A2(G179), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n726), .A2(new_n652), .A3(new_n562), .A4(new_n647), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT31), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n723), .A2(new_n725), .A3(new_n727), .A4(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n686), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT98), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n723), .A2(new_n725), .A3(new_n727), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n687), .A2(new_n728), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n731), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n732), .A2(new_n731), .A3(new_n733), .ZN(new_n736));
  AOI22_X1  g0536(.A1(new_n718), .A2(new_n730), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n717), .B1(new_n737), .B2(new_n690), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n497), .A2(new_n507), .ZN(new_n739));
  INV_X1    g0539(.A(new_n633), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n680), .B1(new_n740), .B2(new_n631), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n672), .A2(new_n741), .A3(new_n673), .A4(new_n625), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n739), .A2(new_n742), .A3(new_n603), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n730), .B1(new_n743), .B2(new_n728), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n735), .A2(new_n736), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n746), .A2(KEYINPUT99), .A3(new_n691), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n738), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n716), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n709), .B1(new_n749), .B2(G1), .ZN(G364));
  AND2_X1   g0550(.A1(new_n208), .A2(G13), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G45), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n705), .A2(G1), .A3(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n703), .A2(new_n274), .ZN(new_n754));
  INV_X1    g0554(.A(new_n229), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G45), .ZN(new_n756));
  INV_X1    g0556(.A(G45), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n242), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n754), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n703), .A2(new_n249), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n760), .A2(G355), .B1(new_n613), .B2(new_n703), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G13), .A2(G33), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(G20), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT100), .Z(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n225), .B1(G20), .B2(new_n403), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n753), .B1(new_n762), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(G20), .A2(G179), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT101), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G200), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n773), .A2(new_n202), .A3(new_n304), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G179), .A2(G200), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n775), .A2(G20), .A3(new_n304), .ZN(new_n776));
  INV_X1    g0576(.A(G159), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT32), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n208), .B1(new_n775), .B2(G190), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G97), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n412), .A2(G179), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n783), .A2(G20), .A3(G190), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G87), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n783), .A2(G20), .A3(new_n304), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n249), .B1(new_n788), .B2(G107), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n779), .A2(new_n782), .A3(new_n786), .A4(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n773), .A2(G190), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n774), .B(new_n790), .C1(G68), .C2(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n772), .B(KEYINPUT102), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(new_n412), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n304), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n794), .A2(G190), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n792), .B1(new_n258), .B2(new_n796), .C1(new_n347), .C2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G294), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n780), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n776), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n788), .A2(G283), .B1(new_n802), .B2(G329), .ZN(new_n803));
  INV_X1    g0603(.A(G303), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n803), .B(new_n249), .C1(new_n804), .C2(new_n784), .ZN(new_n805));
  XNOR2_X1  g0605(.A(KEYINPUT33), .B(G317), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n801), .B(new_n805), .C1(new_n791), .C2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n797), .A2(G311), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n795), .A2(G322), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n773), .A2(new_n304), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(G326), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n807), .A2(new_n808), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n799), .A2(KEYINPUT103), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(new_n768), .ZN(new_n814));
  AOI21_X1  g0614(.A(KEYINPUT103), .B1(new_n799), .B2(new_n812), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n770), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n689), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n816), .B1(new_n817), .B2(new_n767), .ZN(new_n818));
  INV_X1    g0618(.A(new_n753), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n693), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n689), .A2(new_n691), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n818), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(G396));
  NOR3_X1   g0624(.A1(new_n435), .A2(new_n450), .A3(new_n687), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT105), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n451), .B(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n686), .B1(new_n432), .B2(new_n434), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n447), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n825), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n710), .B(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n748), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n753), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n835), .A2(KEYINPUT106), .B1(new_n834), .B2(new_n833), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(KEYINPUT106), .B2(new_n835), .ZN(new_n837));
  INV_X1    g0637(.A(new_n768), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n764), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n819), .B1(G77), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(G283), .ZN(new_n841));
  NOR3_X1   g0641(.A1(new_n773), .A2(G190), .A3(new_n841), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n785), .A2(G107), .B1(new_n802), .B2(G311), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n274), .B1(new_n788), .B2(G87), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n843), .A2(new_n844), .A3(new_n782), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n842), .B(new_n845), .C1(G303), .C2(new_n810), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n846), .B1(new_n798), .B2(new_n613), .C1(new_n800), .C2(new_n796), .ZN(new_n847));
  AOI22_X1  g0647(.A1(G137), .A2(new_n810), .B1(new_n791), .B2(G150), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n798), .B2(new_n777), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(G143), .B2(new_n795), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(KEYINPUT34), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n788), .A2(G68), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n202), .B2(new_n784), .ZN(new_n853));
  XOR2_X1   g0653(.A(new_n853), .B(KEYINPUT104), .Z(new_n854));
  NAND2_X1  g0654(.A1(new_n781), .A2(G58), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n249), .B1(new_n802), .B2(G132), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n847), .B1(new_n851), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n840), .B1(new_n858), .B2(new_n768), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n832), .B2(new_n764), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n837), .A2(new_n860), .ZN(G384));
  NOR2_X1   g0661(.A1(new_n227), .A2(new_n613), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n518), .B2(KEYINPUT35), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(KEYINPUT35), .B2(new_n518), .ZN(new_n864));
  XOR2_X1   g0664(.A(KEYINPUT107), .B(KEYINPUT36), .Z(new_n865));
  XNOR2_X1  g0665(.A(new_n864), .B(new_n865), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n755), .B(G77), .C1(new_n258), .C2(new_n217), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n202), .A2(G68), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n207), .B(G13), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n827), .A2(new_n686), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(new_n710), .B2(new_n832), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n389), .A2(new_n686), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n411), .A2(new_n416), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n873), .B1(new_n411), .B2(new_n416), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n684), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n324), .A2(new_n326), .A3(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT37), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n320), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n331), .A2(new_n879), .A3(new_n882), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n265), .A2(new_n254), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n267), .B(new_n316), .C1(KEYINPUT16), .C2(new_n884), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n885), .A2(new_n319), .B1(new_n329), .B2(new_n684), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n284), .A2(new_n306), .A3(new_n319), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT37), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n883), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n684), .B1(new_n885), .B2(new_n319), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n889), .B1(new_n335), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT38), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI211_X1 g0694(.A(KEYINPUT38), .B(new_n889), .C1(new_n335), .C2(new_n891), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n877), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n644), .A2(new_n684), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n411), .A2(new_n686), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n322), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n284), .A2(new_n325), .A3(new_n319), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n325), .B1(new_n284), .B2(new_n319), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT18), .B1(new_n905), .B2(new_n330), .ZN(new_n906));
  INV_X1    g0706(.A(new_n334), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n902), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n890), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT38), .B1(new_n909), .B2(new_n889), .ZN(new_n910));
  INV_X1    g0710(.A(new_n895), .ZN(new_n911));
  OAI21_X1  g0711(.A(KEYINPUT39), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n641), .A2(new_n320), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n880), .B1(new_n913), .B2(new_n879), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n883), .A2(KEYINPUT108), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT108), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n331), .A2(new_n879), .A3(new_n882), .A4(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n914), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n879), .B1(new_n902), .B2(new_n643), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n893), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT39), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n920), .A2(new_n921), .A3(new_n895), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n901), .B1(new_n912), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n899), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n453), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n716), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n646), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n924), .B(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n914), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n881), .B1(new_n905), .B2(new_n330), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n916), .B1(new_n930), .B2(new_n879), .ZN(new_n931));
  INV_X1    g0731(.A(new_n917), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n919), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n911), .B1(new_n935), .B2(new_n893), .ZN(new_n936));
  INV_X1    g0736(.A(new_n730), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(new_n637), .B2(KEYINPUT31), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n732), .A2(new_n733), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(KEYINPUT109), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT109), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n744), .A2(new_n942), .A3(new_n939), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n876), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n944), .A2(KEYINPUT40), .A3(new_n832), .A4(new_n945), .ZN(new_n946));
  NOR3_X1   g0746(.A1(new_n938), .A2(KEYINPUT109), .A3(new_n940), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n942), .B1(new_n744), .B2(new_n939), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n945), .B(new_n832), .C1(new_n947), .C2(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(new_n894), .B2(new_n895), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n936), .A2(new_n946), .B1(new_n950), .B2(KEYINPUT40), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n925), .A2(new_n944), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n951), .B(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n953), .A2(new_n690), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n928), .A2(new_n954), .B1(new_n207), .B2(new_n751), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n928), .A2(new_n954), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n870), .B1(new_n955), .B2(new_n956), .ZN(G367));
  INV_X1    g0757(.A(new_n754), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n769), .B1(new_n211), .B2(new_n429), .C1(new_n238), .C2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n819), .B1(new_n959), .B2(KEYINPUT112), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(KEYINPUT112), .B2(new_n959), .ZN(new_n961));
  OR3_X1    g0761(.A1(new_n654), .A2(new_n656), .A3(new_n687), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n668), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(new_n659), .B2(new_n963), .ZN(new_n965));
  INV_X1    g0765(.A(G317), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n249), .B1(new_n776), .B2(new_n966), .C1(new_n787), .C2(new_n469), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n784), .A2(new_n613), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT46), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n967), .B(new_n969), .C1(new_n520), .C2(new_n781), .ZN(new_n970));
  AOI22_X1  g0770(.A1(G294), .A2(new_n791), .B1(new_n810), .B2(G311), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n972), .B1(new_n841), .B2(new_n798), .C1(new_n804), .C2(new_n796), .ZN(new_n973));
  NOR3_X1   g0773(.A1(new_n773), .A2(new_n777), .A3(G190), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n785), .A2(G58), .B1(new_n802), .B2(G137), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n249), .B1(new_n788), .B2(G77), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n781), .A2(G68), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  AOI211_X1 g0778(.A(new_n974), .B(new_n978), .C1(G143), .C2(new_n810), .ZN(new_n979));
  INV_X1    g0779(.A(G150), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n979), .B1(new_n798), .B2(new_n202), .C1(new_n980), .C2(new_n796), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n973), .A2(KEYINPUT47), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n768), .ZN(new_n983));
  AOI21_X1  g0783(.A(KEYINPUT47), .B1(new_n973), .B2(new_n981), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n961), .B1(new_n766), .B2(new_n965), .C1(new_n983), .C2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n752), .A2(G1), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n527), .A2(new_n686), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n556), .A2(new_n987), .A3(new_n602), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n649), .A2(new_n686), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n700), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT45), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n700), .A2(new_n990), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT44), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n993), .B(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n992), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(new_n698), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT110), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n674), .A2(new_n687), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n695), .B2(new_n696), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n699), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n998), .B2(new_n1000), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n693), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT111), .Z(new_n1004));
  OR2_X1    g0804(.A1(new_n1002), .A2(new_n693), .ZN(new_n1005));
  AND3_X1   g0805(.A1(new_n749), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n997), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n749), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n704), .B(KEYINPUT41), .Z(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n986), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n699), .A2(new_n990), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT42), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n556), .B1(new_n988), .B2(new_n599), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n687), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1012), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1020), .B(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n698), .A2(new_n990), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1022), .B(new_n1023), .Z(new_n1024));
  OAI21_X1  g0824(.A(new_n985), .B1(new_n1011), .B2(new_n1024), .ZN(G387));
  NOR2_X1   g0825(.A1(new_n1006), .A2(new_n705), .ZN(new_n1026));
  AND2_X1   g0826(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1026), .B1(new_n749), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n986), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n419), .A2(new_n202), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT50), .Z(new_n1031));
  AOI21_X1  g0831(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1031), .A2(new_n706), .A3(new_n1032), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1033), .B(new_n754), .C1(new_n235), .C2(new_n757), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n760), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1034), .B1(G107), .B2(new_n211), .C1(new_n706), .C2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n753), .B1(new_n1036), .B2(new_n769), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n784), .A2(new_n347), .B1(new_n776), .B2(new_n980), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n249), .B(new_n1038), .C1(G97), .C2(new_n788), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n810), .A2(G159), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n791), .A2(new_n312), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n426), .A2(new_n428), .A3(new_n781), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .A4(new_n1042), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n796), .A2(new_n202), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1043), .B(new_n1044), .C1(G68), .C2(new_n797), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G311), .A2(new_n791), .B1(new_n810), .B2(G322), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n798), .B2(new_n804), .C1(new_n966), .C2(new_n796), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT48), .ZN(new_n1048));
  AND2_X1   g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n784), .A2(new_n800), .B1(new_n780), .B2(new_n841), .ZN(new_n1051));
  NOR3_X1   g0851(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n1052), .A2(KEYINPUT49), .ZN(new_n1053));
  INV_X1    g0853(.A(G326), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n249), .B1(new_n776), .B2(new_n1054), .C1(new_n787), .C2(new_n613), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n1052), .B2(KEYINPUT49), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1045), .B1(new_n1053), .B2(new_n1056), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1037), .B1(new_n697), .B2(new_n766), .C1(new_n1057), .C2(new_n838), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1028), .A2(new_n1029), .A3(new_n1058), .ZN(G393));
  OR2_X1    g0859(.A1(new_n997), .A2(new_n1006), .ZN(new_n1060));
  AND3_X1   g0860(.A1(new_n1060), .A2(new_n704), .A3(new_n1007), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(KEYINPUT114), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n990), .A2(new_n767), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n769), .B1(new_n469), .B2(new_n211), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n958), .A2(new_n245), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n819), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n795), .A2(G159), .B1(G150), .B2(new_n810), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT51), .Z(new_n1068));
  AOI22_X1  g0868(.A1(new_n785), .A2(new_n271), .B1(new_n802), .B2(G143), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1069), .A2(KEYINPUT113), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n780), .A2(new_n347), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n249), .B(new_n1071), .C1(G87), .C2(new_n788), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n791), .A2(G50), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1069), .A2(KEYINPUT113), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1070), .A2(new_n1072), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(new_n419), .B2(new_n797), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1068), .A2(new_n1076), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n795), .A2(G311), .B1(G317), .B2(new_n810), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT52), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n785), .A2(G283), .B1(new_n802), .B2(G322), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n274), .B1(new_n788), .B2(G107), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n781), .A2(G116), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(G303), .B2(new_n791), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n798), .B2(new_n800), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1077), .B1(new_n1079), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1066), .B1(new_n1086), .B2(new_n768), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n997), .A2(new_n986), .B1(new_n1063), .B2(new_n1087), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n1062), .A2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1061), .A2(KEYINPUT114), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1089), .A2(new_n1091), .ZN(G390));
  AOI21_X1  g0892(.A(new_n831), .B1(new_n941), .B2(new_n943), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1093), .A2(G330), .A3(new_n945), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n901), .B1(new_n872), .B2(new_n876), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n912), .A2(new_n922), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n920), .A2(new_n895), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n714), .A2(new_n687), .A3(new_n827), .A4(new_n830), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n871), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1097), .B(new_n901), .C1(new_n876), .C2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1094), .B1(new_n1096), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  NOR3_X1   g0904(.A1(new_n737), .A2(new_n717), .A3(new_n690), .ZN(new_n1105));
  AOI21_X1  g0905(.A(KEYINPUT99), .B1(new_n746), .B2(new_n691), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n832), .B(new_n945), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1096), .A2(new_n1102), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1104), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT116), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n831), .B1(new_n738), .B2(new_n747), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1094), .B1(new_n1111), .B2(new_n945), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n872), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1100), .B1(new_n1111), .B2(new_n945), .ZN(new_n1115));
  OAI211_X1 g0915(.A(G330), .B(new_n832), .C1(new_n947), .C2(new_n948), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n876), .ZN(new_n1117));
  AOI21_X1  g0917(.A(KEYINPUT115), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  AND4_X1   g0918(.A1(KEYINPUT115), .A2(new_n1107), .A3(new_n1117), .A4(new_n1101), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1114), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n925), .A2(G330), .A3(new_n944), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n926), .A2(new_n646), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1110), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n705), .B1(new_n1109), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(KEYINPUT116), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n1096), .A2(new_n1102), .A3(new_n1107), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1128), .A2(new_n1103), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1125), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n912), .A2(new_n922), .A3(new_n763), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n819), .B1(new_n312), .B2(new_n839), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n802), .A2(G294), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n786), .A2(new_n852), .A3(new_n249), .A4(new_n1134), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n1071), .B(new_n1135), .C1(G283), .C2(new_n810), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n791), .A2(new_n520), .ZN(new_n1137));
  AND2_X1   g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n1138), .B1(new_n469), .B2(new_n798), .C1(new_n613), .C2(new_n796), .ZN(new_n1139));
  XOR2_X1   g0939(.A(KEYINPUT54), .B(G143), .Z(new_n1140));
  NAND2_X1  g0940(.A1(new_n797), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n795), .A2(G132), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n274), .B1(new_n787), .B2(new_n202), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(KEYINPUT117), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n784), .A2(new_n980), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT53), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n781), .A2(G159), .B1(new_n802), .B2(G125), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n1143), .A2(KEYINPUT117), .ZN(new_n1148));
  AND4_X1   g0948(.A1(new_n1144), .A2(new_n1146), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(G128), .A2(new_n810), .B1(new_n791), .B2(G137), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1141), .A2(new_n1142), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1139), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1133), .B1(new_n1152), .B2(new_n768), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1132), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n986), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1154), .B1(new_n1109), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1131), .A2(new_n1157), .ZN(G378));
  OAI21_X1  g0958(.A(new_n819), .B1(G50), .B2(new_n839), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n791), .A2(G132), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n785), .A2(new_n1140), .B1(new_n781), .B2(G150), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(G125), .B2(new_n810), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n797), .A2(G137), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n795), .A2(G128), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  OR2_X1    g0966(.A1(new_n1166), .A2(KEYINPUT59), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(KEYINPUT59), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n285), .B(new_n286), .C1(new_n787), .C2(new_n777), .ZN(new_n1169));
  XOR2_X1   g0969(.A(KEYINPUT118), .B(G124), .Z(new_n1170));
  AOI21_X1  g0970(.A(new_n1169), .B1(new_n802), .B2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1167), .A2(new_n1168), .A3(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(new_n249), .B2(new_n286), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n810), .A2(G116), .ZN(new_n1175));
  AOI211_X1 g0975(.A(G41), .B(new_n274), .C1(new_n785), .C2(G77), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n788), .A2(G58), .B1(new_n802), .B2(G283), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1175), .A2(new_n977), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G97), .B2(new_n791), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1179), .B1(new_n511), .B2(new_n796), .C1(new_n429), .C2(new_n798), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT58), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1174), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1172), .B(new_n1182), .C1(new_n1181), .C2(new_n1180), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1159), .B1(new_n1183), .B2(new_n768), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n341), .A2(new_n684), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n361), .B(new_n1185), .ZN(new_n1186));
  XOR2_X1   g0986(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1186), .B(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1184), .B1(new_n1190), .B2(new_n764), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT119), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT120), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n899), .B2(new_n923), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n949), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n910), .B2(new_n911), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT40), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n946), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n1197), .A2(new_n1198), .B1(new_n1097), .B2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1190), .B1(new_n1200), .B2(G330), .ZN(new_n1201));
  AOI21_X1  g1001(.A(KEYINPUT40), .B1(new_n896), .B2(new_n1196), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n946), .B1(new_n920), .B2(new_n895), .ZN(new_n1203));
  INV_X1    g1003(.A(G330), .ZN(new_n1204));
  NOR4_X1   g1004(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .A4(new_n1189), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1195), .B1(new_n1201), .B2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1189), .B1(new_n951), .B2(new_n1204), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n920), .A2(new_n921), .A3(new_n895), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n921), .B1(new_n894), .B2(new_n895), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n900), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n877), .A2(new_n896), .B1(new_n644), .B2(new_n684), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1203), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1213), .A2(new_n1214), .A3(G330), .A4(new_n1190), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1207), .A2(new_n1212), .A3(new_n1194), .A4(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1206), .A2(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1193), .B1(new_n1217), .B2(new_n1155), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n924), .B1(new_n1201), .B2(new_n1205), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1207), .A2(new_n1212), .A3(new_n1215), .ZN(new_n1220));
  AND3_X1   g1020(.A1(new_n1219), .A2(KEYINPUT57), .A3(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1120), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1123), .B1(new_n1109), .B2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n705), .B1(new_n1221), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT57), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1122), .B1(new_n1129), .B2(new_n1120), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1225), .B1(new_n1226), .B2(new_n1217), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1218), .B1(new_n1224), .B2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(G375));
  OAI211_X1 g1029(.A(new_n1122), .B(new_n1114), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1126), .A2(new_n1010), .A3(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n876), .A2(new_n763), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n819), .B1(G68), .B2(new_n839), .ZN(new_n1233));
  NOR3_X1   g1033(.A1(new_n773), .A2(new_n613), .A3(G190), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n785), .A2(G97), .B1(new_n802), .B2(G303), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n274), .B1(new_n788), .B2(G77), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1235), .A2(new_n1236), .A3(new_n1042), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n1234), .B(new_n1237), .C1(G294), .C2(new_n810), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1238), .B1(new_n798), .B2(new_n439), .C1(new_n841), .C2(new_n796), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n798), .A2(new_n980), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n795), .A2(G137), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n810), .A2(G132), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n785), .A2(G159), .B1(new_n802), .B2(G128), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n249), .B1(new_n788), .B2(G58), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1243), .B(new_n1244), .C1(new_n202), .C2(new_n780), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(new_n791), .B2(new_n1140), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1241), .A2(new_n1242), .A3(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1239), .B1(new_n1240), .B2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1233), .B1(new_n1248), .B2(new_n768), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1120), .A2(new_n986), .B1(new_n1232), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1231), .A2(new_n1250), .ZN(G381));
  INV_X1    g1051(.A(G387), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1089), .A2(new_n1252), .A3(new_n1091), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1254));
  AND2_X1   g1054(.A1(new_n1254), .A2(KEYINPUT121), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1254), .A2(KEYINPUT121), .ZN(new_n1256));
  NOR4_X1   g1056(.A1(new_n1253), .A2(new_n1255), .A3(new_n1256), .A4(G381), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1257), .B(KEYINPUT122), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(G375), .A2(G378), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  OR2_X1    g1060(.A1(new_n1258), .A2(new_n1260), .ZN(G407));
  OAI211_X1 g1061(.A(G407), .B(G213), .C1(G343), .C2(new_n1260), .ZN(G409));
  INV_X1    g1062(.A(KEYINPUT123), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1219), .A2(new_n986), .A3(new_n1220), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n1191), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1226), .A2(new_n1217), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1265), .B1(new_n1266), .B2(new_n1010), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1263), .B1(new_n1267), .B2(G378), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1156), .B1(new_n1125), .B2(new_n1130), .ZN(new_n1269));
  NOR3_X1   g1069(.A1(new_n1226), .A2(new_n1217), .A3(new_n1009), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1269), .B(KEYINPUT123), .C1(new_n1270), .C2(new_n1265), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1218), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1217), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT57), .B1(new_n1273), .B2(new_n1223), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1219), .A2(KEYINPUT57), .A3(new_n1220), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n704), .B1(new_n1226), .B2(new_n1275), .ZN(new_n1276));
  OAI211_X1 g1076(.A(G378), .B(new_n1272), .C1(new_n1274), .C2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1268), .A2(new_n1271), .A3(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT62), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n685), .A2(G213), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1230), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1281), .B1(new_n1126), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT60), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n704), .B1(new_n1230), .B2(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1250), .B1(new_n1284), .B2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(G384), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  OAI211_X1 g1089(.A(G384), .B(new_n1250), .C1(new_n1284), .C2(new_n1286), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1278), .A2(new_n1279), .A3(new_n1280), .A4(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT61), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1280), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1269), .B1(new_n1270), .B2(new_n1265), .ZN(new_n1295));
  AOI22_X1  g1095(.A1(G378), .A2(new_n1228), .B1(new_n1295), .B2(new_n1263), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1294), .B1(new_n1296), .B2(new_n1271), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT125), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1289), .A2(new_n1298), .A3(new_n1290), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1298), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1294), .A2(G2897), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1299), .B1(new_n1300), .B2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1291), .A2(new_n1298), .A3(new_n1301), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  OAI211_X1 g1105(.A(new_n1292), .B(new_n1293), .C1(new_n1297), .C2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1278), .A2(new_n1280), .A3(new_n1291), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1307), .A2(KEYINPUT62), .ZN(new_n1308));
  OAI21_X1  g1108(.A(KEYINPUT127), .B1(new_n1306), .B2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1062), .A2(new_n1088), .ZN(new_n1310));
  OAI21_X1  g1110(.A(G387), .B1(new_n1310), .B2(new_n1090), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1253), .A2(new_n1311), .ZN(new_n1312));
  XNOR2_X1  g1112(.A(G393), .B(new_n823), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1313), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1253), .A2(new_n1315), .A3(new_n1311), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1314), .A2(new_n1316), .ZN(new_n1317));
  AND2_X1   g1117(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1278), .A2(new_n1280), .ZN(new_n1319));
  AOI21_X1  g1119(.A(KEYINPUT61), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT127), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1307), .A2(KEYINPUT62), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1320), .A2(new_n1321), .A3(new_n1322), .A4(new_n1292), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1309), .A2(new_n1317), .A3(new_n1323), .ZN(new_n1324));
  OAI21_X1  g1124(.A(KEYINPUT126), .B1(new_n1317), .B2(KEYINPUT61), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT126), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1314), .A2(new_n1316), .A3(new_n1326), .A4(new_n1293), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1325), .A2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1307), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(KEYINPUT63), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT63), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1331), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1332));
  OAI211_X1 g1132(.A(new_n1328), .B(new_n1330), .C1(new_n1329), .C2(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1324), .A2(new_n1333), .ZN(G405));
  XNOR2_X1  g1134(.A(new_n1317), .B(new_n1291), .ZN(new_n1335));
  XNOR2_X1  g1135(.A(new_n1228), .B(G378), .ZN(new_n1336));
  XNOR2_X1  g1136(.A(new_n1335), .B(new_n1336), .ZN(G402));
endmodule


