//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 0 0 1 0 0 1 0 0 1 0 0 1 0 0 0 0 1 0 1 0 0 1 1 1 0 1 1 0 1 1 1 0 1 0 0 0 0 0 0 1 1 1 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n631,
    new_n632, new_n633, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n706, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n795, new_n796, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926;
  NAND2_X1  g000(.A1(G29gat), .A2(G36gat), .ZN(new_n202));
  OAI21_X1  g001(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  NOR3_X1   g003(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(G43gat), .B(G50gat), .ZN(new_n206));
  OAI221_X1 g005(.A(new_n202), .B1(new_n204), .B2(new_n205), .C1(new_n206), .C2(KEYINPUT15), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(KEYINPUT15), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n209), .A2(KEYINPUT17), .ZN(new_n210));
  XNOR2_X1  g009(.A(G15gat), .B(G22gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT16), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n211), .B1(new_n212), .B2(G1gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(KEYINPUT90), .A2(G8gat), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n213), .B(new_n214), .C1(G1gat), .C2(new_n211), .ZN(new_n215));
  NOR2_X1   g014(.A1(KEYINPUT90), .A2(G8gat), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n215), .B(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n209), .A2(KEYINPUT17), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n210), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G229gat), .A2(G233gat), .ZN(new_n220));
  INV_X1    g019(.A(new_n217), .ZN(new_n221));
  INV_X1    g020(.A(new_n209), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n219), .A2(new_n220), .A3(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT91), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT18), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT92), .B1(new_n217), .B2(new_n209), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n223), .A2(new_n228), .ZN(new_n229));
  XOR2_X1   g028(.A(new_n220), .B(KEYINPUT13), .Z(new_n230));
  NAND3_X1  g029(.A1(new_n221), .A2(KEYINPUT92), .A3(new_n222), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n225), .A2(new_n226), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n219), .A2(new_n220), .A3(new_n223), .A4(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n227), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT11), .B(G169gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(G197gat), .ZN(new_n237));
  XOR2_X1   g036(.A(G113gat), .B(G141gat), .Z(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n239), .B(KEYINPUT12), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n235), .A2(new_n241), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n227), .A2(new_n240), .A3(new_n232), .A4(new_n234), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G197gat), .B(G204gat), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT22), .ZN(new_n247));
  INV_X1    g046(.A(G211gat), .ZN(new_n248));
  INV_X1    g047(.A(G218gat), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n246), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G211gat), .B(G218gat), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n251), .B(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n255));
  INV_X1    g054(.A(G169gat), .ZN(new_n256));
  INV_X1    g055(.A(G176gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT23), .ZN(new_n259));
  AND2_X1   g058(.A1(new_n259), .A2(KEYINPUT66), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(KEYINPUT66), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n258), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n256), .A2(new_n257), .A3(KEYINPUT23), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n264));
  NAND2_X1  g063(.A1(G169gat), .A2(G176gat), .ZN(new_n265));
  AND3_X1   g064(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n264), .B1(new_n263), .B2(new_n265), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n262), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NOR2_X1   g067(.A1(G183gat), .A2(G190gat), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n269), .B1(new_n270), .B2(KEYINPUT68), .ZN(new_n271));
  NAND2_X1  g070(.A1(G183gat), .A2(G190gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT68), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT24), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT25), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n255), .B1(new_n268), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT65), .B(G176gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n278), .A2(KEYINPUT23), .A3(new_n256), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n269), .A2(KEYINPUT64), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT24), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n272), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT64), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n283), .B1(G183gat), .B2(G190gat), .ZN(new_n284));
  NAND3_X1  g083(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n280), .A2(new_n282), .A3(new_n284), .A4(new_n285), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n279), .A2(new_n286), .A3(new_n262), .A4(new_n265), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT25), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n263), .A2(new_n265), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT67), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n288), .B1(new_n271), .B2(new_n274), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n293), .A2(new_n294), .A3(KEYINPUT69), .A4(new_n262), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n277), .A2(new_n289), .A3(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT27), .B(G183gat), .ZN(new_n297));
  INV_X1    g096(.A(G190gat), .ZN(new_n298));
  AOI21_X1  g097(.A(KEYINPUT70), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT71), .B(KEYINPUT28), .ZN(new_n300));
  OR2_X1    g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n300), .ZN(new_n302));
  OR2_X1    g101(.A1(new_n258), .A2(KEYINPUT26), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n258), .A2(KEYINPUT26), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n303), .A2(new_n304), .A3(new_n265), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n301), .A2(new_n272), .A3(new_n302), .A4(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT29), .B1(new_n296), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(G226gat), .A2(G233gat), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(KEYINPUT76), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n308), .B1(new_n296), .B2(new_n306), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n296), .A2(new_n306), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT29), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n311), .B1(new_n314), .B2(new_n308), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n254), .B(new_n310), .C1(new_n315), .C2(KEYINPUT76), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n254), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n251), .A2(new_n253), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n252), .B1(new_n250), .B2(new_n246), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT75), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n307), .A2(new_n309), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n323), .B1(new_n324), .B2(new_n311), .ZN(new_n325));
  XOR2_X1   g124(.A(G8gat), .B(G36gat), .Z(new_n326));
  XNOR2_X1  g125(.A(new_n326), .B(G64gat), .ZN(new_n327));
  INV_X1    g126(.A(G92gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n327), .B(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n316), .A2(new_n325), .A3(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT77), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT30), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n316), .A2(KEYINPUT77), .A3(new_n325), .A4(new_n330), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(G155gat), .ZN(new_n337));
  INV_X1    g136(.A(G162gat), .ZN(new_n338));
  OAI21_X1  g137(.A(KEYINPUT2), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT78), .ZN(new_n340));
  INV_X1    g139(.A(G141gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n341), .A2(G148gat), .ZN(new_n342));
  INV_X1    g141(.A(G148gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n343), .A2(G141gat), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n339), .B(new_n340), .C1(new_n342), .C2(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G155gat), .B(G162gat), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  XOR2_X1   g147(.A(G141gat), .B(G148gat), .Z(new_n349));
  NAND4_X1  g148(.A1(new_n349), .A2(new_n340), .A3(new_n346), .A4(new_n339), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G127gat), .B(G134gat), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(G120gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(G113gat), .ZN(new_n356));
  INV_X1    g155(.A(G113gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(G120gat), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT1), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n354), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT72), .ZN(new_n361));
  INV_X1    g160(.A(G127gat), .ZN(new_n362));
  NOR3_X1   g161(.A1(new_n361), .A2(new_n362), .A3(G134gat), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n363), .B1(new_n361), .B2(new_n353), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n360), .B1(new_n364), .B2(new_n359), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n352), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n360), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n353), .A2(new_n361), .ZN(new_n368));
  INV_X1    g167(.A(new_n363), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n359), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(new_n351), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n366), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(G225gat), .A2(G233gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n374), .B(KEYINPUT79), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT80), .B(KEYINPUT5), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT4), .B1(new_n371), .B2(new_n351), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT4), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n365), .A2(new_n379), .A3(new_n348), .A4(new_n350), .ZN(new_n380));
  AND2_X1   g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n351), .A2(KEYINPUT3), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT3), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n348), .A2(new_n383), .A3(new_n350), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n382), .A2(new_n371), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n375), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n376), .B(new_n377), .C1(new_n381), .C2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n380), .A2(KEYINPUT81), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT81), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n352), .A2(new_n390), .A3(new_n379), .A4(new_n365), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n389), .A2(new_n391), .A3(new_n378), .ZN(new_n392));
  INV_X1    g191(.A(new_n377), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n392), .A2(new_n386), .A3(new_n393), .A4(new_n385), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n388), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(KEYINPUT0), .B(G57gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n396), .B(G85gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(G1gat), .B(G29gat), .ZN(new_n398));
  XOR2_X1   g197(.A(new_n397), .B(new_n398), .Z(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT82), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n388), .A2(new_n394), .A3(new_n399), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT6), .ZN(new_n404));
  AND2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n399), .B1(new_n388), .B2(new_n394), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT82), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n402), .A2(new_n405), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n406), .A2(KEYINPUT6), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n330), .B1(new_n316), .B2(new_n325), .ZN(new_n412));
  AND3_X1   g211(.A1(new_n316), .A2(new_n325), .A3(new_n330), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n412), .B1(new_n413), .B2(KEYINPUT30), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n336), .A2(new_n411), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(G227gat), .ZN(new_n416));
  INV_X1    g215(.A(G233gat), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n296), .A2(new_n365), .A3(new_n306), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n365), .B1(new_n296), .B2(new_n306), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n418), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT33), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n422), .B1(KEYINPUT32), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G15gat), .B(G43gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(G71gat), .ZN(new_n426));
  INV_X1    g225(.A(G99gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT73), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT32), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n312), .A2(new_n371), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n419), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n431), .B1(new_n433), .B2(new_n418), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n428), .A2(KEYINPUT33), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n430), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AND4_X1   g235(.A1(new_n430), .A2(new_n422), .A3(KEYINPUT32), .A4(new_n435), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n429), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  XNOR2_X1  g237(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n420), .A2(new_n421), .ZN(new_n441));
  INV_X1    g240(.A(new_n418), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NOR3_X1   g242(.A1(new_n433), .A2(new_n418), .A3(new_n439), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n438), .A2(new_n446), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n445), .B(new_n429), .C1(new_n436), .C2(new_n437), .ZN(new_n448));
  XNOR2_X1  g247(.A(G78gat), .B(G106gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n449), .B(KEYINPUT31), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n450), .B(G50gat), .ZN(new_n451));
  XOR2_X1   g250(.A(new_n451), .B(KEYINPUT83), .Z(new_n452));
  AOI22_X1  g251(.A1(new_n318), .A2(new_n322), .B1(new_n313), .B2(new_n384), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n313), .B1(new_n319), .B2(new_n320), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n352), .B1(new_n383), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(G228gat), .A2(G233gat), .ZN(new_n456));
  NOR3_X1   g255(.A1(new_n453), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n455), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n384), .A2(new_n313), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n321), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT84), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT84), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n459), .A2(new_n462), .A3(new_n321), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n458), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n457), .B1(new_n456), .B2(new_n464), .ZN(new_n465));
  XOR2_X1   g264(.A(KEYINPUT85), .B(G22gat), .Z(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  AOI211_X1 g267(.A(new_n466), .B(new_n457), .C1(new_n456), .C2(new_n464), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n452), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n465), .A2(new_n467), .ZN(new_n471));
  INV_X1    g270(.A(G22gat), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n471), .B(new_n451), .C1(new_n472), .C2(new_n465), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n447), .A2(new_n448), .A3(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT35), .B1(new_n415), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT89), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT89), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n478), .B(KEYINPUT35), .C1(new_n415), .C2(new_n475), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n336), .A2(new_n414), .ZN(new_n481));
  INV_X1    g280(.A(new_n410), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n482), .B1(new_n401), .B2(new_n405), .ZN(new_n483));
  OR4_X1    g282(.A1(KEYINPUT35), .A2(new_n481), .A3(new_n475), .A4(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n333), .A2(new_n335), .ZN(new_n486));
  XNOR2_X1  g285(.A(KEYINPUT86), .B(KEYINPUT38), .ZN(new_n487));
  XNOR2_X1  g286(.A(KEYINPUT87), .B(KEYINPUT37), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n316), .A2(new_n325), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n329), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT37), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n491), .B1(new_n316), .B2(new_n325), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n487), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT76), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n494), .B1(new_n324), .B2(new_n311), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n254), .B1(new_n495), .B2(new_n310), .ZN(new_n496));
  NOR3_X1   g295(.A1(new_n324), .A2(new_n311), .A3(new_n323), .ZN(new_n497));
  OAI21_X1  g296(.A(KEYINPUT37), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n487), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n498), .A2(new_n329), .A3(new_n499), .A4(new_n489), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n486), .A2(new_n493), .A3(new_n483), .A4(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(new_n474), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n386), .B1(new_n392), .B2(new_n385), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT39), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n373), .A2(new_n375), .ZN(new_n505));
  OR3_X1    g304(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n400), .B1(new_n503), .B2(new_n504), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT40), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n508), .A2(new_n509), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(new_n401), .ZN(new_n512));
  AOI211_X1 g311(.A(new_n510), .B(new_n512), .C1(new_n336), .C2(new_n414), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT88), .B1(new_n502), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT36), .ZN(new_n515));
  INV_X1    g314(.A(new_n447), .ZN(new_n516));
  INV_X1    g315(.A(new_n448), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n447), .A2(KEYINPUT36), .A3(new_n448), .ZN(new_n519));
  INV_X1    g318(.A(new_n474), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n518), .A2(new_n519), .B1(new_n415), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n510), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n481), .A2(new_n401), .A3(new_n511), .A4(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT88), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n523), .A2(new_n524), .A3(new_n474), .A4(new_n501), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n514), .A2(new_n521), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n245), .B1(new_n485), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT97), .ZN(new_n528));
  XNOR2_X1  g327(.A(G120gat), .B(G148gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(new_n257), .ZN(new_n530));
  XOR2_X1   g329(.A(new_n530), .B(G204gat), .Z(new_n531));
  XNOR2_X1  g330(.A(G57gat), .B(G64gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(KEYINPUT93), .ZN(new_n533));
  NAND2_X1  g332(.A1(G71gat), .A2(G78gat), .ZN(new_n534));
  OR2_X1    g333(.A1(G71gat), .A2(G78gat), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT9), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n534), .B(new_n535), .C1(new_n532), .C2(new_n536), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G99gat), .A2(G106gat), .ZN(new_n541));
  INV_X1    g340(.A(G85gat), .ZN(new_n542));
  AOI22_X1  g341(.A1(KEYINPUT8), .A2(new_n541), .B1(new_n542), .B2(new_n328), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT7), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n544), .B1(new_n542), .B2(new_n328), .ZN(new_n545));
  NAND3_X1  g344(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n543), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G99gat), .B(G106gat), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n547), .B(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT94), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n547), .B(new_n548), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n553), .A2(KEYINPUT94), .ZN(new_n554));
  OAI211_X1 g353(.A(KEYINPUT10), .B(new_n540), .C1(new_n552), .C2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT96), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n550), .B(new_n551), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n558), .A2(KEYINPUT96), .A3(KEYINPUT10), .A4(new_n540), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n547), .A2(KEYINPUT95), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n540), .A2(new_n553), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT10), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n538), .A2(new_n560), .A3(new_n539), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(new_n550), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n557), .A2(new_n559), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G230gat), .A2(G233gat), .ZN(new_n567));
  AND2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n567), .B1(new_n561), .B2(new_n564), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n528), .B(new_n531), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n531), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n569), .B1(new_n566), .B2(new_n567), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n571), .B1(new_n572), .B2(KEYINPUT97), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  AND2_X1   g374(.A1(G232gat), .A2(G233gat), .ZN(new_n576));
  AOI22_X1  g375(.A1(new_n558), .A2(new_n222), .B1(KEYINPUT41), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n210), .A2(new_n218), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n577), .B1(new_n578), .B2(new_n558), .ZN(new_n579));
  XNOR2_X1  g378(.A(G134gat), .B(G162gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n576), .A2(KEYINPUT41), .ZN(new_n582));
  XNOR2_X1  g381(.A(G190gat), .B(G218gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n580), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n577), .B(new_n585), .C1(new_n578), .C2(new_n558), .ZN(new_n586));
  AND3_X1   g385(.A1(new_n581), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n584), .B1(new_n581), .B2(new_n586), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n540), .A2(KEYINPUT21), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n592));
  XOR2_X1   g391(.A(new_n591), .B(new_n592), .Z(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n540), .A2(KEYINPUT21), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(new_n217), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(G183gat), .ZN(new_n597));
  AND2_X1   g396(.A1(G231gat), .A2(G233gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G127gat), .B(G155gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(G211gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n599), .A2(new_n601), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n594), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n604), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n606), .A2(new_n593), .A3(new_n602), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n590), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n527), .A2(new_n575), .A3(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n609), .A2(new_n411), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n610), .B(G1gat), .Z(G1324gat));
  INV_X1    g410(.A(KEYINPUT42), .ZN(new_n612));
  INV_X1    g411(.A(new_n481), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n612), .B1(new_n615), .B2(G8gat), .ZN(new_n616));
  XOR2_X1   g415(.A(KEYINPUT16), .B(G8gat), .Z(new_n617));
  NAND2_X1  g416(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n617), .A2(KEYINPUT98), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n617), .B1(KEYINPUT98), .B2(KEYINPUT42), .ZN(new_n621));
  AOI22_X1  g420(.A1(new_n616), .A2(new_n618), .B1(new_n620), .B2(new_n621), .ZN(G1325gat));
  INV_X1    g421(.A(G15gat), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n516), .A2(new_n517), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n623), .B1(new_n609), .B2(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n626), .B(KEYINPUT99), .Z(new_n627));
  NAND2_X1  g426(.A1(new_n518), .A2(new_n519), .ZN(new_n628));
  NOR3_X1   g427(.A1(new_n609), .A2(new_n623), .A3(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n627), .A2(new_n629), .ZN(G1326gat));
  NOR2_X1   g429(.A1(new_n609), .A2(new_n474), .ZN(new_n631));
  XOR2_X1   g430(.A(KEYINPUT43), .B(G22gat), .Z(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT100), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n631), .B(new_n633), .ZN(G1327gat));
  AND2_X1   g433(.A1(new_n605), .A2(new_n607), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n636), .A2(new_n574), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(KEYINPUT101), .B1(new_n638), .B2(new_n589), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT101), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n637), .A2(new_n640), .A3(new_n590), .ZN(new_n641));
  AND3_X1   g440(.A1(new_n527), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(G29gat), .ZN(new_n643));
  INV_X1    g442(.A(new_n411), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT45), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n589), .B(KEYINPUT103), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n647), .A2(KEYINPUT44), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n485), .A2(new_n526), .A3(KEYINPUT102), .ZN(new_n649));
  AOI21_X1  g448(.A(KEYINPUT102), .B1(new_n485), .B2(new_n526), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n485), .A2(new_n526), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(new_n590), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(KEYINPUT44), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n636), .A2(new_n574), .A3(new_n245), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(G29gat), .B1(new_n657), .B2(new_n411), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n646), .A2(new_n658), .ZN(G1328gat));
  INV_X1    g458(.A(new_n642), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n660), .A2(G36gat), .A3(new_n613), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT46), .ZN(new_n662));
  OAI21_X1  g461(.A(G36gat), .B1(new_n657), .B2(new_n613), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(G1329gat));
  INV_X1    g463(.A(new_n628), .ZN(new_n665));
  INV_X1    g464(.A(new_n648), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT102), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n485), .A2(new_n526), .A3(KEYINPUT102), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n666), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n589), .B1(new_n485), .B2(new_n526), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT44), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OAI211_X1 g472(.A(new_n665), .B(new_n656), .C1(new_n670), .C2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(G43gat), .ZN(new_n675));
  AOI21_X1  g474(.A(KEYINPUT47), .B1(new_n675), .B2(KEYINPUT105), .ZN(new_n676));
  INV_X1    g475(.A(G43gat), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n642), .A2(KEYINPUT104), .A3(new_n677), .A4(new_n624), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT104), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n527), .A2(new_n639), .A3(new_n624), .A4(new_n641), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n679), .B1(new_n680), .B2(G43gat), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n675), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n676), .A2(new_n683), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n682), .B(new_n675), .C1(KEYINPUT105), .C2(KEYINPUT47), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(G1330gat));
  NAND4_X1  g485(.A1(new_n655), .A2(G50gat), .A3(new_n520), .A4(new_n656), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n660), .A2(new_n474), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n687), .B1(G50gat), .B2(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g489(.A1(new_n668), .A2(new_n669), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n608), .A2(new_n574), .A3(new_n245), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n692), .B(KEYINPUT106), .Z(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(new_n644), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g496(.A1(new_n694), .A2(new_n613), .ZN(new_n698));
  NOR2_X1   g497(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n699));
  AND2_X1   g498(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n701), .B1(new_n698), .B2(new_n699), .ZN(G1333gat));
  NAND3_X1  g501(.A1(new_n695), .A2(G71gat), .A3(new_n665), .ZN(new_n703));
  INV_X1    g502(.A(G71gat), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n704), .B1(new_n694), .B2(new_n625), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g506(.A1(new_n695), .A2(new_n520), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(G78gat), .ZN(G1335gat));
  INV_X1    g508(.A(KEYINPUT107), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n636), .A2(new_n244), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n655), .A2(new_n574), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n710), .B1(new_n712), .B2(new_n411), .ZN(new_n713));
  INV_X1    g512(.A(new_n711), .ZN(new_n714));
  AOI211_X1 g513(.A(new_n575), .B(new_n714), .C1(new_n651), .C2(new_n654), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n715), .A2(KEYINPUT107), .A3(new_n644), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n713), .A2(new_n716), .A3(G85gat), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n652), .A2(new_n590), .A3(new_n711), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT51), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n671), .A2(KEYINPUT51), .A3(new_n711), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n720), .A2(KEYINPUT108), .A3(new_n721), .ZN(new_n722));
  OR3_X1    g521(.A1(new_n718), .A2(KEYINPUT108), .A3(new_n719), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n724), .A2(new_n575), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n725), .A2(new_n542), .A3(new_n644), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n717), .A2(new_n726), .ZN(G1336gat));
  AOI21_X1  g526(.A(new_n328), .B1(new_n715), .B2(new_n481), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n613), .A2(G92gat), .ZN(new_n729));
  AND4_X1   g528(.A1(KEYINPUT51), .A2(new_n652), .A3(new_n590), .A4(new_n711), .ZN(new_n730));
  XOR2_X1   g529(.A(KEYINPUT109), .B(KEYINPUT51), .Z(new_n731));
  AOI21_X1  g530(.A(new_n731), .B1(new_n671), .B2(new_n711), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n574), .B(new_n729), .C1(new_n730), .C2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT110), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n731), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n718), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n721), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n738), .A2(KEYINPUT110), .A3(new_n574), .A4(new_n729), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(KEYINPUT52), .B1(new_n728), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(G92gat), .B1(new_n712), .B2(new_n613), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT52), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n722), .A2(new_n723), .A3(new_n574), .A4(new_n729), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n741), .A2(new_n745), .ZN(G1337gat));
  NAND3_X1  g545(.A1(new_n725), .A2(new_n427), .A3(new_n624), .ZN(new_n747));
  OAI21_X1  g546(.A(G99gat), .B1(new_n712), .B2(new_n628), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(G1338gat));
  NAND4_X1  g548(.A1(new_n655), .A2(new_n574), .A3(new_n520), .A4(new_n711), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n575), .A2(G106gat), .A3(new_n474), .ZN(new_n751));
  AOI22_X1  g550(.A1(new_n750), .A2(G106gat), .B1(new_n738), .B2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT53), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n750), .A2(G106gat), .ZN(new_n754));
  INV_X1    g553(.A(new_n751), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n753), .B1(new_n724), .B2(new_n755), .ZN(new_n756));
  OAI22_X1  g555(.A1(new_n752), .A2(new_n753), .B1(new_n754), .B2(new_n756), .ZN(G1339gat));
  NAND3_X1  g556(.A1(new_n608), .A2(new_n575), .A3(new_n245), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n566), .A2(new_n567), .ZN(new_n759));
  INV_X1    g558(.A(new_n567), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n557), .A2(new_n559), .A3(new_n760), .A4(new_n565), .ZN(new_n761));
  AND3_X1   g560(.A1(new_n759), .A2(KEYINPUT54), .A3(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n531), .B1(new_n759), .B2(KEYINPUT54), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AOI22_X1  g563(.A1(new_n764), .A2(KEYINPUT55), .B1(new_n572), .B2(new_n571), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT54), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n571), .B1(new_n568), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n759), .A2(KEYINPUT54), .A3(new_n761), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT55), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n230), .B1(new_n229), .B2(new_n231), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n220), .B1(new_n219), .B2(new_n223), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n239), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(KEYINPUT111), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT111), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n775), .B(new_n239), .C1(new_n771), .C2(new_n772), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n774), .A2(new_n243), .A3(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n765), .A2(new_n770), .A3(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n778), .A2(new_n647), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n574), .ZN(new_n780));
  OR2_X1    g579(.A1(new_n780), .A2(KEYINPUT112), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n765), .A2(new_n244), .A3(new_n770), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(KEYINPUT112), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n779), .B1(new_n784), .B2(new_n647), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n758), .B1(new_n785), .B2(new_n636), .ZN(new_n786));
  INV_X1    g585(.A(new_n475), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n786), .A2(new_n644), .A3(new_n613), .A4(new_n787), .ZN(new_n788));
  OR2_X1    g587(.A1(new_n788), .A2(KEYINPUT113), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(KEYINPUT113), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n245), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n244), .A2(new_n357), .ZN(new_n792));
  XOR2_X1   g591(.A(new_n792), .B(KEYINPUT114), .Z(new_n793));
  OAI22_X1  g592(.A1(new_n791), .A2(new_n357), .B1(new_n788), .B2(new_n793), .ZN(G1340gat));
  AOI21_X1  g593(.A(new_n575), .B1(new_n789), .B2(new_n790), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n574), .A2(new_n355), .ZN(new_n796));
  OAI22_X1  g595(.A1(new_n795), .A2(new_n355), .B1(new_n788), .B2(new_n796), .ZN(G1341gat));
  INV_X1    g596(.A(KEYINPUT115), .ZN(new_n798));
  OR3_X1    g597(.A1(new_n788), .A2(G127gat), .A3(new_n635), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n635), .B1(new_n789), .B2(new_n790), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n798), .B(new_n799), .C1(new_n800), .C2(new_n362), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n788), .A2(KEYINPUT113), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n788), .A2(KEYINPUT113), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n636), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(G127gat), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n798), .B1(new_n806), .B2(new_n799), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n802), .A2(new_n807), .ZN(G1342gat));
  NOR3_X1   g607(.A1(new_n788), .A2(G134gat), .A3(new_n589), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT56), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n811), .B(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n590), .B1(new_n803), .B2(new_n804), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(G134gat), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n813), .B(new_n815), .C1(new_n810), .C2(new_n809), .ZN(G1343gat));
  INV_X1    g615(.A(KEYINPUT58), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n786), .A2(new_n644), .A3(new_n520), .A4(new_n628), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n818), .A2(new_n481), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n819), .A2(new_n341), .A3(new_n244), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT118), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n817), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT57), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n786), .A2(new_n823), .A3(new_n520), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n767), .A2(KEYINPUT55), .A3(new_n768), .ZN(new_n825));
  XOR2_X1   g624(.A(KEYINPUT117), .B(KEYINPUT55), .Z(new_n826));
  OAI21_X1  g625(.A(new_n826), .B1(new_n762), .B2(new_n763), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n572), .A2(new_n571), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n244), .A2(new_n825), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n590), .B1(new_n829), .B2(new_n780), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n635), .B1(new_n779), .B2(new_n830), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n831), .A2(new_n758), .ZN(new_n832));
  OAI21_X1  g631(.A(KEYINPUT57), .B1(new_n832), .B2(new_n474), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n665), .A2(new_n411), .A3(new_n481), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n824), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(G141gat), .B1(new_n835), .B2(new_n245), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n820), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n822), .B(new_n837), .ZN(G1344gat));
  NAND3_X1  g637(.A1(new_n819), .A2(new_n343), .A3(new_n574), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT59), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n828), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n774), .A2(new_n243), .A3(new_n776), .ZN(new_n842));
  NOR4_X1   g641(.A1(new_n841), .A2(new_n769), .A3(new_n589), .A4(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n635), .B1(new_n830), .B2(new_n843), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n844), .A2(KEYINPUT119), .A3(new_n758), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT119), .B1(new_n844), .B2(new_n758), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n845), .A2(new_n846), .A3(new_n474), .ZN(new_n847));
  OAI21_X1  g646(.A(KEYINPUT120), .B1(new_n847), .B2(KEYINPUT57), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n786), .A2(KEYINPUT57), .A3(new_n520), .ZN(new_n849));
  INV_X1    g648(.A(new_n846), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n844), .A2(KEYINPUT119), .A3(new_n758), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n850), .A2(new_n520), .A3(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n852), .A2(new_n853), .A3(new_n823), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n848), .A2(new_n849), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n574), .A3(new_n834), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n840), .B1(new_n856), .B2(G148gat), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n840), .B1(new_n835), .B2(new_n575), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n858), .A2(new_n343), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n839), .B1(new_n857), .B2(new_n859), .ZN(G1345gat));
  OAI21_X1  g659(.A(G155gat), .B1(new_n835), .B2(new_n635), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n819), .A2(new_n337), .A3(new_n636), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(G1346gat));
  OAI21_X1  g662(.A(G162gat), .B1(new_n835), .B2(new_n647), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n819), .A2(new_n338), .A3(new_n590), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(G1347gat));
  AND2_X1   g665(.A1(new_n786), .A2(new_n411), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n613), .A2(new_n475), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(G169gat), .B1(new_n869), .B2(new_n245), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(KEYINPUT121), .B1(new_n613), .B2(new_n475), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n786), .A2(new_n411), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n875), .A2(G169gat), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n871), .B1(new_n876), .B2(new_n244), .ZN(new_n877));
  NOR4_X1   g676(.A1(new_n875), .A2(KEYINPUT122), .A3(G169gat), .A4(new_n245), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n870), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n879), .B(new_n880), .ZN(G1348gat));
  NOR3_X1   g680(.A1(new_n869), .A2(new_n575), .A3(new_n278), .ZN(new_n882));
  INV_X1    g681(.A(new_n875), .ZN(new_n883));
  AOI21_X1  g682(.A(G176gat), .B1(new_n883), .B2(new_n574), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n882), .A2(new_n884), .ZN(G1349gat));
  OAI21_X1  g684(.A(G183gat), .B1(new_n869), .B2(new_n635), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n636), .A2(new_n297), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n886), .B1(new_n875), .B2(new_n887), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g688(.A(G190gat), .B1(new_n869), .B2(new_n589), .ZN(new_n890));
  XOR2_X1   g689(.A(KEYINPUT124), .B(KEYINPUT61), .Z(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  OR2_X1    g691(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n647), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n883), .A2(new_n298), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n890), .A2(new_n892), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n893), .A2(new_n895), .A3(new_n896), .ZN(G1351gat));
  NOR2_X1   g696(.A1(new_n665), .A2(new_n613), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n411), .ZN(new_n899));
  XOR2_X1   g698(.A(new_n899), .B(KEYINPUT126), .Z(new_n900));
  NAND3_X1  g699(.A1(new_n855), .A2(new_n244), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(G197gat), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n665), .A2(new_n613), .A3(new_n474), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(KEYINPUT125), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n903), .A2(KEYINPUT125), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n867), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n906), .A2(G197gat), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n902), .B1(new_n245), .B2(new_n907), .ZN(G1352gat));
  NOR3_X1   g707(.A1(new_n906), .A2(G204gat), .A3(new_n575), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(KEYINPUT62), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n855), .A2(new_n574), .A3(new_n900), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(G204gat), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(G1353gat));
  NAND3_X1  g712(.A1(new_n855), .A2(new_n636), .A3(new_n900), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(G211gat), .ZN(new_n915));
  NAND2_X1  g714(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT127), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT63), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n915), .A2(new_n916), .A3(new_n919), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n914), .A2(new_n917), .A3(new_n918), .A4(G211gat), .ZN(new_n921));
  INV_X1    g720(.A(new_n906), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(new_n248), .A3(new_n636), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n920), .A2(new_n921), .A3(new_n923), .ZN(G1354gat));
  NAND3_X1  g723(.A1(new_n922), .A2(new_n249), .A3(new_n894), .ZN(new_n925));
  AND3_X1   g724(.A1(new_n855), .A2(new_n590), .A3(new_n900), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n926), .B2(new_n249), .ZN(G1355gat));
endmodule


