//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 1 0 1 0 1 0 1 0 1 0 1 0 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1 0 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 0 0 0 1 1 0 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1188, new_n1189,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G77), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR3_X1   g0009(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  AOI22_X1  g0012(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G226), .ZN(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT66), .B(G77), .ZN(new_n215));
  INV_X1    g0015(.A(G244), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n213), .B1(new_n201), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  OR2_X1    g0017(.A1(new_n217), .A2(KEYINPUT67), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G58), .A2(G232), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(KEYINPUT67), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G87), .A2(G250), .ZN(new_n221));
  NAND4_X1  g0021(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n222), .B1(G97), .B2(G257), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G107), .A2(G264), .ZN(new_n224));
  AOI22_X1  g0024(.A1(new_n223), .A2(new_n224), .B1(G1), .B2(G20), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT1), .Z(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G20), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT65), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n202), .A2(new_n203), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G50), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n212), .B(new_n226), .C1(new_n230), .C2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  INV_X1    g0040(.A(G264), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G270), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n239), .B(new_n243), .Z(G358));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(new_n201), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G58), .ZN(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(KEYINPUT10), .ZN(new_n252));
  INV_X1    g0052(.A(G200), .ZN(new_n253));
  OR2_X1    g0053(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n254));
  NAND2_X1  g0054(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT3), .B(G33), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n256), .A2(new_n257), .A3(G222), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G1698), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT70), .ZN(new_n266));
  XNOR2_X1  g0066(.A(new_n265), .B(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G223), .ZN(new_n268));
  OAI221_X1 g0068(.A(new_n258), .B1(new_n215), .B2(new_n257), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G41), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n228), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n274));
  INV_X1    g0074(.A(G274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT68), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n227), .B1(new_n277), .B2(new_n270), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n278), .B1(new_n277), .B2(new_n270), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n274), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n276), .B1(new_n281), .B2(G226), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n253), .B1(new_n273), .B2(new_n282), .ZN(new_n283));
  AND2_X1   g0083(.A1(new_n273), .A2(new_n282), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n283), .B1(G190), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n227), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT8), .B(G58), .ZN(new_n289));
  NOR3_X1   g0089(.A1(new_n289), .A2(G20), .A3(new_n259), .ZN(new_n290));
  NOR2_X1   g0090(.A1(G20), .A2(G33), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n290), .B1(G150), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n205), .A2(G20), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n288), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n208), .A2(G20), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n288), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n294), .B1(G50), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G13), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n201), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT9), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n298), .A2(new_n301), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT9), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n252), .B1(new_n285), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n304), .A2(KEYINPUT73), .A3(new_n306), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(KEYINPUT73), .B1(new_n304), .B2(new_n306), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT75), .ZN(new_n313));
  XNOR2_X1  g0113(.A(KEYINPUT74), .B(KEYINPUT10), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n312), .A2(new_n313), .A3(new_n285), .A4(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT73), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n307), .A2(new_n316), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n317), .A2(new_n285), .A3(new_n314), .A4(new_n309), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT75), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n308), .B1(new_n315), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n215), .ZN(new_n321));
  XOR2_X1   g0121(.A(KEYINPUT15), .B(G87), .Z(new_n322));
  NOR2_X1   g0122(.A1(new_n259), .A2(G20), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n321), .A2(G20), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n289), .B(KEYINPUT71), .ZN(new_n325));
  INV_X1    g0125(.A(new_n291), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n327), .A2(new_n287), .B1(G77), .B2(new_n297), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n300), .A2(new_n215), .ZN(new_n329));
  XOR2_X1   g0129(.A(new_n329), .B(KEYINPUT72), .Z(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n256), .A2(new_n257), .A3(G232), .ZN(new_n332));
  INV_X1    g0132(.A(G238), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n332), .B1(new_n267), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G107), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n257), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n272), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n276), .B1(new_n281), .B2(G244), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n331), .B1(new_n340), .B2(G190), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(new_n253), .B2(new_n340), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n284), .A2(G169), .ZN(new_n344));
  INV_X1    g0144(.A(G179), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n344), .B1(new_n345), .B2(new_n284), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n346), .A2(new_n305), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n340), .A2(new_n345), .ZN(new_n348));
  INV_X1    g0148(.A(G169), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n339), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n348), .A2(new_n331), .A3(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NOR4_X1   g0152(.A1(new_n320), .A2(new_n343), .A3(new_n347), .A4(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT76), .ZN(new_n354));
  INV_X1    g0154(.A(G97), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n259), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  AND2_X1   g0157(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n358));
  NOR2_X1   g0158(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n359));
  OAI21_X1  g0159(.A(G226), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G232), .A2(G1698), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n354), .B(new_n357), .C1(new_n362), .C2(new_n263), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n263), .B1(new_n360), .B2(new_n361), .ZN(new_n364));
  OAI21_X1  g0164(.A(KEYINPUT76), .B1(new_n364), .B2(new_n356), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n363), .A2(new_n365), .A3(new_n272), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT13), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n276), .B1(new_n281), .B2(G238), .ZN(new_n368));
  AND3_X1   g0168(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n367), .B1(new_n366), .B2(new_n368), .ZN(new_n370));
  OAI21_X1  g0170(.A(G169), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(KEYINPUT14), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n369), .A2(new_n370), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(G179), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT14), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n375), .B(G169), .C1(new_n369), .C2(new_n370), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n372), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n300), .A2(new_n203), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT12), .B1(new_n378), .B2(KEYINPUT77), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(KEYINPUT77), .ZN(new_n380));
  XNOR2_X1  g0180(.A(new_n379), .B(new_n380), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n323), .A2(G77), .B1(new_n291), .B2(G50), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n382), .B1(new_n209), .B2(G68), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n287), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT11), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n384), .A2(new_n385), .B1(G68), .B2(new_n297), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n381), .B(new_n386), .C1(new_n385), .C2(new_n384), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n377), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n387), .B1(new_n373), .B2(G190), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n253), .B2(new_n373), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  XOR2_X1   g0191(.A(new_n391), .B(KEYINPUT78), .Z(new_n392));
  NAND2_X1  g0192(.A1(new_n256), .A2(G223), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(new_n214), .B2(new_n264), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n261), .A2(G33), .ZN(new_n395));
  OAI21_X1  g0195(.A(KEYINPUT79), .B1(new_n259), .B2(KEYINPUT3), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT79), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n397), .A2(new_n261), .A3(G33), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n395), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n394), .A2(new_n399), .B1(G33), .B2(G87), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n400), .A2(new_n271), .ZN(new_n401));
  OAI22_X1  g0201(.A1(new_n280), .A2(new_n236), .B1(new_n275), .B2(new_n274), .ZN(new_n402));
  OAI21_X1  g0202(.A(G169), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n402), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(new_n271), .B2(new_n400), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n403), .B1(new_n345), .B2(new_n405), .ZN(new_n406));
  XNOR2_X1  g0206(.A(KEYINPUT82), .B(KEYINPUT18), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n397), .B1(new_n261), .B2(G33), .ZN(new_n408));
  NOR3_X1   g0208(.A1(new_n259), .A2(KEYINPUT79), .A3(KEYINPUT3), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n260), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT7), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(new_n411), .A3(new_n209), .ZN(new_n412));
  OAI21_X1  g0212(.A(KEYINPUT7), .B1(new_n399), .B2(G20), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(new_n413), .A3(G68), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT80), .B1(new_n202), .B2(new_n203), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT80), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n416), .A2(G58), .A3(G68), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(new_n231), .A3(new_n417), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n418), .A2(G20), .B1(G159), .B2(new_n291), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n414), .A2(KEYINPUT16), .A3(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT16), .ZN(new_n421));
  INV_X1    g0221(.A(new_n419), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n411), .B1(new_n257), .B2(G20), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n263), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n203), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n421), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n420), .A2(new_n287), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT81), .ZN(new_n428));
  INV_X1    g0228(.A(new_n300), .ZN(new_n429));
  MUX2_X1   g0229(.A(new_n296), .B(new_n429), .S(new_n289), .Z(new_n430));
  AND3_X1   g0230(.A1(new_n427), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n428), .B1(new_n427), .B2(new_n430), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n406), .B(new_n407), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n406), .B1(new_n431), .B2(new_n432), .ZN(new_n434));
  INV_X1    g0234(.A(new_n407), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT17), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n427), .A2(new_n430), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT83), .ZN(new_n439));
  OAI21_X1  g0239(.A(G200), .B1(new_n401), .B2(new_n402), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n404), .B(G190), .C1(new_n271), .C2(new_n400), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n438), .A2(new_n439), .A3(new_n440), .A4(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n440), .A2(new_n427), .A3(new_n441), .A4(new_n430), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(KEYINPUT83), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n437), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n443), .A2(KEYINPUT17), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n433), .B(new_n436), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n392), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n353), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(G116), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n300), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n208), .A2(G33), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n287), .B1(KEYINPUT84), .B2(new_n453), .ZN(new_n454));
  OR2_X1    g0254(.A1(new_n453), .A2(KEYINPUT84), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n454), .A2(new_n429), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(G20), .B1(G33), .B2(G283), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n457), .B1(G33), .B2(new_n355), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n458), .B(new_n287), .C1(new_n209), .C2(G116), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT20), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n459), .A2(new_n460), .ZN(new_n462));
  OAI221_X1 g0262(.A(new_n452), .B1(new_n456), .B2(new_n451), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(G45), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(G1), .ZN(new_n465));
  AND2_X1   g0265(.A1(KEYINPUT5), .A2(G41), .ZN(new_n466));
  NOR2_X1   g0266(.A1(KEYINPUT5), .A2(G41), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n279), .A2(G270), .A3(new_n468), .ZN(new_n469));
  OR2_X1    g0269(.A1(new_n468), .A2(new_n275), .ZN(new_n470));
  INV_X1    g0270(.A(G303), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n257), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(G257), .B1(new_n358), .B2(new_n359), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n473), .B1(new_n241), .B2(new_n264), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n472), .B1(new_n474), .B2(new_n399), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n469), .B(new_n470), .C1(new_n475), .C2(new_n271), .ZN(new_n476));
  XNOR2_X1  g0276(.A(new_n476), .B(KEYINPUT87), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n463), .B1(new_n477), .B2(G200), .ZN(new_n478));
  INV_X1    g0278(.A(G190), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n478), .B1(new_n479), .B2(new_n477), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n396), .A2(new_n398), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n481), .A2(KEYINPUT22), .A3(G87), .A4(new_n260), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G116), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n209), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n257), .A2(new_n209), .A3(G87), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT22), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n209), .A2(G107), .ZN(new_n489));
  XNOR2_X1  g0289(.A(new_n489), .B(KEYINPUT23), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n485), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT24), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n485), .A2(KEYINPUT24), .A3(new_n488), .A4(new_n490), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n493), .A2(new_n287), .A3(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n456), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G107), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n300), .A2(new_n335), .ZN(new_n498));
  XOR2_X1   g0298(.A(new_n498), .B(KEYINPUT25), .Z(new_n499));
  NAND3_X1  g0299(.A1(new_n495), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n256), .A2(G250), .B1(G257), .B2(G1698), .ZN(new_n501));
  INV_X1    g0301(.A(G294), .ZN(new_n502));
  OAI22_X1  g0302(.A1(new_n501), .A2(new_n410), .B1(new_n259), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n272), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n279), .A2(G264), .A3(new_n468), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n504), .A2(new_n470), .A3(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n506), .A2(G179), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n507), .B1(new_n349), .B2(new_n506), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n500), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n477), .A2(KEYINPUT21), .A3(G169), .A4(new_n463), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n476), .A2(new_n345), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n463), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n474), .A2(new_n399), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n272), .B1(new_n514), .B2(new_n472), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n515), .A2(KEYINPUT87), .A3(new_n469), .A4(new_n470), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT87), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n476), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n516), .A2(G169), .A3(new_n518), .A4(new_n463), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT21), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n511), .A2(new_n513), .A3(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n510), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n456), .A2(new_n355), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n423), .A2(new_n424), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(G107), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n291), .A2(G77), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n335), .A2(KEYINPUT6), .A3(G97), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n355), .A2(new_n335), .ZN(new_n529));
  NOR2_X1   g0329(.A1(G97), .A2(G107), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n528), .B1(new_n531), .B2(KEYINPUT6), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(G20), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n526), .A2(new_n527), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n524), .B1(new_n534), .B2(new_n287), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(G97), .B2(new_n429), .ZN(new_n536));
  AND3_X1   g0336(.A1(new_n279), .A2(G257), .A3(new_n468), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n265), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT4), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n256), .A2(G244), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n539), .B1(new_n410), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n263), .A2(new_n539), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT85), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n542), .A2(new_n543), .A3(G244), .A4(new_n256), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n257), .A2(KEYINPUT4), .ZN(new_n545));
  OAI21_X1  g0345(.A(KEYINPUT85), .B1(new_n540), .B2(new_n545), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n538), .A2(new_n541), .A3(new_n544), .A4(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n537), .B1(new_n547), .B2(new_n272), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n548), .A2(new_n345), .A3(new_n470), .ZN(new_n549));
  INV_X1    g0349(.A(new_n470), .ZN(new_n550));
  AOI211_X1 g0350(.A(new_n550), .B(new_n537), .C1(new_n547), .C2(new_n272), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n536), .B(new_n549), .C1(G169), .C2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n548), .A2(G190), .A3(new_n470), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n429), .A2(G97), .ZN(new_n554));
  AOI211_X1 g0354(.A(new_n554), .B(new_n524), .C1(new_n534), .C2(new_n287), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n553), .B(new_n555), .C1(new_n253), .C2(new_n551), .ZN(new_n556));
  MUX2_X1   g0356(.A(G250), .B(G274), .S(new_n465), .Z(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n279), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n399), .A2(G244), .A3(G1698), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(KEYINPUT86), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n399), .A2(G238), .A3(new_n256), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT86), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n399), .A2(new_n563), .A3(G244), .A4(G1698), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n561), .A2(new_n483), .A3(new_n562), .A4(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n559), .B1(new_n565), .B2(new_n272), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n345), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n399), .A2(new_n209), .A3(G68), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT19), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(new_n357), .B2(G20), .ZN(new_n570));
  AOI21_X1  g0370(.A(G20), .B1(new_n356), .B2(KEYINPUT19), .ZN(new_n571));
  NOR3_X1   g0371(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n568), .B(new_n570), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n322), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n573), .A2(new_n287), .B1(new_n574), .B2(new_n300), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n574), .B2(new_n456), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n567), .B(new_n576), .C1(G169), .C2(new_n566), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n496), .A2(G87), .ZN(new_n578));
  AND2_X1   g0378(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n565), .A2(new_n272), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n580), .A2(G190), .A3(new_n558), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n579), .B(new_n581), .C1(new_n253), .C2(new_n566), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n552), .A2(new_n556), .A3(new_n577), .A4(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n506), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n584), .A2(new_n253), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n506), .A2(new_n479), .ZN(new_n586));
  NOR3_X1   g0386(.A1(new_n500), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n450), .A2(new_n480), .A3(new_n523), .A4(new_n588), .ZN(new_n589));
  XNOR2_X1  g0389(.A(new_n589), .B(KEYINPUT88), .ZN(G372));
  NAND2_X1  g0390(.A1(new_n427), .A2(new_n430), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n406), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g0392(.A(new_n592), .B(KEYINPUT18), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n442), .A2(new_n444), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n446), .B1(new_n595), .B2(KEYINPUT17), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n596), .B1(new_n351), .B2(new_n388), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n390), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n320), .B1(new_n594), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n588), .B1(new_n522), .B2(new_n510), .ZN(new_n600));
  INV_X1    g0400(.A(new_n577), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n577), .A2(new_n582), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n552), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n601), .B1(new_n605), .B2(KEYINPUT26), .ZN(new_n606));
  XNOR2_X1  g0406(.A(KEYINPUT89), .B(KEYINPUT26), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n600), .B(new_n606), .C1(new_n605), .C2(new_n607), .ZN(new_n608));
  AOI211_X1 g0408(.A(new_n347), .B(new_n599), .C1(new_n450), .C2(new_n608), .ZN(new_n609));
  XOR2_X1   g0409(.A(new_n609), .B(KEYINPUT90), .Z(G369));
  NOR2_X1   g0410(.A1(new_n299), .A2(G20), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n208), .ZN(new_n612));
  OR2_X1    g0412(.A1(new_n612), .A2(KEYINPUT27), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(KEYINPUT27), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(G213), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(G343), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n463), .A2(new_n617), .ZN(new_n618));
  OR2_X1    g0418(.A1(new_n522), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n522), .A2(new_n618), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(new_n480), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(G330), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OR3_X1    g0423(.A1(new_n500), .A2(new_n585), .A3(new_n586), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n500), .A2(new_n617), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n510), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n509), .A2(new_n617), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n617), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n522), .A2(new_n630), .ZN(new_n631));
  OAI22_X1  g0431(.A1(new_n626), .A2(new_n631), .B1(new_n509), .B2(new_n617), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n629), .A2(new_n633), .ZN(G399));
  INV_X1    g0434(.A(new_n210), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n635), .A2(G41), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(G1), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n572), .A2(new_n451), .ZN(new_n639));
  OAI22_X1  g0439(.A1(new_n638), .A2(new_n639), .B1(new_n232), .B2(new_n637), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n640), .B(KEYINPUT28), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n608), .A2(new_n630), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n642), .A2(KEYINPUT29), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n605), .A2(new_n607), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n601), .A2(KEYINPUT92), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n602), .A2(new_n552), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT26), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n601), .A2(KEYINPUT92), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n644), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(KEYINPUT93), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT93), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n644), .A2(new_n648), .A3(new_n652), .A4(new_n649), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n651), .A2(new_n600), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n630), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n643), .B1(new_n655), .B2(KEYINPUT29), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n584), .A2(new_n566), .A3(new_n512), .A4(new_n548), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT30), .ZN(new_n658));
  XNOR2_X1  g0458(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n548), .A2(new_n470), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n477), .A2(new_n506), .A3(new_n660), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n661), .A2(G179), .A3(new_n566), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n617), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT31), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n665), .A2(KEYINPUT91), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n588), .A2(new_n523), .A3(new_n480), .A4(new_n630), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n477), .A2(new_n660), .ZN(new_n668));
  INV_X1    g0468(.A(new_n566), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n668), .A2(new_n345), .A3(new_n506), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n657), .B(KEYINPUT30), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n630), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(KEYINPUT91), .B1(new_n672), .B2(KEYINPUT31), .ZN(new_n673));
  INV_X1    g0473(.A(new_n665), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n666), .B(new_n667), .C1(new_n673), .C2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G330), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n656), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n641), .B1(new_n678), .B2(G1), .ZN(G364));
  NOR2_X1   g0479(.A1(new_n209), .A2(G190), .ZN(new_n680));
  XOR2_X1   g0480(.A(new_n680), .B(KEYINPUT95), .Z(new_n681));
  NAND3_X1  g0481(.A1(new_n681), .A2(new_n345), .A3(new_n253), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n209), .A2(new_n479), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n345), .A2(new_n253), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n683), .A2(G329), .B1(G326), .B2(new_n687), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n479), .A2(G179), .A3(G200), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(new_n209), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n688), .B1(new_n502), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n253), .A2(G179), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n684), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n691), .B1(G303), .B2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n345), .A2(G200), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n684), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G322), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n681), .A2(new_n692), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(G283), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n696), .A2(new_n680), .ZN(new_n703));
  INV_X1    g0503(.A(G311), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n263), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n685), .A2(new_n680), .ZN(new_n706));
  INV_X1    g0506(.A(G317), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n706), .B1(KEYINPUT33), .B2(new_n707), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n707), .A2(KEYINPUT33), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n705), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n695), .A2(new_n699), .A3(new_n702), .A4(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n690), .ZN(new_n712));
  AOI22_X1  g0512(.A1(new_n712), .A2(G97), .B1(new_n694), .B2(G87), .ZN(new_n713));
  OAI221_X1 g0513(.A(new_n713), .B1(new_n202), .B2(new_n697), .C1(new_n203), .C2(new_n706), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n683), .A2(G159), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT32), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n716), .B1(new_n215), .B2(new_n703), .ZN(new_n717));
  AOI211_X1 g0517(.A(new_n714), .B(new_n717), .C1(G50), .C2(new_n687), .ZN(new_n718));
  OAI221_X1 g0518(.A(new_n718), .B1(KEYINPUT32), .B2(new_n715), .C1(new_n335), .C2(new_n700), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n711), .B1(new_n719), .B2(new_n263), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n227), .B1(G20), .B2(new_n349), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n635), .A2(new_n263), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G355), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n247), .A2(new_n464), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n399), .A2(new_n635), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(G45), .B2(new_n232), .ZN(new_n727));
  OAI221_X1 g0527(.A(new_n724), .B1(G116), .B2(new_n210), .C1(new_n725), .C2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(G13), .A2(G33), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(G20), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(new_n721), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n728), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n638), .B1(G45), .B2(new_n611), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n735), .B1(new_n621), .B2(new_n731), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n722), .A2(new_n733), .A3(new_n736), .ZN(new_n737));
  XOR2_X1   g0537(.A(new_n737), .B(KEYINPUT96), .Z(new_n738));
  NAND2_X1  g0538(.A1(new_n621), .A2(new_n622), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n623), .A2(KEYINPUT94), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n623), .A2(KEYINPUT94), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n735), .B(new_n739), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n738), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(G396));
  NOR2_X1   g0545(.A1(new_n351), .A2(new_n617), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n331), .A2(new_n617), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n342), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n747), .B1(new_n749), .B2(new_n352), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT99), .ZN(new_n751));
  MUX2_X1   g0551(.A(new_n750), .B(new_n751), .S(new_n642), .Z(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(new_n676), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n735), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n750), .A2(new_n729), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n721), .A2(new_n729), .ZN(new_n756));
  INV_X1    g0556(.A(G77), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n703), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n701), .A2(G87), .B1(G116), .B2(new_n759), .ZN(new_n760));
  XNOR2_X1  g0560(.A(KEYINPUT97), .B(G283), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI221_X1 g0562(.A(new_n760), .B1(new_n704), .B2(new_n682), .C1(new_n706), .C2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n686), .A2(new_n471), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n263), .B1(new_n693), .B2(new_n335), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT98), .Z(new_n766));
  OAI22_X1  g0566(.A1(new_n690), .A2(new_n355), .B1(new_n697), .B2(new_n502), .ZN(new_n767));
  NOR4_X1   g0567(.A1(new_n763), .A2(new_n764), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(G132), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n682), .A2(new_n769), .B1(new_n201), .B2(new_n693), .ZN(new_n770));
  AOI211_X1 g0570(.A(new_n410), .B(new_n770), .C1(G58), .C2(new_n712), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n701), .A2(G68), .ZN(new_n772));
  INV_X1    g0572(.A(new_n706), .ZN(new_n773));
  AOI22_X1  g0573(.A1(G143), .A2(new_n698), .B1(new_n773), .B2(G150), .ZN(new_n774));
  INV_X1    g0574(.A(G137), .ZN(new_n775));
  INV_X1    g0575(.A(G159), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n774), .B1(new_n775), .B2(new_n686), .C1(new_n776), .C2(new_n703), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT34), .ZN(new_n778));
  AND3_X1   g0578(.A1(new_n771), .A2(new_n772), .A3(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n721), .B1(new_n768), .B2(new_n779), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n755), .A2(new_n734), .A3(new_n758), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n754), .A2(new_n781), .ZN(G384));
  NOR2_X1   g0582(.A1(new_n388), .A2(new_n617), .ZN(new_n783));
  AND2_X1   g0583(.A1(new_n595), .A2(new_n434), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n431), .A2(new_n432), .ZN(new_n785));
  INV_X1    g0585(.A(new_n615), .ZN(new_n786));
  AOI21_X1  g0586(.A(KEYINPUT37), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n420), .A2(new_n287), .ZN(new_n788));
  AOI21_X1  g0588(.A(KEYINPUT16), .B1(new_n414), .B2(new_n419), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n430), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(new_n786), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n406), .A2(new_n790), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n595), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n784), .A2(new_n787), .B1(new_n793), .B2(KEYINPUT37), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n791), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n436), .A2(new_n433), .ZN(new_n797));
  OAI211_X1 g0597(.A(KEYINPUT102), .B(new_n796), .C1(new_n596), .C2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(KEYINPUT102), .B1(new_n447), .B2(new_n796), .ZN(new_n800));
  OAI211_X1 g0600(.A(KEYINPUT38), .B(new_n795), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  AND2_X1   g0601(.A1(new_n785), .A2(new_n786), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n592), .A2(new_n443), .ZN(new_n803));
  OAI21_X1  g0603(.A(KEYINPUT37), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n784), .A2(new_n787), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n802), .B1(new_n596), .B2(new_n593), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT38), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT39), .ZN(new_n811));
  AND3_X1   g0611(.A1(new_n801), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n796), .B1(new_n596), .B2(new_n797), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT102), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(new_n798), .ZN(new_n816));
  AOI21_X1  g0616(.A(KEYINPUT38), .B1(new_n816), .B2(new_n795), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n809), .B(new_n794), .C1(new_n815), .C2(new_n798), .ZN(new_n818));
  OAI21_X1  g0618(.A(KEYINPUT39), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n812), .B1(new_n819), .B2(KEYINPUT103), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n801), .A2(new_n810), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT103), .ZN(new_n822));
  NOR3_X1   g0622(.A1(new_n821), .A2(new_n822), .A3(KEYINPUT39), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n783), .B1(new_n820), .B2(new_n823), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n746), .A2(KEYINPUT100), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n746), .A2(KEYINPUT100), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n825), .B(new_n826), .C1(new_n642), .C2(new_n750), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n387), .A2(new_n617), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n388), .A2(new_n390), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n377), .A2(new_n387), .A3(new_n617), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT101), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n829), .A2(KEYINPUT101), .A3(new_n830), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n827), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n817), .A2(new_n818), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n836), .A2(new_n837), .B1(new_n594), .B2(new_n786), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n824), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n599), .A2(new_n347), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n656), .B2(new_n449), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n840), .B(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n672), .A2(KEYINPUT31), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n667), .A2(new_n665), .A3(new_n844), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n450), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n342), .A2(new_n748), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n746), .B1(new_n847), .B2(new_n351), .ZN(new_n848));
  AND3_X1   g0648(.A1(new_n829), .A2(KEYINPUT101), .A3(new_n830), .ZN(new_n849));
  AOI21_X1  g0649(.A(KEYINPUT101), .B1(new_n829), .B2(new_n830), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n845), .B(new_n848), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT104), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OR2_X1    g0653(.A1(KEYINPUT104), .A2(KEYINPUT40), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n835), .A2(new_n848), .A3(new_n845), .A4(new_n854), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n853), .B(new_n855), .C1(new_n818), .C2(new_n817), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT38), .B1(new_n806), .B2(new_n807), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n794), .B1(new_n815), .B2(new_n798), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n857), .B1(new_n858), .B2(KEYINPUT38), .ZN(new_n859));
  OAI21_X1  g0659(.A(KEYINPUT40), .B1(new_n859), .B2(new_n851), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n846), .B(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n862), .A2(new_n622), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n843), .B(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n208), .B2(new_n611), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n451), .B1(new_n532), .B2(KEYINPUT35), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n866), .B(new_n230), .C1(KEYINPUT35), .C2(new_n532), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(KEYINPUT36), .ZN(new_n868));
  OAI21_X1  g0668(.A(G50), .B1(new_n418), .B2(new_n215), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n201), .A2(new_n203), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n869), .A2(G1), .A3(new_n299), .A4(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n865), .A2(new_n868), .A3(new_n871), .ZN(G367));
  NOR3_X1   g0672(.A1(new_n626), .A2(new_n627), .A3(new_n631), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n552), .A2(new_n556), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n536), .A2(new_n617), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT42), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n604), .B1(new_n877), .B2(new_n510), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n878), .A2(KEYINPUT42), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT106), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR3_X1   g0683(.A1(new_n878), .A2(KEYINPUT106), .A3(KEYINPUT42), .ZN(new_n884));
  OAI221_X1 g0684(.A(new_n879), .B1(new_n617), .B2(new_n880), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT107), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n579), .A2(new_n630), .ZN(new_n887));
  XOR2_X1   g0687(.A(new_n887), .B(KEYINPUT105), .Z(new_n888));
  NOR2_X1   g0688(.A1(new_n888), .A2(new_n603), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(new_n577), .B2(new_n888), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n885), .A2(new_n886), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n891), .B1(new_n885), .B2(new_n886), .ZN(new_n893));
  OAI211_X1 g0693(.A(KEYINPUT43), .B(new_n885), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n893), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT43), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n885), .A2(new_n886), .A3(new_n891), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n604), .A2(new_n617), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n876), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n629), .A2(new_n901), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n894), .A2(new_n898), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n902), .B1(new_n894), .B2(new_n898), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n636), .B(KEYINPUT41), .Z(new_n906));
  INV_X1    g0706(.A(KEYINPUT108), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n633), .A2(KEYINPUT45), .A3(new_n900), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT45), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n632), .B2(new_n901), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  OR3_X1    g0711(.A1(new_n633), .A2(KEYINPUT44), .A3(new_n900), .ZN(new_n912));
  OAI21_X1  g0712(.A(KEYINPUT44), .B1(new_n633), .B2(new_n900), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n629), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n914), .A2(new_n915), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n907), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n631), .B1(new_n626), .B2(new_n627), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT109), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(new_n873), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n623), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n740), .A2(new_n741), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n923), .B1(new_n924), .B2(new_n922), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n677), .A2(new_n925), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n918), .B(new_n926), .C1(new_n907), .C2(new_n916), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n906), .B1(new_n927), .B2(new_n678), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n208), .B1(new_n611), .B2(G45), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n905), .A2(new_n931), .ZN(new_n932));
  AOI22_X1  g0732(.A1(G58), .A2(new_n694), .B1(new_n698), .B2(G150), .ZN(new_n933));
  OAI221_X1 g0733(.A(new_n933), .B1(new_n201), .B2(new_n703), .C1(new_n776), .C2(new_n706), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n934), .B1(G68), .B2(new_n712), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n263), .B1(new_n687), .B2(G143), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n935), .B(new_n936), .C1(new_n775), .C2(new_n682), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(new_n321), .B2(new_n701), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n410), .B1(new_n502), .B2(new_n706), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n701), .B2(G97), .ZN(new_n940));
  OAI221_X1 g0740(.A(new_n940), .B1(new_n335), .B2(new_n690), .C1(new_n703), .C2(new_n762), .ZN(new_n941));
  XOR2_X1   g0741(.A(KEYINPUT110), .B(G317), .Z(new_n942));
  NOR2_X1   g0742(.A1(new_n682), .A2(new_n942), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n686), .A2(new_n704), .B1(new_n697), .B2(new_n471), .ZN(new_n944));
  NOR3_X1   g0744(.A1(new_n941), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n694), .A2(G116), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT46), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n938), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT47), .Z(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n721), .ZN(new_n950));
  INV_X1    g0750(.A(new_n726), .ZN(new_n951));
  OAI221_X1 g0751(.A(new_n732), .B1(new_n210), .B2(new_n574), .C1(new_n243), .C2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n950), .A2(new_n734), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n731), .B2(new_n891), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n932), .A2(new_n955), .ZN(G387));
  AOI21_X1  g0756(.A(new_n637), .B1(new_n677), .B2(new_n925), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n677), .B2(new_n925), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n698), .A2(G50), .ZN(new_n959));
  INV_X1    g0759(.A(G150), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n959), .B1(new_n700), .B2(new_n355), .C1(new_n960), .C2(new_n682), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n693), .A2(new_n215), .B1(new_n703), .B2(new_n203), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n399), .B1(new_n776), .B2(new_n686), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n574), .A2(new_n690), .B1(new_n289), .B2(new_n706), .ZN(new_n964));
  NOR4_X1   g0764(.A1(new_n961), .A2(new_n962), .A3(new_n963), .A4(new_n964), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT111), .Z(new_n966));
  AOI22_X1  g0766(.A1(new_n687), .A2(G322), .B1(new_n759), .B2(G303), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n967), .B1(new_n704), .B2(new_n706), .C1(new_n697), .C2(new_n942), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT48), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n969), .B1(new_n502), .B2(new_n693), .C1(new_n690), .C2(new_n762), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT49), .Z(new_n971));
  AOI21_X1  g0771(.A(new_n399), .B1(new_n683), .B2(G326), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n451), .B2(new_n700), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n966), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n721), .ZN(new_n975));
  INV_X1    g0775(.A(new_n325), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n201), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT50), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n203), .A2(new_n757), .ZN(new_n979));
  NOR4_X1   g0779(.A1(new_n978), .A2(G45), .A3(new_n979), .A4(new_n639), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n951), .B1(new_n239), .B2(G45), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(new_n639), .B2(new_n723), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n980), .A2(new_n982), .B1(G107), .B2(new_n210), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n732), .ZN(new_n984));
  INV_X1    g0784(.A(new_n731), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n975), .B(new_n984), .C1(new_n628), .C2(new_n985), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n958), .B1(new_n735), .B2(new_n986), .C1(new_n929), .C2(new_n925), .ZN(G393));
  OR2_X1    g0787(.A1(new_n916), .A2(new_n917), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n988), .A2(new_n929), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n901), .A2(new_n731), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n686), .A2(new_n707), .B1(new_n697), .B2(new_n704), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT52), .Z(new_n992));
  AOI21_X1  g0792(.A(new_n257), .B1(new_n694), .B2(new_n761), .ZN(new_n993));
  INV_X1    g0793(.A(G322), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n993), .B1(new_n700), .B2(new_n335), .C1(new_n994), .C2(new_n682), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT114), .Z(new_n996));
  AOI211_X1 g0796(.A(new_n992), .B(new_n996), .C1(G116), .C2(new_n712), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n997), .B1(new_n502), .B2(new_n703), .C1(new_n471), .C2(new_n706), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n690), .A2(new_n757), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(new_n976), .B2(new_n759), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n201), .B2(new_n706), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n1002), .A2(KEYINPUT113), .B1(G87), .B2(new_n701), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n686), .A2(new_n960), .B1(new_n697), .B2(new_n776), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT51), .Z(new_n1005));
  INV_X1    g0805(.A(G143), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n682), .A2(new_n1006), .B1(new_n203), .B2(new_n693), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n410), .B(new_n1005), .C1(KEYINPUT112), .C2(new_n1007), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n1003), .A2(new_n1008), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(KEYINPUT112), .B2(new_n1007), .C1(KEYINPUT113), .C2(new_n1002), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n998), .A2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT115), .Z(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n721), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n732), .B1(new_n355), .B2(new_n210), .C1(new_n250), .C2(new_n951), .ZN(new_n1014));
  AND3_X1   g0814(.A1(new_n1013), .A2(new_n734), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n989), .B1(new_n990), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n988), .B1(new_n677), .B2(new_n925), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n927), .A2(new_n1017), .A3(new_n636), .ZN(new_n1018));
  AOI21_X1  g0818(.A(KEYINPUT116), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1016), .A2(KEYINPUT116), .A3(new_n1018), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(G390));
  INV_X1    g0822(.A(new_n783), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n821), .A2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n749), .A2(new_n352), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n747), .B1(new_n655), .B2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1024), .B1(new_n1026), .B2(new_n835), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n819), .A2(KEYINPUT103), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n859), .A2(new_n811), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n823), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n836), .A2(new_n1023), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1027), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n851), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(G330), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n795), .B1(new_n799), .B2(new_n800), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n809), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n811), .B1(new_n1037), .B2(new_n801), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1029), .B1(new_n1038), .B2(new_n822), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n823), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1039), .A2(new_n1040), .A3(new_n1031), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1027), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n675), .A2(G330), .A3(new_n848), .A4(new_n835), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  NOR3_X1   g0845(.A1(new_n1035), .A2(new_n1045), .A3(new_n929), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1030), .A2(new_n729), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n703), .A2(new_n355), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n683), .A2(G294), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n257), .B(new_n999), .C1(G107), .C2(new_n773), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G283), .A2(new_n687), .B1(new_n694), .B2(G87), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1049), .A2(new_n772), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1048), .B(new_n1052), .C1(G116), .C2(new_n698), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n693), .A2(new_n960), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT53), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(G132), .A2(new_n698), .B1(new_n773), .B2(G137), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n687), .A2(G128), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1055), .A2(new_n257), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(G125), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n682), .A2(new_n1059), .B1(new_n700), .B2(new_n201), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n690), .A2(new_n776), .ZN(new_n1061));
  XOR2_X1   g0861(.A(KEYINPUT54), .B(G143), .Z(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1063), .A2(new_n703), .ZN(new_n1064));
  NOR4_X1   g0864(.A1(new_n1058), .A2(new_n1060), .A3(new_n1061), .A4(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n721), .B1(new_n1053), .B2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1047), .A2(new_n734), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n289), .B2(new_n756), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1046), .A2(new_n1068), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n353), .A2(G330), .A3(new_n448), .A4(new_n845), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1070), .B(new_n841), .C1(new_n656), .C2(new_n449), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n835), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n676), .B2(new_n750), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n1034), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n827), .ZN(new_n1075));
  AND2_X1   g0875(.A1(new_n654), .A2(new_n630), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1025), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n746), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n751), .A2(G330), .A3(new_n845), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n1072), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1078), .A2(new_n1080), .A3(new_n1043), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1071), .B1(new_n1075), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n1035), .B2(new_n1045), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1044), .B(new_n1082), .C1(new_n1032), .C2(new_n1034), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1084), .A2(new_n636), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1069), .A2(new_n1086), .ZN(G378));
  INV_X1    g0887(.A(new_n1071), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT119), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n1037), .A2(new_n801), .B1(new_n852), .B2(new_n851), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n821), .A2(new_n1033), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n1091), .A2(new_n855), .B1(new_n1092), .B2(KEYINPUT40), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1090), .B1(new_n1093), .B2(new_n622), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1094), .A2(new_n824), .A3(new_n839), .ZN(new_n1095));
  AOI21_X1  g0895(.A(KEYINPUT119), .B1(new_n861), .B2(G330), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1023), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1096), .B1(new_n1097), .B2(new_n838), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n861), .A2(KEYINPUT119), .A3(G330), .ZN(new_n1100));
  XOR2_X1   g0900(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1101));
  OR3_X1    g0901(.A1(new_n320), .A2(new_n347), .A3(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1101), .B1(new_n320), .B2(new_n347), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n302), .A2(new_n615), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1104), .B(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1100), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1099), .A2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1095), .A2(new_n1098), .A3(new_n1100), .A4(new_n1107), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1089), .A2(new_n1109), .A3(KEYINPUT57), .A4(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n636), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT120), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1089), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT57), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1111), .A2(KEYINPUT120), .A3(new_n636), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1114), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1109), .A2(new_n930), .A3(new_n1110), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n735), .B1(new_n1107), .B2(new_n729), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n756), .A2(new_n201), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n701), .A2(G58), .B1(new_n322), .B2(new_n759), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n355), .B2(new_n706), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(G283), .B2(new_n683), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n203), .B2(new_n690), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n410), .B1(new_n451), .B2(new_n686), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n335), .A2(new_n697), .B1(new_n693), .B2(new_n215), .ZN(new_n1128));
  NOR4_X1   g0928(.A1(new_n1126), .A2(G41), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  XOR2_X1   g0929(.A(new_n1129), .B(KEYINPUT58), .Z(new_n1130));
  AOI21_X1  g0930(.A(new_n259), .B1(new_n396), .B2(new_n398), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n201), .B1(new_n1131), .B2(G41), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n712), .A2(G150), .B1(new_n698), .B2(G128), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(G125), .A2(new_n687), .B1(new_n773), .B2(G132), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n1135), .B1(new_n775), .B2(new_n703), .C1(new_n693), .C2(new_n1063), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT59), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(G33), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1140));
  AOI21_X1  g0940(.A(G41), .B1(new_n683), .B2(G124), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1140), .B(new_n1141), .C1(new_n776), .C2(new_n700), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1130), .B(new_n1132), .C1(new_n1139), .C2(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT117), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n721), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT118), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1121), .A2(new_n1122), .A3(new_n1146), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n1120), .A2(new_n1147), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1119), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(G375));
  NAND3_X1  g0950(.A1(new_n1075), .A2(new_n1071), .A3(new_n1081), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n906), .B(KEYINPUT121), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1083), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n263), .B1(new_n700), .B2(new_n757), .ZN(new_n1154));
  XOR2_X1   g0954(.A(new_n1154), .B(KEYINPUT122), .Z(new_n1155));
  NAND2_X1  g0955(.A1(new_n698), .A2(G283), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n687), .A2(G294), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n682), .A2(new_n471), .B1(new_n355), .B2(new_n693), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n574), .A2(new_n690), .B1(new_n335), .B2(new_n703), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .A4(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(G116), .B2(new_n773), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n410), .B1(new_n701), .B2(G58), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1163), .A2(KEYINPUT123), .B1(G159), .B2(new_n694), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(G137), .A2(new_n698), .B1(new_n759), .B2(G150), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1164), .B(new_n1165), .C1(new_n769), .C2(new_n686), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n690), .A2(new_n201), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1063), .A2(new_n706), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n683), .A2(G128), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n1163), .B2(KEYINPUT123), .ZN(new_n1170));
  NOR4_X1   g0970(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .A4(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n721), .B1(new_n1162), .B2(new_n1171), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n734), .B(new_n1172), .C1(new_n835), .C2(new_n730), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(new_n203), .B2(new_n756), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1075), .A2(new_n1081), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1174), .B1(new_n1175), .B2(new_n930), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1153), .A2(new_n1176), .ZN(G381));
  AND3_X1   g0977(.A1(new_n1069), .A2(new_n1086), .A3(KEYINPUT125), .ZN(new_n1178));
  AOI21_X1  g0978(.A(KEYINPUT125), .B1(new_n1069), .B2(new_n1086), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(G375), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1021), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1182), .A2(new_n1019), .ZN(new_n1183));
  NOR3_X1   g0983(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1184), .B(KEYINPUT124), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(G387), .A2(G381), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1181), .A2(new_n1183), .A3(new_n1185), .A4(new_n1186), .ZN(G407));
  INV_X1    g0987(.A(G213), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(new_n1181), .B2(new_n616), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(G407), .ZN(G409));
  NAND2_X1  g0990(.A1(G387), .A2(new_n1183), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n954), .B1(new_n905), .B2(new_n931), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(G390), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT126), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(G393), .B(new_n744), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1191), .A2(new_n1193), .A3(new_n1194), .A4(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(KEYINPUT126), .B1(new_n1192), .B2(G390), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n1199), .A2(new_n1196), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1188), .A2(G343), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT60), .ZN(new_n1203));
  OR2_X1    g1003(.A1(new_n1151), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1151), .A2(new_n1203), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1204), .A2(new_n636), .A3(new_n1083), .A4(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1206), .A2(G384), .A3(new_n1176), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(G384), .B1(new_n1206), .B2(new_n1176), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1119), .A2(G378), .A3(new_n1148), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1152), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1148), .B1(new_n1115), .B2(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1202), .B(new_n1211), .C1(new_n1212), .C2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT62), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1202), .B1(new_n1212), .B2(new_n1215), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1202), .A2(G2897), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1210), .B(new_n1219), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n1216), .A2(new_n1217), .B1(new_n1218), .B2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1212), .A2(new_n1215), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1202), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1222), .A2(new_n1217), .A3(new_n1223), .A4(new_n1210), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT61), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1201), .B1(new_n1221), .B2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(KEYINPUT63), .B1(new_n1218), .B2(new_n1220), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1218), .A2(new_n1210), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1201), .A2(KEYINPUT61), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1216), .A2(KEYINPUT63), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1227), .A2(new_n1233), .ZN(G405));
  INV_X1    g1034(.A(KEYINPUT127), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1199), .A2(new_n1196), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1239), .A2(KEYINPUT127), .A3(new_n1197), .ZN(new_n1240));
  AND3_X1   g1040(.A1(new_n1236), .A2(new_n1211), .A3(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1211), .B1(new_n1236), .B2(new_n1240), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1212), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1149), .A2(new_n1180), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n1241), .A2(new_n1242), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1236), .A2(new_n1240), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n1210), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1244), .A2(new_n1243), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1236), .A2(new_n1240), .A3(new_n1211), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1247), .A2(new_n1248), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1245), .A2(new_n1250), .ZN(G402));
endmodule


