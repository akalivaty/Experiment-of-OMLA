

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584;

  INV_X1 U320 ( .A(KEYINPUT11), .ZN(n383) );
  XNOR2_X1 U321 ( .A(n349), .B(n348), .ZN(n571) );
  XNOR2_X1 U322 ( .A(n347), .B(n346), .ZN(n348) );
  INV_X1 U323 ( .A(KEYINPUT45), .ZN(n393) );
  XNOR2_X1 U324 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U325 ( .A(n396), .B(n395), .ZN(n398) );
  XOR2_X1 U326 ( .A(G85GAT), .B(G92GAT), .Z(n372) );
  XNOR2_X1 U327 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U328 ( .A(n339), .B(n338), .ZN(n341) );
  XNOR2_X1 U329 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U330 ( .A(KEYINPUT55), .B(KEYINPUT119), .ZN(n438) );
  XNOR2_X1 U331 ( .A(n386), .B(n385), .ZN(n389) );
  XNOR2_X1 U332 ( .A(KEYINPUT96), .B(KEYINPUT36), .ZN(n392) );
  XNOR2_X1 U333 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U334 ( .A(n450), .B(n392), .ZN(n582) );
  INV_X1 U335 ( .A(G134GAT), .ZN(n451) );
  XNOR2_X1 U336 ( .A(n441), .B(G176GAT), .ZN(n442) );
  XNOR2_X1 U337 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U338 ( .A(n443), .B(n442), .ZN(G1349GAT) );
  XOR2_X1 U339 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n291) );
  XOR2_X1 U340 ( .A(G113GAT), .B(G15GAT), .Z(n325) );
  NAND2_X1 U341 ( .A1(G227GAT), .A2(G233GAT), .ZN(n288) );
  XOR2_X1 U342 ( .A(G43GAT), .B(G134GAT), .Z(n382) );
  XNOR2_X1 U343 ( .A(n288), .B(n382), .ZN(n289) );
  XNOR2_X1 U344 ( .A(n325), .B(n289), .ZN(n290) );
  XNOR2_X1 U345 ( .A(n291), .B(n290), .ZN(n294) );
  XOR2_X1 U346 ( .A(G127GAT), .B(KEYINPUT0), .Z(n293) );
  XNOR2_X1 U347 ( .A(KEYINPUT80), .B(KEYINPUT81), .ZN(n292) );
  XNOR2_X1 U348 ( .A(n293), .B(n292), .ZN(n434) );
  XOR2_X1 U349 ( .A(n294), .B(n434), .Z(n302) );
  XOR2_X1 U350 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n296) );
  XNOR2_X1 U351 ( .A(G190GAT), .B(KEYINPUT19), .ZN(n295) );
  XNOR2_X1 U352 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U353 ( .A(n297), .B(G183GAT), .Z(n299) );
  XNOR2_X1 U354 ( .A(G169GAT), .B(G176GAT), .ZN(n298) );
  XNOR2_X1 U355 ( .A(n299), .B(n298), .ZN(n312) );
  XNOR2_X1 U356 ( .A(G99GAT), .B(G71GAT), .ZN(n300) );
  XNOR2_X1 U357 ( .A(n300), .B(G120GAT), .ZN(n345) );
  XNOR2_X1 U358 ( .A(n312), .B(n345), .ZN(n301) );
  XNOR2_X1 U359 ( .A(n302), .B(n301), .ZN(n458) );
  XOR2_X1 U360 ( .A(G204GAT), .B(G64GAT), .Z(n331) );
  XOR2_X1 U361 ( .A(n331), .B(G92GAT), .Z(n307) );
  XOR2_X1 U362 ( .A(KEYINPUT84), .B(G218GAT), .Z(n304) );
  XNOR2_X1 U363 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n303) );
  XNOR2_X1 U364 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U365 ( .A(G197GAT), .B(n305), .Z(n417) );
  XNOR2_X1 U366 ( .A(G36GAT), .B(n417), .ZN(n306) );
  XNOR2_X1 U367 ( .A(n307), .B(n306), .ZN(n311) );
  XOR2_X1 U368 ( .A(KEYINPUT87), .B(KEYINPUT88), .Z(n309) );
  NAND2_X1 U369 ( .A1(G226GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U370 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U371 ( .A(n311), .B(n310), .Z(n314) );
  XNOR2_X1 U372 ( .A(G8GAT), .B(n312), .ZN(n313) );
  XNOR2_X1 U373 ( .A(n314), .B(n313), .ZN(n459) );
  XOR2_X1 U374 ( .A(KEYINPUT66), .B(G197GAT), .Z(n316) );
  XNOR2_X1 U375 ( .A(G169GAT), .B(G141GAT), .ZN(n315) );
  XNOR2_X1 U376 ( .A(n316), .B(n315), .ZN(n330) );
  XOR2_X1 U377 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n318) );
  NAND2_X1 U378 ( .A1(G229GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U379 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U380 ( .A(n319), .B(KEYINPUT67), .Z(n324) );
  XOR2_X1 U381 ( .A(G29GAT), .B(G36GAT), .Z(n321) );
  XNOR2_X1 U382 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n320) );
  XNOR2_X1 U383 ( .A(n321), .B(n320), .ZN(n387) );
  XNOR2_X1 U384 ( .A(G22GAT), .B(G1GAT), .ZN(n322) );
  XNOR2_X1 U385 ( .A(n322), .B(G8GAT), .ZN(n354) );
  XNOR2_X1 U386 ( .A(n387), .B(n354), .ZN(n323) );
  XNOR2_X1 U387 ( .A(n324), .B(n323), .ZN(n326) );
  XOR2_X1 U388 ( .A(n326), .B(n325), .Z(n328) );
  XNOR2_X1 U389 ( .A(G43GAT), .B(G50GAT), .ZN(n327) );
  XNOR2_X1 U390 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U391 ( .A(n330), .B(n329), .Z(n503) );
  INV_X1 U392 ( .A(n503), .ZN(n568) );
  XOR2_X1 U393 ( .A(KEYINPUT32), .B(n372), .Z(n333) );
  XNOR2_X1 U394 ( .A(G176GAT), .B(n331), .ZN(n332) );
  XNOR2_X1 U395 ( .A(n333), .B(n332), .ZN(n339) );
  XOR2_X1 U396 ( .A(KEYINPUT72), .B(KEYINPUT33), .Z(n335) );
  XNOR2_X1 U397 ( .A(KEYINPUT71), .B(KEYINPUT31), .ZN(n334) );
  XOR2_X1 U398 ( .A(n335), .B(n334), .Z(n337) );
  NAND2_X1 U399 ( .A1(G230GAT), .A2(G233GAT), .ZN(n336) );
  INV_X1 U400 ( .A(KEYINPUT70), .ZN(n340) );
  XNOR2_X1 U401 ( .A(n341), .B(n340), .ZN(n349) );
  XNOR2_X1 U402 ( .A(G106GAT), .B(G78GAT), .ZN(n342) );
  XNOR2_X1 U403 ( .A(n342), .B(G148GAT), .ZN(n409) );
  XOR2_X1 U404 ( .A(KEYINPUT13), .B(KEYINPUT68), .Z(n344) );
  XNOR2_X1 U405 ( .A(G57GAT), .B(KEYINPUT69), .ZN(n343) );
  XNOR2_X1 U406 ( .A(n344), .B(n343), .ZN(n353) );
  XNOR2_X1 U407 ( .A(n409), .B(n353), .ZN(n347) );
  XNOR2_X1 U408 ( .A(n345), .B(KEYINPUT73), .ZN(n346) );
  XOR2_X1 U409 ( .A(n571), .B(KEYINPUT41), .Z(n546) );
  AND2_X1 U410 ( .A1(n568), .A2(n546), .ZN(n350) );
  XNOR2_X1 U411 ( .A(n350), .B(KEYINPUT46), .ZN(n370) );
  XOR2_X1 U412 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n352) );
  XNOR2_X1 U413 ( .A(KEYINPUT12), .B(KEYINPUT14), .ZN(n351) );
  XNOR2_X1 U414 ( .A(n352), .B(n351), .ZN(n369) );
  XNOR2_X1 U415 ( .A(n354), .B(n353), .ZN(n367) );
  XOR2_X1 U416 ( .A(G127GAT), .B(G71GAT), .Z(n356) );
  XNOR2_X1 U417 ( .A(G15GAT), .B(G183GAT), .ZN(n355) );
  XNOR2_X1 U418 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U419 ( .A(G64GAT), .B(G155GAT), .Z(n358) );
  XNOR2_X1 U420 ( .A(G211GAT), .B(G78GAT), .ZN(n357) );
  XNOR2_X1 U421 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U422 ( .A(n360), .B(n359), .Z(n365) );
  XOR2_X1 U423 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n362) );
  NAND2_X1 U424 ( .A1(G231GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U425 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U426 ( .A(KEYINPUT15), .B(n363), .ZN(n364) );
  XNOR2_X1 U427 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U428 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U429 ( .A(n369), .B(n368), .ZN(n575) );
  NOR2_X1 U430 ( .A1(n370), .A2(n575), .ZN(n371) );
  XNOR2_X1 U431 ( .A(n371), .B(KEYINPUT108), .ZN(n390) );
  XOR2_X1 U432 ( .A(G50GAT), .B(G162GAT), .Z(n413) );
  XOR2_X1 U433 ( .A(n372), .B(n413), .Z(n374) );
  NAND2_X1 U434 ( .A1(G232GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U435 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U436 ( .A(KEYINPUT10), .B(KEYINPUT74), .Z(n376) );
  XNOR2_X1 U437 ( .A(G99GAT), .B(G106GAT), .ZN(n375) );
  XNOR2_X1 U438 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U439 ( .A(n378), .B(n377), .Z(n386) );
  XOR2_X1 U440 ( .A(KEYINPUT9), .B(KEYINPUT65), .Z(n380) );
  XNOR2_X1 U441 ( .A(G190GAT), .B(G218GAT), .ZN(n379) );
  XNOR2_X1 U442 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U443 ( .A(n382), .B(n381), .ZN(n384) );
  XNOR2_X1 U444 ( .A(n387), .B(KEYINPUT75), .ZN(n388) );
  XNOR2_X1 U445 ( .A(n389), .B(n388), .ZN(n450) );
  NAND2_X1 U446 ( .A1(n390), .A2(n450), .ZN(n391) );
  XNOR2_X1 U447 ( .A(n391), .B(KEYINPUT47), .ZN(n401) );
  INV_X1 U448 ( .A(n575), .ZN(n487) );
  NOR2_X1 U449 ( .A1(n582), .A2(n487), .ZN(n396) );
  XNOR2_X1 U450 ( .A(KEYINPUT64), .B(KEYINPUT109), .ZN(n394) );
  INV_X1 U451 ( .A(n571), .ZN(n397) );
  NAND2_X1 U452 ( .A1(n398), .A2(n397), .ZN(n399) );
  NOR2_X1 U453 ( .A1(n568), .A2(n399), .ZN(n400) );
  NOR2_X1 U454 ( .A1(n401), .A2(n400), .ZN(n402) );
  XNOR2_X1 U455 ( .A(n402), .B(KEYINPUT48), .ZN(n445) );
  NOR2_X1 U456 ( .A1(n459), .A2(n445), .ZN(n403) );
  XNOR2_X1 U457 ( .A(n403), .B(KEYINPUT54), .ZN(n564) );
  XOR2_X1 U458 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n405) );
  NAND2_X1 U459 ( .A1(G228GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U460 ( .A(n405), .B(n404), .ZN(n408) );
  XOR2_X1 U461 ( .A(G155GAT), .B(KEYINPUT2), .Z(n407) );
  XNOR2_X1 U462 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n406) );
  XNOR2_X1 U463 ( .A(n407), .B(n406), .ZN(n433) );
  XOR2_X1 U464 ( .A(n408), .B(n433), .Z(n411) );
  XNOR2_X1 U465 ( .A(G22GAT), .B(n409), .ZN(n410) );
  XNOR2_X1 U466 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U467 ( .A(n412), .B(KEYINPUT24), .Z(n415) );
  XNOR2_X1 U468 ( .A(n413), .B(G204GAT), .ZN(n414) );
  XNOR2_X1 U469 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U470 ( .A(n417), .B(n416), .ZN(n462) );
  XOR2_X1 U471 ( .A(G85GAT), .B(G162GAT), .Z(n419) );
  XNOR2_X1 U472 ( .A(G29GAT), .B(G134GAT), .ZN(n418) );
  XNOR2_X1 U473 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U474 ( .A(KEYINPUT1), .B(G148GAT), .Z(n421) );
  XNOR2_X1 U475 ( .A(G113GAT), .B(G120GAT), .ZN(n420) );
  XNOR2_X1 U476 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U477 ( .A(n423), .B(n422), .Z(n428) );
  XOR2_X1 U478 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n425) );
  NAND2_X1 U479 ( .A1(G225GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U480 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U481 ( .A(KEYINPUT86), .B(n426), .ZN(n427) );
  XNOR2_X1 U482 ( .A(n428), .B(n427), .ZN(n432) );
  XOR2_X1 U483 ( .A(KEYINPUT6), .B(KEYINPUT85), .Z(n430) );
  XNOR2_X1 U484 ( .A(G1GAT), .B(G57GAT), .ZN(n429) );
  XNOR2_X1 U485 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U486 ( .A(n432), .B(n431), .Z(n436) );
  XNOR2_X1 U487 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U488 ( .A(n436), .B(n435), .ZN(n517) );
  INV_X1 U489 ( .A(n517), .ZN(n563) );
  AND2_X1 U490 ( .A1(n462), .A2(n563), .ZN(n437) );
  NAND2_X1 U491 ( .A1(n564), .A2(n437), .ZN(n439) );
  NOR2_X1 U492 ( .A1(n458), .A2(n440), .ZN(n557) );
  NAND2_X1 U493 ( .A1(n557), .A2(n546), .ZN(n443) );
  XOR2_X1 U494 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n441) );
  XNOR2_X1 U495 ( .A(KEYINPUT28), .B(n462), .ZN(n482) );
  XOR2_X1 U496 ( .A(n459), .B(KEYINPUT89), .Z(n444) );
  XNOR2_X1 U497 ( .A(KEYINPUT27), .B(n444), .ZN(n465) );
  NOR2_X1 U498 ( .A1(n445), .A2(n465), .ZN(n446) );
  NAND2_X1 U499 ( .A1(n517), .A2(n446), .ZN(n447) );
  XNOR2_X1 U500 ( .A(KEYINPUT110), .B(n447), .ZN(n541) );
  NOR2_X1 U501 ( .A1(n458), .A2(n541), .ZN(n448) );
  NAND2_X1 U502 ( .A1(n482), .A2(n448), .ZN(n449) );
  XNOR2_X1 U503 ( .A(KEYINPUT111), .B(n449), .ZN(n535) );
  INV_X1 U504 ( .A(n450), .ZN(n556) );
  NAND2_X1 U505 ( .A1(n535), .A2(n556), .ZN(n454) );
  XOR2_X1 U506 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n452) );
  XNOR2_X1 U507 ( .A(n454), .B(n453), .ZN(G1343GAT) );
  NOR2_X1 U508 ( .A1(n503), .A2(n571), .ZN(n489) );
  XNOR2_X1 U509 ( .A(KEYINPUT83), .B(n458), .ZN(n455) );
  NOR2_X1 U510 ( .A1(n465), .A2(n455), .ZN(n456) );
  NAND2_X1 U511 ( .A1(n482), .A2(n456), .ZN(n457) );
  NAND2_X1 U512 ( .A1(n457), .A2(n517), .ZN(n470) );
  INV_X1 U513 ( .A(n458), .ZN(n523) );
  INV_X1 U514 ( .A(n459), .ZN(n521) );
  NAND2_X1 U515 ( .A1(n523), .A2(n521), .ZN(n460) );
  NAND2_X1 U516 ( .A1(n462), .A2(n460), .ZN(n461) );
  XOR2_X1 U517 ( .A(KEYINPUT25), .B(n461), .Z(n468) );
  NOR2_X1 U518 ( .A1(n523), .A2(n462), .ZN(n464) );
  XNOR2_X1 U519 ( .A(KEYINPUT26), .B(KEYINPUT90), .ZN(n463) );
  XNOR2_X1 U520 ( .A(n464), .B(n463), .ZN(n566) );
  INV_X1 U521 ( .A(n566), .ZN(n540) );
  NOR2_X1 U522 ( .A1(n540), .A2(n465), .ZN(n466) );
  NOR2_X1 U523 ( .A1(n517), .A2(n466), .ZN(n467) );
  NAND2_X1 U524 ( .A1(n468), .A2(n467), .ZN(n469) );
  NAND2_X1 U525 ( .A1(n470), .A2(n469), .ZN(n471) );
  XOR2_X1 U526 ( .A(KEYINPUT91), .B(n471), .Z(n485) );
  NOR2_X1 U527 ( .A1(n487), .A2(n556), .ZN(n472) );
  XOR2_X1 U528 ( .A(KEYINPUT16), .B(n472), .Z(n473) );
  NOR2_X1 U529 ( .A1(n485), .A2(n473), .ZN(n505) );
  NAND2_X1 U530 ( .A1(n489), .A2(n505), .ZN(n474) );
  XOR2_X1 U531 ( .A(KEYINPUT92), .B(n474), .Z(n483) );
  NAND2_X1 U532 ( .A1(n483), .A2(n517), .ZN(n475) );
  XNOR2_X1 U533 ( .A(n475), .B(KEYINPUT34), .ZN(n476) );
  XNOR2_X1 U534 ( .A(G1GAT), .B(n476), .ZN(G1324GAT) );
  XOR2_X1 U535 ( .A(G8GAT), .B(KEYINPUT93), .Z(n478) );
  NAND2_X1 U536 ( .A1(n483), .A2(n521), .ZN(n477) );
  XNOR2_X1 U537 ( .A(n478), .B(n477), .ZN(G1325GAT) );
  XOR2_X1 U538 ( .A(KEYINPUT94), .B(KEYINPUT35), .Z(n480) );
  NAND2_X1 U539 ( .A1(n483), .A2(n523), .ZN(n479) );
  XNOR2_X1 U540 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U541 ( .A(G15GAT), .B(n481), .ZN(G1326GAT) );
  INV_X1 U542 ( .A(n482), .ZN(n525) );
  NAND2_X1 U543 ( .A1(n483), .A2(n525), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n484), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U545 ( .A1(n582), .A2(n485), .ZN(n486) );
  NAND2_X1 U546 ( .A1(n487), .A2(n486), .ZN(n488) );
  XNOR2_X1 U547 ( .A(KEYINPUT37), .B(n488), .ZN(n515) );
  NAND2_X1 U548 ( .A1(n515), .A2(n489), .ZN(n490) );
  XNOR2_X1 U549 ( .A(n490), .B(KEYINPUT97), .ZN(n491) );
  XNOR2_X1 U550 ( .A(KEYINPUT38), .B(n491), .ZN(n499) );
  NAND2_X1 U551 ( .A1(n499), .A2(n517), .ZN(n494) );
  XNOR2_X1 U552 ( .A(G29GAT), .B(KEYINPUT95), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n492), .B(KEYINPUT39), .ZN(n493) );
  XNOR2_X1 U554 ( .A(n494), .B(n493), .ZN(G1328GAT) );
  NAND2_X1 U555 ( .A1(n499), .A2(n521), .ZN(n495) );
  XNOR2_X1 U556 ( .A(n495), .B(KEYINPUT98), .ZN(n496) );
  XNOR2_X1 U557 ( .A(G36GAT), .B(n496), .ZN(G1329GAT) );
  NAND2_X1 U558 ( .A1(n499), .A2(n523), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n497), .B(KEYINPUT40), .ZN(n498) );
  XNOR2_X1 U560 ( .A(G43GAT), .B(n498), .ZN(G1330GAT) );
  NAND2_X1 U561 ( .A1(n525), .A2(n499), .ZN(n500) );
  XNOR2_X1 U562 ( .A(G50GAT), .B(n500), .ZN(G1331GAT) );
  XNOR2_X1 U563 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n501), .B(KEYINPUT102), .ZN(n502) );
  XOR2_X1 U565 ( .A(KEYINPUT99), .B(n502), .Z(n508) );
  NAND2_X1 U566 ( .A1(n546), .A2(n503), .ZN(n504) );
  XOR2_X1 U567 ( .A(n504), .B(KEYINPUT100), .Z(n516) );
  NAND2_X1 U568 ( .A1(n505), .A2(n516), .ZN(n506) );
  XNOR2_X1 U569 ( .A(KEYINPUT101), .B(n506), .ZN(n512) );
  NAND2_X1 U570 ( .A1(n512), .A2(n517), .ZN(n507) );
  XNOR2_X1 U571 ( .A(n508), .B(n507), .ZN(G1332GAT) );
  NAND2_X1 U572 ( .A1(n521), .A2(n512), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n509), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U574 ( .A(G71GAT), .B(KEYINPUT103), .Z(n511) );
  NAND2_X1 U575 ( .A1(n512), .A2(n523), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(G1334GAT) );
  XOR2_X1 U577 ( .A(G78GAT), .B(KEYINPUT43), .Z(n514) );
  NAND2_X1 U578 ( .A1(n512), .A2(n525), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n514), .B(n513), .ZN(G1335GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n519) );
  AND2_X1 U581 ( .A1(n516), .A2(n515), .ZN(n526) );
  NAND2_X1 U582 ( .A1(n526), .A2(n517), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U584 ( .A(G85GAT), .B(n520), .ZN(G1336GAT) );
  NAND2_X1 U585 ( .A1(n521), .A2(n526), .ZN(n522) );
  XNOR2_X1 U586 ( .A(n522), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U587 ( .A1(n523), .A2(n526), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n524), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(KEYINPUT106), .ZN(n530) );
  XOR2_X1 U590 ( .A(KEYINPUT107), .B(KEYINPUT44), .Z(n528) );
  NAND2_X1 U591 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U593 ( .A(n530), .B(n529), .ZN(G1339GAT) );
  NAND2_X1 U594 ( .A1(n568), .A2(n535), .ZN(n531) );
  XNOR2_X1 U595 ( .A(n531), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT112), .B(KEYINPUT49), .Z(n533) );
  NAND2_X1 U597 ( .A1(n535), .A2(n546), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U599 ( .A(G120GAT), .B(n534), .ZN(G1341GAT) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(KEYINPUT113), .ZN(n539) );
  XOR2_X1 U601 ( .A(KEYINPUT114), .B(KEYINPUT50), .Z(n537) );
  NAND2_X1 U602 ( .A1(n535), .A2(n575), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(G1342GAT) );
  NOR2_X1 U605 ( .A1(n541), .A2(n540), .ZN(n551) );
  NAND2_X1 U606 ( .A1(n551), .A2(n568), .ZN(n542) );
  XNOR2_X1 U607 ( .A(G141GAT), .B(n542), .ZN(G1344GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT53), .B(KEYINPUT117), .Z(n544) );
  XNOR2_X1 U609 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U611 ( .A(KEYINPUT116), .B(n545), .Z(n548) );
  NAND2_X1 U612 ( .A1(n551), .A2(n546), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(G1345GAT) );
  NAND2_X1 U614 ( .A1(n575), .A2(n551), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n549), .B(KEYINPUT118), .ZN(n550) );
  XNOR2_X1 U616 ( .A(G155GAT), .B(n550), .ZN(G1346GAT) );
  NAND2_X1 U617 ( .A1(n556), .A2(n551), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n552), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U619 ( .A(G169GAT), .B(KEYINPUT120), .ZN(n554) );
  NAND2_X1 U620 ( .A1(n557), .A2(n568), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(G1348GAT) );
  NAND2_X1 U622 ( .A1(n575), .A2(n557), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n555), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U624 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n559) );
  NAND2_X1 U625 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1351GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n561) );
  XNOR2_X1 U628 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n560) );
  XNOR2_X1 U629 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U630 ( .A(KEYINPUT60), .B(n562), .Z(n570) );
  AND2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n565) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(KEYINPUT121), .ZN(n580) );
  NAND2_X1 U634 ( .A1(n580), .A2(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n573) );
  NAND2_X1 U637 ( .A1(n580), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(G204GAT), .B(n574), .ZN(G1353GAT) );
  XOR2_X1 U640 ( .A(G211GAT), .B(KEYINPUT125), .Z(n577) );
  NAND2_X1 U641 ( .A1(n580), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1354GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n579) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n584) );
  INV_X1 U646 ( .A(n580), .ZN(n581) );
  NOR2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U648 ( .A(n584), .B(n583), .Z(G1355GAT) );
endmodule

