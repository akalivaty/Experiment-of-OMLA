

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603;

  XNOR2_X1 U324 ( .A(n487), .B(KEYINPUT96), .ZN(n498) );
  XOR2_X1 U325 ( .A(n347), .B(n351), .Z(n596) );
  XNOR2_X1 U326 ( .A(n365), .B(n364), .ZN(n368) );
  XNOR2_X1 U327 ( .A(n399), .B(n398), .ZN(n538) );
  XOR2_X1 U328 ( .A(n460), .B(n459), .Z(n553) );
  OR2_X1 U329 ( .A1(n478), .A2(n541), .ZN(n292) );
  OR2_X1 U330 ( .A1(n536), .A2(n486), .ZN(n293) );
  NOR2_X1 U331 ( .A1(n480), .A2(n536), .ZN(n294) );
  XNOR2_X1 U332 ( .A(KEYINPUT22), .B(G204GAT), .ZN(n404) );
  XNOR2_X1 U333 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U334 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U335 ( .A(n389), .B(n388), .ZN(n390) );
  NAND2_X1 U336 ( .A1(n292), .A2(n293), .ZN(n487) );
  XNOR2_X1 U337 ( .A(n340), .B(n339), .ZN(n345) );
  XNOR2_X1 U338 ( .A(n460), .B(n390), .ZN(n391) );
  XNOR2_X1 U339 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U340 ( .A(n372), .B(KEYINPUT36), .ZN(n373) );
  XNOR2_X1 U341 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U342 ( .A(n414), .B(n413), .ZN(n416) );
  XNOR2_X1 U343 ( .A(n579), .B(n373), .ZN(n600) );
  NOR2_X1 U344 ( .A1(n461), .A2(n553), .ZN(n462) );
  INV_X1 U345 ( .A(G211GAT), .ZN(n472) );
  XNOR2_X1 U346 ( .A(n462), .B(KEYINPUT120), .ZN(n588) );
  NOR2_X1 U347 ( .A1(n535), .A2(n534), .ZN(n544) );
  XOR2_X1 U348 ( .A(n480), .B(KEYINPUT28), .Z(n551) );
  XNOR2_X1 U349 ( .A(n472), .B(KEYINPUT126), .ZN(n473) );
  XNOR2_X1 U350 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U351 ( .A(n494), .B(G43GAT), .ZN(n495) );
  XNOR2_X1 U352 ( .A(n474), .B(n473), .ZN(G1354GAT) );
  XNOR2_X1 U353 ( .A(n466), .B(n465), .ZN(G1349GAT) );
  XNOR2_X1 U354 ( .A(n496), .B(n495), .ZN(G1330GAT) );
  XOR2_X1 U355 ( .A(KEYINPUT47), .B(KEYINPUT111), .Z(n371) );
  XOR2_X1 U356 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n296) );
  XNOR2_X1 U357 ( .A(G8GAT), .B(KEYINPUT79), .ZN(n295) );
  XNOR2_X1 U358 ( .A(n296), .B(n295), .ZN(n308) );
  XOR2_X1 U359 ( .A(G211GAT), .B(G71GAT), .Z(n298) );
  XNOR2_X1 U360 ( .A(G183GAT), .B(G127GAT), .ZN(n297) );
  XNOR2_X1 U361 ( .A(n298), .B(n297), .ZN(n306) );
  XOR2_X1 U362 ( .A(KEYINPUT76), .B(KEYINPUT77), .Z(n300) );
  XNOR2_X1 U363 ( .A(KEYINPUT15), .B(KEYINPUT78), .ZN(n299) );
  XNOR2_X1 U364 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U365 ( .A(G64GAT), .B(G155GAT), .Z(n302) );
  XNOR2_X1 U366 ( .A(G22GAT), .B(G78GAT), .ZN(n301) );
  XNOR2_X1 U367 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U368 ( .A(n304), .B(n303), .Z(n305) );
  XNOR2_X1 U369 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U370 ( .A(n308), .B(n307), .ZN(n313) );
  XNOR2_X1 U371 ( .A(G57GAT), .B(KEYINPUT68), .ZN(n309) );
  XNOR2_X1 U372 ( .A(n309), .B(KEYINPUT13), .ZN(n343) );
  XOR2_X1 U373 ( .A(G15GAT), .B(G1GAT), .Z(n320) );
  XOR2_X1 U374 ( .A(n343), .B(n320), .Z(n311) );
  NAND2_X1 U375 ( .A1(G231GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U376 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U377 ( .A(n313), .B(n312), .Z(n575) );
  INV_X1 U378 ( .A(n575), .ZN(n584) );
  XOR2_X1 U379 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n315) );
  XNOR2_X1 U380 ( .A(G43GAT), .B(G29GAT), .ZN(n314) );
  XNOR2_X1 U381 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U382 ( .A(KEYINPUT67), .B(n316), .ZN(n366) );
  XOR2_X1 U383 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n318) );
  XNOR2_X1 U384 ( .A(G113GAT), .B(G197GAT), .ZN(n317) );
  XNOR2_X1 U385 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U386 ( .A(G141GAT), .B(G22GAT), .Z(n410) );
  XNOR2_X1 U387 ( .A(n319), .B(n410), .ZN(n324) );
  XOR2_X1 U388 ( .A(n320), .B(KEYINPUT66), .Z(n322) );
  NAND2_X1 U389 ( .A1(G229GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U390 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U391 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U392 ( .A(G169GAT), .B(G8GAT), .Z(n389) );
  XOR2_X1 U393 ( .A(n325), .B(n389), .Z(n327) );
  XNOR2_X1 U394 ( .A(G50GAT), .B(G36GAT), .ZN(n326) );
  XNOR2_X1 U395 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U396 ( .A(n366), .B(n328), .Z(n581) );
  INV_X1 U397 ( .A(n581), .ZN(n591) );
  XOR2_X1 U398 ( .A(G120GAT), .B(G71GAT), .Z(n446) );
  INV_X1 U399 ( .A(G148GAT), .ZN(n329) );
  NAND2_X1 U400 ( .A1(G78GAT), .A2(n329), .ZN(n332) );
  INV_X1 U401 ( .A(G78GAT), .ZN(n330) );
  NAND2_X1 U402 ( .A1(n330), .A2(G148GAT), .ZN(n331) );
  NAND2_X1 U403 ( .A1(n332), .A2(n331), .ZN(n334) );
  XNOR2_X1 U404 ( .A(G106GAT), .B(KEYINPUT69), .ZN(n333) );
  XNOR2_X1 U405 ( .A(n334), .B(n333), .ZN(n401) );
  XNOR2_X1 U406 ( .A(n401), .B(KEYINPUT71), .ZN(n340) );
  XOR2_X1 U407 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n336) );
  XNOR2_X1 U408 ( .A(KEYINPUT33), .B(KEYINPUT70), .ZN(n335) );
  XNOR2_X1 U409 ( .A(n336), .B(n335), .ZN(n338) );
  AND2_X1 U410 ( .A1(G230GAT), .A2(G233GAT), .ZN(n337) );
  XOR2_X1 U411 ( .A(G64GAT), .B(G92GAT), .Z(n342) );
  XNOR2_X1 U412 ( .A(G176GAT), .B(G204GAT), .ZN(n341) );
  XNOR2_X1 U413 ( .A(n342), .B(n341), .ZN(n397) );
  XOR2_X1 U414 ( .A(n343), .B(n397), .Z(n344) );
  XNOR2_X1 U415 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U416 ( .A(n446), .B(n346), .ZN(n347) );
  XNOR2_X1 U417 ( .A(G99GAT), .B(G85GAT), .ZN(n351) );
  XOR2_X1 U418 ( .A(KEYINPUT41), .B(n596), .Z(n569) );
  NOR2_X1 U419 ( .A1(n591), .A2(n569), .ZN(n348) );
  XNOR2_X1 U420 ( .A(n348), .B(KEYINPUT46), .ZN(n349) );
  NOR2_X1 U421 ( .A1(n584), .A2(n349), .ZN(n369) );
  XOR2_X1 U422 ( .A(G50GAT), .B(G162GAT), .Z(n411) );
  NAND2_X1 U423 ( .A1(G232GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U424 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U425 ( .A(G36GAT), .B(G190GAT), .Z(n392) );
  XNOR2_X1 U426 ( .A(n352), .B(n392), .ZN(n353) );
  XNOR2_X1 U427 ( .A(n411), .B(n353), .ZN(n365) );
  XOR2_X1 U428 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n355) );
  XNOR2_X1 U429 ( .A(G218GAT), .B(KEYINPUT74), .ZN(n354) );
  XNOR2_X1 U430 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U431 ( .A(KEYINPUT64), .B(G92GAT), .Z(n357) );
  XNOR2_X1 U432 ( .A(KEYINPUT65), .B(KEYINPUT10), .ZN(n356) );
  XNOR2_X1 U433 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U434 ( .A(n359), .B(n358), .Z(n363) );
  XOR2_X1 U435 ( .A(KEYINPUT73), .B(KEYINPUT75), .Z(n361) );
  XNOR2_X1 U436 ( .A(G134GAT), .B(G106GAT), .ZN(n360) );
  XNOR2_X1 U437 ( .A(n361), .B(n360), .ZN(n362) );
  INV_X1 U438 ( .A(n366), .ZN(n367) );
  XOR2_X1 U439 ( .A(n368), .B(n367), .Z(n579) );
  NAND2_X1 U440 ( .A1(n369), .A2(n579), .ZN(n370) );
  XNOR2_X1 U441 ( .A(n371), .B(n370), .ZN(n379) );
  INV_X1 U442 ( .A(KEYINPUT101), .ZN(n372) );
  NOR2_X1 U443 ( .A1(n575), .A2(n600), .ZN(n374) );
  XNOR2_X1 U444 ( .A(n374), .B(KEYINPUT45), .ZN(n375) );
  NAND2_X1 U445 ( .A1(n375), .A2(n596), .ZN(n376) );
  NOR2_X1 U446 ( .A1(n581), .A2(n376), .ZN(n377) );
  XNOR2_X1 U447 ( .A(n377), .B(KEYINPUT112), .ZN(n378) );
  NOR2_X1 U448 ( .A1(n379), .A2(n378), .ZN(n380) );
  XNOR2_X1 U449 ( .A(KEYINPUT48), .B(n380), .ZN(n549) );
  XNOR2_X1 U450 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n386) );
  INV_X1 U451 ( .A(KEYINPUT83), .ZN(n381) );
  NAND2_X1 U452 ( .A1(KEYINPUT19), .A2(n381), .ZN(n384) );
  INV_X1 U453 ( .A(KEYINPUT19), .ZN(n382) );
  NAND2_X1 U454 ( .A1(n382), .A2(KEYINPUT83), .ZN(n383) );
  NAND2_X1 U455 ( .A1(n384), .A2(n383), .ZN(n385) );
  XNOR2_X1 U456 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U457 ( .A(KEYINPUT18), .B(n387), .Z(n460) );
  XOR2_X1 U458 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n388) );
  XOR2_X1 U459 ( .A(n392), .B(n391), .Z(n394) );
  NAND2_X1 U460 ( .A1(G226GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U461 ( .A(n394), .B(n393), .ZN(n399) );
  XOR2_X1 U462 ( .A(G211GAT), .B(KEYINPUT21), .Z(n396) );
  XNOR2_X1 U463 ( .A(G197GAT), .B(G218GAT), .ZN(n395) );
  XNOR2_X1 U464 ( .A(n396), .B(n395), .ZN(n405) );
  XNOR2_X1 U465 ( .A(n405), .B(n397), .ZN(n398) );
  INV_X1 U466 ( .A(n538), .ZN(n516) );
  NOR2_X1 U467 ( .A1(n549), .A2(n516), .ZN(n400) );
  XNOR2_X1 U468 ( .A(n400), .B(KEYINPUT54), .ZN(n469) );
  XOR2_X1 U469 ( .A(G155GAT), .B(KEYINPUT2), .Z(n403) );
  XNOR2_X1 U470 ( .A(KEYINPUT84), .B(KEYINPUT3), .ZN(n402) );
  XNOR2_X1 U471 ( .A(n403), .B(n402), .ZN(n427) );
  XNOR2_X1 U472 ( .A(n401), .B(n427), .ZN(n407) );
  XNOR2_X1 U473 ( .A(n407), .B(n406), .ZN(n409) );
  INV_X1 U474 ( .A(KEYINPUT23), .ZN(n408) );
  XNOR2_X1 U475 ( .A(n409), .B(n408), .ZN(n414) );
  XOR2_X1 U476 ( .A(n410), .B(KEYINPUT24), .Z(n412) );
  NAND2_X1 U477 ( .A1(G228GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U478 ( .A(n416), .B(n415), .ZN(n480) );
  XOR2_X1 U479 ( .A(KEYINPUT6), .B(KEYINPUT85), .Z(n418) );
  XNOR2_X1 U480 ( .A(G1GAT), .B(KEYINPUT89), .ZN(n417) );
  XNOR2_X1 U481 ( .A(n418), .B(n417), .ZN(n431) );
  XOR2_X1 U482 ( .A(KEYINPUT1), .B(KEYINPUT90), .Z(n420) );
  XNOR2_X1 U483 ( .A(G57GAT), .B(KEYINPUT88), .ZN(n419) );
  XNOR2_X1 U484 ( .A(n420), .B(n419), .ZN(n424) );
  XOR2_X1 U485 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n422) );
  XNOR2_X1 U486 ( .A(KEYINPUT86), .B(KEYINPUT87), .ZN(n421) );
  XNOR2_X1 U487 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U488 ( .A(n424), .B(n423), .Z(n429) );
  XOR2_X1 U489 ( .A(G127GAT), .B(KEYINPUT0), .Z(n426) );
  XNOR2_X1 U490 ( .A(G113GAT), .B(G134GAT), .ZN(n425) );
  XNOR2_X1 U491 ( .A(n426), .B(n425), .ZN(n454) );
  XNOR2_X1 U492 ( .A(n454), .B(n427), .ZN(n428) );
  XNOR2_X1 U493 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U494 ( .A(n431), .B(n430), .ZN(n439) );
  NAND2_X1 U495 ( .A1(G225GAT), .A2(G233GAT), .ZN(n437) );
  XOR2_X1 U496 ( .A(G148GAT), .B(G162GAT), .Z(n433) );
  XNOR2_X1 U497 ( .A(G141GAT), .B(G120GAT), .ZN(n432) );
  XNOR2_X1 U498 ( .A(n433), .B(n432), .ZN(n435) );
  XOR2_X1 U499 ( .A(G29GAT), .B(G85GAT), .Z(n434) );
  XNOR2_X1 U500 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U501 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U502 ( .A(n439), .B(n438), .Z(n536) );
  AND2_X1 U503 ( .A1(n469), .A2(n294), .ZN(n440) );
  XNOR2_X1 U504 ( .A(n440), .B(KEYINPUT55), .ZN(n461) );
  XOR2_X1 U505 ( .A(KEYINPUT81), .B(G176GAT), .Z(n442) );
  XNOR2_X1 U506 ( .A(G169GAT), .B(G15GAT), .ZN(n441) );
  XOR2_X1 U507 ( .A(n442), .B(n441), .Z(n458) );
  XOR2_X1 U508 ( .A(G190GAT), .B(KEYINPUT20), .Z(n444) );
  XNOR2_X1 U509 ( .A(G43GAT), .B(G99GAT), .ZN(n443) );
  XNOR2_X1 U510 ( .A(n444), .B(n443), .ZN(n447) );
  INV_X1 U511 ( .A(n447), .ZN(n445) );
  NAND2_X1 U512 ( .A1(n446), .A2(n445), .ZN(n450) );
  INV_X1 U513 ( .A(n446), .ZN(n448) );
  NAND2_X1 U514 ( .A1(n448), .A2(n447), .ZN(n449) );
  NAND2_X1 U515 ( .A1(n450), .A2(n449), .ZN(n452) );
  NAND2_X1 U516 ( .A1(G227GAT), .A2(G233GAT), .ZN(n451) );
  XNOR2_X1 U517 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X1 U518 ( .A(n453), .B(KEYINPUT82), .Z(n456) );
  XNOR2_X1 U519 ( .A(n454), .B(KEYINPUT80), .ZN(n455) );
  XNOR2_X1 U520 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U521 ( .A(n458), .B(n457), .ZN(n459) );
  INV_X1 U522 ( .A(n569), .ZN(n556) );
  NAND2_X1 U523 ( .A1(n588), .A2(n556), .ZN(n466) );
  XOR2_X1 U524 ( .A(G176GAT), .B(KEYINPUT122), .Z(n464) );
  XNOR2_X1 U525 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n463) );
  XOR2_X1 U526 ( .A(KEYINPUT26), .B(KEYINPUT95), .Z(n468) );
  NAND2_X1 U527 ( .A1(n480), .A2(n553), .ZN(n467) );
  XOR2_X1 U528 ( .A(n468), .B(n467), .Z(n565) );
  INV_X1 U529 ( .A(n565), .ZN(n483) );
  INV_X1 U530 ( .A(n536), .ZN(n513) );
  NAND2_X1 U531 ( .A1(n469), .A2(n513), .ZN(n470) );
  NOR2_X1 U532 ( .A1(n483), .A2(n470), .ZN(n471) );
  XOR2_X1 U533 ( .A(KEYINPUT124), .B(n471), .Z(n599) );
  NOR2_X1 U534 ( .A1(n575), .A2(n599), .ZN(n474) );
  XOR2_X1 U535 ( .A(KEYINPUT27), .B(n538), .Z(n482) );
  NOR2_X1 U536 ( .A1(n513), .A2(n482), .ZN(n475) );
  XNOR2_X1 U537 ( .A(n475), .B(KEYINPUT93), .ZN(n548) );
  INV_X1 U538 ( .A(n551), .ZN(n528) );
  NOR2_X1 U539 ( .A1(n548), .A2(n528), .ZN(n477) );
  INV_X1 U540 ( .A(KEYINPUT94), .ZN(n476) );
  XNOR2_X1 U541 ( .A(n477), .B(n476), .ZN(n478) );
  INV_X1 U542 ( .A(n553), .ZN(n541) );
  NOR2_X1 U543 ( .A1(n553), .A2(n516), .ZN(n479) );
  NOR2_X1 U544 ( .A1(n480), .A2(n479), .ZN(n481) );
  XOR2_X1 U545 ( .A(KEYINPUT25), .B(n481), .Z(n485) );
  NOR2_X1 U546 ( .A1(n483), .A2(n482), .ZN(n484) );
  NOR2_X1 U547 ( .A1(n485), .A2(n484), .ZN(n486) );
  NOR2_X1 U548 ( .A1(n584), .A2(n600), .ZN(n488) );
  NAND2_X1 U549 ( .A1(n498), .A2(n488), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n489), .B(KEYINPUT102), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n490), .B(KEYINPUT37), .ZN(n533) );
  AND2_X1 U552 ( .A1(n596), .A2(n581), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n491), .B(KEYINPUT72), .ZN(n500) );
  NAND2_X1 U554 ( .A1(n533), .A2(n500), .ZN(n493) );
  XOR2_X1 U555 ( .A(KEYINPUT103), .B(KEYINPUT38), .Z(n492) );
  XNOR2_X1 U556 ( .A(n493), .B(n492), .ZN(n518) );
  NOR2_X1 U557 ( .A1(n553), .A2(n518), .ZN(n496) );
  INV_X1 U558 ( .A(KEYINPUT40), .ZN(n494) );
  INV_X1 U559 ( .A(n579), .ZN(n587) );
  NOR2_X1 U560 ( .A1(n587), .A2(n575), .ZN(n497) );
  XNOR2_X1 U561 ( .A(KEYINPUT16), .B(n497), .ZN(n499) );
  NAND2_X1 U562 ( .A1(n499), .A2(n498), .ZN(n521) );
  INV_X1 U563 ( .A(n521), .ZN(n501) );
  NAND2_X1 U564 ( .A1(n501), .A2(n500), .ZN(n510) );
  NOR2_X1 U565 ( .A1(n513), .A2(n510), .ZN(n503) );
  XNOR2_X1 U566 ( .A(KEYINPUT97), .B(KEYINPUT34), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U568 ( .A(G1GAT), .B(n504), .ZN(G1324GAT) );
  NOR2_X1 U569 ( .A1(n516), .A2(n510), .ZN(n505) );
  XOR2_X1 U570 ( .A(G8GAT), .B(n505), .Z(G1325GAT) );
  NOR2_X1 U571 ( .A1(n510), .A2(n553), .ZN(n509) );
  XOR2_X1 U572 ( .A(KEYINPUT98), .B(KEYINPUT35), .Z(n507) );
  XNOR2_X1 U573 ( .A(G15GAT), .B(KEYINPUT99), .ZN(n506) );
  XNOR2_X1 U574 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n509), .B(n508), .ZN(G1326GAT) );
  NOR2_X1 U576 ( .A1(n551), .A2(n510), .ZN(n511) );
  XOR2_X1 U577 ( .A(KEYINPUT100), .B(n511), .Z(n512) );
  XNOR2_X1 U578 ( .A(G22GAT), .B(n512), .ZN(G1327GAT) );
  NOR2_X1 U579 ( .A1(n518), .A2(n513), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n514), .B(KEYINPUT39), .ZN(n515) );
  XNOR2_X1 U581 ( .A(G29GAT), .B(n515), .ZN(G1328GAT) );
  NOR2_X1 U582 ( .A1(n518), .A2(n516), .ZN(n517) );
  XOR2_X1 U583 ( .A(G36GAT), .B(n517), .Z(G1329GAT) );
  NOR2_X1 U584 ( .A1(n551), .A2(n518), .ZN(n519) );
  XOR2_X1 U585 ( .A(G50GAT), .B(n519), .Z(G1331GAT) );
  NAND2_X1 U586 ( .A1(n556), .A2(n591), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n520), .B(KEYINPUT104), .ZN(n534) );
  NOR2_X1 U588 ( .A1(n534), .A2(n521), .ZN(n522) );
  XOR2_X1 U589 ( .A(KEYINPUT105), .B(n522), .Z(n529) );
  NAND2_X1 U590 ( .A1(n529), .A2(n536), .ZN(n523) );
  XNOR2_X1 U591 ( .A(n523), .B(KEYINPUT42), .ZN(n524) );
  XNOR2_X1 U592 ( .A(G57GAT), .B(n524), .ZN(G1332GAT) );
  NAND2_X1 U593 ( .A1(n538), .A2(n529), .ZN(n525) );
  XNOR2_X1 U594 ( .A(G64GAT), .B(n525), .ZN(G1333GAT) );
  NAND2_X1 U595 ( .A1(n541), .A2(n529), .ZN(n526) );
  XNOR2_X1 U596 ( .A(n526), .B(KEYINPUT106), .ZN(n527) );
  XNOR2_X1 U597 ( .A(G71GAT), .B(n527), .ZN(G1334GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n531) );
  NAND2_X1 U599 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U600 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U601 ( .A(G78GAT), .B(n532), .Z(G1335GAT) );
  INV_X1 U602 ( .A(n533), .ZN(n535) );
  NAND2_X1 U603 ( .A1(n536), .A2(n544), .ZN(n537) );
  XNOR2_X1 U604 ( .A(G85GAT), .B(n537), .ZN(G1336GAT) );
  NAND2_X1 U605 ( .A1(n544), .A2(n538), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n539), .B(KEYINPUT108), .ZN(n540) );
  XNOR2_X1 U607 ( .A(G92GAT), .B(n540), .ZN(G1337GAT) );
  XOR2_X1 U608 ( .A(G99GAT), .B(KEYINPUT109), .Z(n543) );
  NAND2_X1 U609 ( .A1(n544), .A2(n541), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(G1338GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT44), .B(KEYINPUT110), .Z(n546) );
  NAND2_X1 U612 ( .A1(n544), .A2(n528), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U614 ( .A(n547), .B(G106GAT), .Z(G1339GAT) );
  XNOR2_X1 U615 ( .A(G113GAT), .B(KEYINPUT114), .ZN(n555) );
  NOR2_X1 U616 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U617 ( .A(KEYINPUT113), .B(n550), .Z(n566) );
  NAND2_X1 U618 ( .A1(n551), .A2(n566), .ZN(n552) );
  NOR2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n562) );
  NAND2_X1 U620 ( .A1(n562), .A2(n581), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(G1340GAT) );
  XOR2_X1 U622 ( .A(G120GAT), .B(KEYINPUT49), .Z(n558) );
  NAND2_X1 U623 ( .A1(n562), .A2(n556), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1341GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n560) );
  NAND2_X1 U626 ( .A1(n562), .A2(n584), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(G127GAT), .B(n561), .ZN(G1342GAT) );
  XOR2_X1 U629 ( .A(G134GAT), .B(KEYINPUT51), .Z(n564) );
  NAND2_X1 U630 ( .A1(n562), .A2(n587), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(G1343GAT) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n578) );
  NOR2_X1 U633 ( .A1(n591), .A2(n578), .ZN(n567) );
  XOR2_X1 U634 ( .A(G141GAT), .B(n567), .Z(n568) );
  XNOR2_X1 U635 ( .A(KEYINPUT116), .B(n568), .ZN(G1344GAT) );
  NOR2_X1 U636 ( .A1(n569), .A2(n578), .ZN(n574) );
  XOR2_X1 U637 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n571) );
  XNOR2_X1 U638 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n570) );
  XNOR2_X1 U639 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U640 ( .A(KEYINPUT117), .B(n572), .ZN(n573) );
  XNOR2_X1 U641 ( .A(n574), .B(n573), .ZN(G1345GAT) );
  NOR2_X1 U642 ( .A1(n575), .A2(n578), .ZN(n577) );
  XNOR2_X1 U643 ( .A(G155GAT), .B(KEYINPUT119), .ZN(n576) );
  XNOR2_X1 U644 ( .A(n577), .B(n576), .ZN(G1346GAT) );
  NOR2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U646 ( .A(G162GAT), .B(n580), .Z(G1347GAT) );
  XOR2_X1 U647 ( .A(G169GAT), .B(KEYINPUT121), .Z(n583) );
  NAND2_X1 U648 ( .A1(n588), .A2(n581), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(G1348GAT) );
  XOR2_X1 U650 ( .A(G183GAT), .B(KEYINPUT123), .Z(n586) );
  NAND2_X1 U651 ( .A1(n588), .A2(n584), .ZN(n585) );
  XNOR2_X1 U652 ( .A(n586), .B(n585), .ZN(G1350GAT) );
  NAND2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n589), .B(KEYINPUT58), .ZN(n590) );
  XNOR2_X1 U655 ( .A(G190GAT), .B(n590), .ZN(G1351GAT) );
  NOR2_X1 U656 ( .A1(n599), .A2(n591), .ZN(n595) );
  XOR2_X1 U657 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n593) );
  XNOR2_X1 U658 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n592) );
  XNOR2_X1 U659 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U660 ( .A(n595), .B(n594), .ZN(G1352GAT) );
  XNOR2_X1 U661 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n598) );
  NOR2_X1 U662 ( .A1(n596), .A2(n599), .ZN(n597) );
  XNOR2_X1 U663 ( .A(n598), .B(n597), .ZN(G1353GAT) );
  XNOR2_X1 U664 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n602) );
  NOR2_X1 U665 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U666 ( .A(n602), .B(n601), .ZN(n603) );
  XNOR2_X1 U667 ( .A(G218GAT), .B(n603), .ZN(G1355GAT) );
endmodule

