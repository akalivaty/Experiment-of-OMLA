

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X2 U551 ( .A1(G8), .A2(n727), .ZN(n781) );
  NOR2_X1 U552 ( .A1(G2104), .A2(n526), .ZN(n890) );
  NOR2_X1 U553 ( .A1(G2105), .A2(G2104), .ZN(n522) );
  OR2_X1 U554 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U555 ( .A(n716), .B(n715), .ZN(n745) );
  NOR2_X1 U556 ( .A1(n530), .A2(n529), .ZN(G164) );
  XNOR2_X2 U557 ( .A(n525), .B(KEYINPUT65), .ZN(n561) );
  NOR2_X1 U558 ( .A1(n814), .A2(n517), .ZN(n515) );
  XOR2_X1 U559 ( .A(G543), .B(KEYINPUT0), .Z(n516) );
  AND2_X1 U560 ( .A1(n931), .A2(n828), .ZN(n517) );
  XOR2_X1 U561 ( .A(KEYINPUT94), .B(n782), .Z(n518) );
  AND2_X1 U562 ( .A1(n698), .A2(n697), .ZN(n519) );
  NAND2_X1 U563 ( .A1(n924), .A2(n707), .ZN(n520) );
  XNOR2_X1 U564 ( .A(KEYINPUT96), .B(KEYINPUT27), .ZN(n703) );
  XNOR2_X1 U565 ( .A(n704), .B(n703), .ZN(n706) );
  OR2_X1 U566 ( .A1(n710), .A2(n709), .ZN(n714) );
  INV_X1 U567 ( .A(KEYINPUT29), .ZN(n715) );
  INV_X1 U568 ( .A(KEYINPUT101), .ZN(n740) );
  INV_X1 U569 ( .A(KEYINPUT102), .ZN(n761) );
  XNOR2_X1 U570 ( .A(n762), .B(n761), .ZN(n767) );
  INV_X1 U571 ( .A(KEYINPUT17), .ZN(n521) );
  NOR2_X1 U572 ( .A1(G164), .A2(G1384), .ZN(n801) );
  XOR2_X1 U573 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NOR2_X1 U574 ( .A1(n552), .A2(n551), .ZN(G171) );
  XNOR2_X1 U575 ( .A(n522), .B(n521), .ZN(n553) );
  BUF_X1 U576 ( .A(n553), .Z(n885) );
  NAND2_X1 U577 ( .A1(G138), .A2(n885), .ZN(n524) );
  INV_X1 U578 ( .A(G2105), .ZN(n526) );
  AND2_X1 U579 ( .A1(n526), .A2(G2104), .ZN(n886) );
  NAND2_X1 U580 ( .A1(G102), .A2(n886), .ZN(n523) );
  NAND2_X1 U581 ( .A1(n524), .A2(n523), .ZN(n530) );
  NAND2_X1 U582 ( .A1(G2104), .A2(G2105), .ZN(n525) );
  NAND2_X1 U583 ( .A1(G114), .A2(n561), .ZN(n528) );
  NAND2_X1 U584 ( .A1(G126), .A2(n890), .ZN(n527) );
  NAND2_X1 U585 ( .A1(n528), .A2(n527), .ZN(n529) );
  INV_X1 U586 ( .A(G651), .ZN(n537) );
  NOR2_X1 U587 ( .A1(G543), .A2(n537), .ZN(n531) );
  XOR2_X1 U588 ( .A(KEYINPUT1), .B(n531), .Z(n651) );
  NAND2_X1 U589 ( .A1(G63), .A2(n651), .ZN(n533) );
  XNOR2_X1 U590 ( .A(KEYINPUT68), .B(n516), .ZN(n536) );
  NOR2_X1 U591 ( .A1(G651), .A2(n536), .ZN(n589) );
  BUF_X1 U592 ( .A(n589), .Z(n659) );
  NAND2_X1 U593 ( .A1(G51), .A2(n659), .ZN(n532) );
  NAND2_X1 U594 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U595 ( .A(KEYINPUT6), .B(n534), .ZN(n542) );
  NOR2_X1 U596 ( .A1(G651), .A2(G543), .ZN(n652) );
  NAND2_X1 U597 ( .A1(n652), .A2(G89), .ZN(n535) );
  XNOR2_X1 U598 ( .A(n535), .B(KEYINPUT4), .ZN(n539) );
  NOR2_X4 U599 ( .A1(n537), .A2(n536), .ZN(n655) );
  NAND2_X1 U600 ( .A1(G76), .A2(n655), .ZN(n538) );
  NAND2_X1 U601 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U602 ( .A(n540), .B(KEYINPUT5), .Z(n541) );
  NOR2_X1 U603 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U604 ( .A(KEYINPUT78), .B(n543), .Z(n544) );
  XNOR2_X2 U605 ( .A(KEYINPUT7), .B(n544), .ZN(G168) );
  NAND2_X1 U606 ( .A1(G64), .A2(n651), .ZN(n546) );
  NAND2_X1 U607 ( .A1(G52), .A2(n659), .ZN(n545) );
  NAND2_X1 U608 ( .A1(n546), .A2(n545), .ZN(n552) );
  NAND2_X1 U609 ( .A1(G77), .A2(n655), .ZN(n548) );
  NAND2_X1 U610 ( .A1(G90), .A2(n652), .ZN(n547) );
  NAND2_X1 U611 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U612 ( .A(KEYINPUT69), .B(n549), .ZN(n550) );
  XNOR2_X1 U613 ( .A(KEYINPUT9), .B(n550), .ZN(n551) );
  NAND2_X1 U614 ( .A1(n553), .A2(G137), .ZN(n554) );
  XNOR2_X1 U615 ( .A(n554), .B(KEYINPUT66), .ZN(n556) );
  NAND2_X1 U616 ( .A1(G113), .A2(n561), .ZN(n555) );
  NAND2_X1 U617 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U618 ( .A(n557), .B(KEYINPUT67), .ZN(n559) );
  NAND2_X1 U619 ( .A1(G125), .A2(n890), .ZN(n558) );
  AND2_X1 U620 ( .A1(n559), .A2(n558), .ZN(n688) );
  NAND2_X1 U621 ( .A1(G101), .A2(n886), .ZN(n560) );
  XOR2_X1 U622 ( .A(KEYINPUT23), .B(n560), .Z(n687) );
  AND2_X1 U623 ( .A1(n688), .A2(n687), .ZN(G160) );
  AND2_X1 U624 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U625 ( .A1(n886), .A2(G99), .ZN(n568) );
  NAND2_X1 U626 ( .A1(G135), .A2(n885), .ZN(n563) );
  NAND2_X1 U627 ( .A1(G111), .A2(n561), .ZN(n562) );
  NAND2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n566) );
  NAND2_X1 U629 ( .A1(n890), .A2(G123), .ZN(n564) );
  XOR2_X1 U630 ( .A(KEYINPUT18), .B(n564), .Z(n565) );
  NOR2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U632 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U633 ( .A(KEYINPUT83), .B(n569), .Z(n987) );
  XNOR2_X1 U634 ( .A(G2096), .B(n987), .ZN(n570) );
  OR2_X1 U635 ( .A1(G2100), .A2(n570), .ZN(G156) );
  INV_X1 U636 ( .A(G132), .ZN(G219) );
  INV_X1 U637 ( .A(G82), .ZN(G220) );
  INV_X1 U638 ( .A(G57), .ZN(G237) );
  XOR2_X1 U639 ( .A(KEYINPUT10), .B(KEYINPUT71), .Z(n572) );
  NAND2_X1 U640 ( .A1(G7), .A2(G661), .ZN(n571) );
  XNOR2_X1 U641 ( .A(n572), .B(n571), .ZN(G223) );
  INV_X1 U642 ( .A(G223), .ZN(n833) );
  NAND2_X1 U643 ( .A1(n833), .A2(G567), .ZN(n573) );
  XOR2_X1 U644 ( .A(KEYINPUT11), .B(n573), .Z(G234) );
  XOR2_X1 U645 ( .A(KEYINPUT12), .B(KEYINPUT73), .Z(n575) );
  NAND2_X1 U646 ( .A1(G81), .A2(n652), .ZN(n574) );
  XNOR2_X1 U647 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U648 ( .A(KEYINPUT72), .B(n576), .ZN(n579) );
  NAND2_X1 U649 ( .A1(n655), .A2(G68), .ZN(n577) );
  XNOR2_X1 U650 ( .A(KEYINPUT74), .B(n577), .ZN(n578) );
  NAND2_X1 U651 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U652 ( .A(n580), .B(KEYINPUT13), .ZN(n582) );
  NAND2_X1 U653 ( .A1(G43), .A2(n659), .ZN(n581) );
  NAND2_X1 U654 ( .A1(n582), .A2(n581), .ZN(n585) );
  NAND2_X1 U655 ( .A1(n651), .A2(G56), .ZN(n583) );
  XOR2_X1 U656 ( .A(KEYINPUT14), .B(n583), .Z(n584) );
  NOR2_X1 U657 ( .A1(n585), .A2(n584), .ZN(n934) );
  NAND2_X1 U658 ( .A1(n934), .A2(G860), .ZN(G153) );
  INV_X1 U659 ( .A(G868), .ZN(n617) );
  NOR2_X1 U660 ( .A1(n617), .A2(G171), .ZN(n586) );
  XNOR2_X1 U661 ( .A(n586), .B(KEYINPUT75), .ZN(n598) );
  NAND2_X1 U662 ( .A1(G92), .A2(n652), .ZN(n594) );
  NAND2_X1 U663 ( .A1(G66), .A2(n651), .ZN(n588) );
  NAND2_X1 U664 ( .A1(G79), .A2(n655), .ZN(n587) );
  NAND2_X1 U665 ( .A1(n588), .A2(n587), .ZN(n592) );
  NAND2_X1 U666 ( .A1(n589), .A2(G54), .ZN(n590) );
  XOR2_X1 U667 ( .A(KEYINPUT76), .B(n590), .Z(n591) );
  NOR2_X1 U668 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U669 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U670 ( .A(n595), .B(KEYINPUT15), .ZN(n596) );
  XNOR2_X1 U671 ( .A(KEYINPUT77), .B(n596), .ZN(n614) );
  NAND2_X1 U672 ( .A1(n617), .A2(n614), .ZN(n597) );
  NAND2_X1 U673 ( .A1(n598), .A2(n597), .ZN(G284) );
  NAND2_X1 U674 ( .A1(G65), .A2(n651), .ZN(n600) );
  NAND2_X1 U675 ( .A1(G91), .A2(n652), .ZN(n599) );
  NAND2_X1 U676 ( .A1(n600), .A2(n599), .ZN(n603) );
  NAND2_X1 U677 ( .A1(n655), .A2(G78), .ZN(n601) );
  XOR2_X1 U678 ( .A(KEYINPUT70), .B(n601), .Z(n602) );
  NOR2_X1 U679 ( .A1(n603), .A2(n602), .ZN(n605) );
  NAND2_X1 U680 ( .A1(n659), .A2(G53), .ZN(n604) );
  NAND2_X1 U681 ( .A1(n605), .A2(n604), .ZN(G299) );
  NOR2_X1 U682 ( .A1(G286), .A2(n617), .ZN(n607) );
  NOR2_X1 U683 ( .A1(G868), .A2(G299), .ZN(n606) );
  NOR2_X1 U684 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U685 ( .A(KEYINPUT79), .B(n608), .Z(G297) );
  INV_X1 U686 ( .A(G559), .ZN(n609) );
  NOR2_X1 U687 ( .A1(G860), .A2(n609), .ZN(n610) );
  XNOR2_X1 U688 ( .A(n610), .B(KEYINPUT80), .ZN(n611) );
  NOR2_X1 U689 ( .A1(n614), .A2(n611), .ZN(n612) );
  XNOR2_X1 U690 ( .A(n612), .B(KEYINPUT16), .ZN(n613) );
  XNOR2_X1 U691 ( .A(n613), .B(KEYINPUT81), .ZN(G148) );
  INV_X1 U692 ( .A(n614), .ZN(n924) );
  NAND2_X1 U693 ( .A1(n924), .A2(G868), .ZN(n615) );
  NOR2_X1 U694 ( .A1(G559), .A2(n615), .ZN(n616) );
  XNOR2_X1 U695 ( .A(n616), .B(KEYINPUT82), .ZN(n619) );
  AND2_X1 U696 ( .A1(n934), .A2(n617), .ZN(n618) );
  NOR2_X1 U697 ( .A1(n619), .A2(n618), .ZN(G282) );
  NAND2_X1 U698 ( .A1(G67), .A2(n651), .ZN(n621) );
  NAND2_X1 U699 ( .A1(G55), .A2(n659), .ZN(n620) );
  NAND2_X1 U700 ( .A1(n621), .A2(n620), .ZN(n625) );
  NAND2_X1 U701 ( .A1(G80), .A2(n655), .ZN(n623) );
  NAND2_X1 U702 ( .A1(G93), .A2(n652), .ZN(n622) );
  NAND2_X1 U703 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U704 ( .A1(n625), .A2(n624), .ZN(n667) );
  NAND2_X1 U705 ( .A1(G559), .A2(n924), .ZN(n626) );
  XOR2_X1 U706 ( .A(n934), .B(n626), .Z(n670) );
  XNOR2_X1 U707 ( .A(KEYINPUT84), .B(n670), .ZN(n627) );
  NOR2_X1 U708 ( .A1(G860), .A2(n627), .ZN(n628) );
  XNOR2_X1 U709 ( .A(n667), .B(n628), .ZN(G145) );
  AND2_X1 U710 ( .A1(n651), .A2(G60), .ZN(n632) );
  NAND2_X1 U711 ( .A1(G72), .A2(n655), .ZN(n630) );
  NAND2_X1 U712 ( .A1(G85), .A2(n652), .ZN(n629) );
  NAND2_X1 U713 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U714 ( .A1(n632), .A2(n631), .ZN(n634) );
  NAND2_X1 U715 ( .A1(n659), .A2(G47), .ZN(n633) );
  NAND2_X1 U716 ( .A1(n634), .A2(n633), .ZN(G290) );
  NAND2_X1 U717 ( .A1(G62), .A2(n651), .ZN(n636) );
  NAND2_X1 U718 ( .A1(G75), .A2(n655), .ZN(n635) );
  NAND2_X1 U719 ( .A1(n636), .A2(n635), .ZN(n642) );
  NAND2_X1 U720 ( .A1(G50), .A2(n659), .ZN(n637) );
  XNOR2_X1 U721 ( .A(n637), .B(KEYINPUT88), .ZN(n640) );
  NAND2_X1 U722 ( .A1(G88), .A2(n652), .ZN(n638) );
  XOR2_X1 U723 ( .A(KEYINPUT89), .B(n638), .Z(n639) );
  NAND2_X1 U724 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U725 ( .A1(n642), .A2(n641), .ZN(G166) );
  NAND2_X1 U726 ( .A1(G651), .A2(G74), .ZN(n643) );
  XOR2_X1 U727 ( .A(KEYINPUT85), .B(n643), .Z(n645) );
  NAND2_X1 U728 ( .A1(n659), .A2(G49), .ZN(n644) );
  NAND2_X1 U729 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U730 ( .A(KEYINPUT86), .B(n646), .ZN(n647) );
  NOR2_X1 U731 ( .A1(n651), .A2(n647), .ZN(n648) );
  XOR2_X1 U732 ( .A(KEYINPUT87), .B(n648), .Z(n650) );
  NAND2_X1 U733 ( .A1(G87), .A2(n536), .ZN(n649) );
  NAND2_X1 U734 ( .A1(n650), .A2(n649), .ZN(G288) );
  NAND2_X1 U735 ( .A1(G61), .A2(n651), .ZN(n654) );
  NAND2_X1 U736 ( .A1(G86), .A2(n652), .ZN(n653) );
  NAND2_X1 U737 ( .A1(n654), .A2(n653), .ZN(n658) );
  NAND2_X1 U738 ( .A1(n655), .A2(G73), .ZN(n656) );
  XOR2_X1 U739 ( .A(KEYINPUT2), .B(n656), .Z(n657) );
  NOR2_X1 U740 ( .A1(n658), .A2(n657), .ZN(n661) );
  NAND2_X1 U741 ( .A1(n659), .A2(G48), .ZN(n660) );
  NAND2_X1 U742 ( .A1(n661), .A2(n660), .ZN(G305) );
  NOR2_X1 U743 ( .A1(G868), .A2(n667), .ZN(n662) );
  XNOR2_X1 U744 ( .A(n662), .B(KEYINPUT91), .ZN(n673) );
  XOR2_X1 U745 ( .A(KEYINPUT19), .B(KEYINPUT90), .Z(n663) );
  XNOR2_X1 U746 ( .A(G290), .B(n663), .ZN(n666) );
  XNOR2_X1 U747 ( .A(G166), .B(G288), .ZN(n664) );
  XNOR2_X1 U748 ( .A(n664), .B(G299), .ZN(n665) );
  XNOR2_X1 U749 ( .A(n666), .B(n665), .ZN(n669) );
  XNOR2_X1 U750 ( .A(G305), .B(n667), .ZN(n668) );
  XNOR2_X1 U751 ( .A(n669), .B(n668), .ZN(n901) );
  XNOR2_X1 U752 ( .A(n901), .B(n670), .ZN(n671) );
  NAND2_X1 U753 ( .A1(G868), .A2(n671), .ZN(n672) );
  NAND2_X1 U754 ( .A1(n673), .A2(n672), .ZN(G295) );
  NAND2_X1 U755 ( .A1(G2078), .A2(G2084), .ZN(n674) );
  XOR2_X1 U756 ( .A(KEYINPUT20), .B(n674), .Z(n675) );
  NAND2_X1 U757 ( .A1(G2090), .A2(n675), .ZN(n676) );
  XNOR2_X1 U758 ( .A(KEYINPUT21), .B(n676), .ZN(n677) );
  NAND2_X1 U759 ( .A1(n677), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U760 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U761 ( .A1(G120), .A2(G108), .ZN(n678) );
  NOR2_X1 U762 ( .A1(G237), .A2(n678), .ZN(n679) );
  NAND2_X1 U763 ( .A1(G69), .A2(n679), .ZN(n838) );
  NAND2_X1 U764 ( .A1(G567), .A2(n838), .ZN(n680) );
  XNOR2_X1 U765 ( .A(n680), .B(KEYINPUT92), .ZN(n685) );
  NOR2_X1 U766 ( .A1(G220), .A2(G219), .ZN(n681) );
  XOR2_X1 U767 ( .A(KEYINPUT22), .B(n681), .Z(n682) );
  NOR2_X1 U768 ( .A1(G218), .A2(n682), .ZN(n683) );
  NAND2_X1 U769 ( .A1(G96), .A2(n683), .ZN(n839) );
  NAND2_X1 U770 ( .A1(G2106), .A2(n839), .ZN(n684) );
  NAND2_X1 U771 ( .A1(n685), .A2(n684), .ZN(n840) );
  NAND2_X1 U772 ( .A1(G483), .A2(G661), .ZN(n686) );
  NOR2_X1 U773 ( .A1(n840), .A2(n686), .ZN(n835) );
  NAND2_X1 U774 ( .A1(n835), .A2(G36), .ZN(G176) );
  INV_X1 U775 ( .A(G166), .ZN(G303) );
  XOR2_X1 U776 ( .A(G1996), .B(KEYINPUT97), .Z(n958) );
  XNOR2_X1 U777 ( .A(KEYINPUT64), .B(KEYINPUT26), .ZN(n695) );
  NOR2_X1 U778 ( .A1(n958), .A2(n695), .ZN(n702) );
  AND2_X1 U779 ( .A1(G40), .A2(n687), .ZN(n689) );
  AND2_X1 U780 ( .A1(n689), .A2(n688), .ZN(n799) );
  NAND2_X2 U781 ( .A1(n801), .A2(n799), .ZN(n727) );
  NAND2_X1 U782 ( .A1(G1348), .A2(n727), .ZN(n690) );
  XNOR2_X1 U783 ( .A(n690), .B(KEYINPUT98), .ZN(n692) );
  INV_X1 U784 ( .A(n727), .ZN(n717) );
  NAND2_X1 U785 ( .A1(n717), .A2(G2067), .ZN(n691) );
  NAND2_X1 U786 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U787 ( .A(KEYINPUT99), .B(n693), .ZN(n707) );
  NOR2_X1 U788 ( .A1(n924), .A2(n707), .ZN(n700) );
  INV_X1 U789 ( .A(G1341), .ZN(n1005) );
  NAND2_X1 U790 ( .A1(n1005), .A2(n695), .ZN(n694) );
  NAND2_X1 U791 ( .A1(n694), .A2(n727), .ZN(n698) );
  AND2_X1 U792 ( .A1(n717), .A2(n958), .ZN(n696) );
  NAND2_X1 U793 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U794 ( .A1(n519), .A2(n934), .ZN(n699) );
  OR2_X1 U795 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U796 ( .A1(n702), .A2(n701), .ZN(n710) );
  NAND2_X1 U797 ( .A1(G2072), .A2(n717), .ZN(n704) );
  AND2_X1 U798 ( .A1(n727), .A2(G1956), .ZN(n705) );
  NOR2_X1 U799 ( .A1(n706), .A2(n705), .ZN(n711) );
  INV_X1 U800 ( .A(G299), .ZN(n929) );
  NAND2_X1 U801 ( .A1(n711), .A2(n929), .ZN(n708) );
  NAND2_X1 U802 ( .A1(n708), .A2(n520), .ZN(n709) );
  NOR2_X1 U803 ( .A1(n711), .A2(n929), .ZN(n712) );
  XOR2_X1 U804 ( .A(n712), .B(KEYINPUT28), .Z(n713) );
  NAND2_X1 U805 ( .A1(n714), .A2(n713), .ZN(n716) );
  XNOR2_X1 U806 ( .A(KEYINPUT95), .B(G1961), .ZN(n1014) );
  NAND2_X1 U807 ( .A1(n727), .A2(n1014), .ZN(n719) );
  XNOR2_X1 U808 ( .A(KEYINPUT25), .B(G2078), .ZN(n957) );
  NAND2_X1 U809 ( .A1(n717), .A2(n957), .ZN(n718) );
  NAND2_X1 U810 ( .A1(n719), .A2(n718), .ZN(n731) );
  NAND2_X1 U811 ( .A1(n731), .A2(G171), .ZN(n746) );
  NOR2_X1 U812 ( .A1(G1971), .A2(n781), .ZN(n720) );
  XNOR2_X1 U813 ( .A(n720), .B(KEYINPUT100), .ZN(n722) );
  NOR2_X1 U814 ( .A1(n727), .A2(G2090), .ZN(n721) );
  NOR2_X1 U815 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U816 ( .A1(n723), .A2(G303), .ZN(n735) );
  INV_X1 U817 ( .A(n735), .ZN(n724) );
  OR2_X1 U818 ( .A1(n724), .A2(G286), .ZN(n726) );
  AND2_X1 U819 ( .A1(n746), .A2(n726), .ZN(n725) );
  NAND2_X1 U820 ( .A1(n745), .A2(n725), .ZN(n739) );
  INV_X1 U821 ( .A(n726), .ZN(n737) );
  NOR2_X1 U822 ( .A1(G1966), .A2(n781), .ZN(n750) );
  NOR2_X1 U823 ( .A1(G2084), .A2(n727), .ZN(n744) );
  NOR2_X1 U824 ( .A1(n750), .A2(n744), .ZN(n728) );
  NAND2_X1 U825 ( .A1(G8), .A2(n728), .ZN(n729) );
  XNOR2_X1 U826 ( .A(KEYINPUT30), .B(n729), .ZN(n730) );
  NOR2_X1 U827 ( .A1(G168), .A2(n730), .ZN(n733) );
  NOR2_X1 U828 ( .A1(G171), .A2(n731), .ZN(n732) );
  NOR2_X1 U829 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U830 ( .A(KEYINPUT31), .B(n734), .Z(n747) );
  AND2_X1 U831 ( .A1(n747), .A2(n735), .ZN(n736) );
  NAND2_X1 U832 ( .A1(n739), .A2(n738), .ZN(n741) );
  XNOR2_X1 U833 ( .A(n741), .B(n740), .ZN(n742) );
  NAND2_X1 U834 ( .A1(n742), .A2(G8), .ZN(n743) );
  XNOR2_X1 U835 ( .A(n743), .B(KEYINPUT32), .ZN(n770) );
  NAND2_X1 U836 ( .A1(G8), .A2(n744), .ZN(n752) );
  NAND2_X1 U837 ( .A1(n746), .A2(n745), .ZN(n748) );
  AND2_X1 U838 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U839 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U840 ( .A1(n752), .A2(n751), .ZN(n771) );
  NAND2_X1 U841 ( .A1(G1976), .A2(G288), .ZN(n935) );
  INV_X1 U842 ( .A(n781), .ZN(n753) );
  NAND2_X1 U843 ( .A1(n935), .A2(n753), .ZN(n757) );
  INV_X1 U844 ( .A(n757), .ZN(n754) );
  AND2_X1 U845 ( .A1(n771), .A2(n754), .ZN(n755) );
  NAND2_X1 U846 ( .A1(n770), .A2(n755), .ZN(n760) );
  NOR2_X1 U847 ( .A1(G1976), .A2(G288), .ZN(n763) );
  NOR2_X1 U848 ( .A1(G1971), .A2(G303), .ZN(n756) );
  NOR2_X1 U849 ( .A1(n763), .A2(n756), .ZN(n944) );
  NOR2_X1 U850 ( .A1(n757), .A2(n944), .ZN(n758) );
  NOR2_X1 U851 ( .A1(n758), .A2(KEYINPUT33), .ZN(n759) );
  NAND2_X1 U852 ( .A1(n760), .A2(n759), .ZN(n762) );
  NAND2_X1 U853 ( .A1(n763), .A2(KEYINPUT33), .ZN(n764) );
  NOR2_X1 U854 ( .A1(n781), .A2(n764), .ZN(n765) );
  XOR2_X1 U855 ( .A(KEYINPUT103), .B(n765), .Z(n766) );
  NOR2_X2 U856 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U857 ( .A(n768), .B(KEYINPUT104), .ZN(n769) );
  XOR2_X1 U858 ( .A(G1981), .B(G305), .Z(n941) );
  NAND2_X1 U859 ( .A1(n769), .A2(n941), .ZN(n777) );
  NAND2_X1 U860 ( .A1(n771), .A2(n770), .ZN(n774) );
  NOR2_X1 U861 ( .A1(G2090), .A2(G303), .ZN(n772) );
  NAND2_X1 U862 ( .A1(G8), .A2(n772), .ZN(n773) );
  NAND2_X1 U863 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U864 ( .A1(n781), .A2(n775), .ZN(n776) );
  NAND2_X1 U865 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U866 ( .A(n778), .B(KEYINPUT105), .ZN(n783) );
  NOR2_X1 U867 ( .A1(G1981), .A2(G305), .ZN(n779) );
  XOR2_X1 U868 ( .A(n779), .B(KEYINPUT24), .Z(n780) );
  NOR2_X1 U869 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U870 ( .A1(n783), .A2(n518), .ZN(n815) );
  NAND2_X1 U871 ( .A1(G131), .A2(n885), .ZN(n785) );
  NAND2_X1 U872 ( .A1(G107), .A2(n561), .ZN(n784) );
  NAND2_X1 U873 ( .A1(n785), .A2(n784), .ZN(n789) );
  NAND2_X1 U874 ( .A1(G95), .A2(n886), .ZN(n787) );
  NAND2_X1 U875 ( .A1(G119), .A2(n890), .ZN(n786) );
  NAND2_X1 U876 ( .A1(n787), .A2(n786), .ZN(n788) );
  NOR2_X1 U877 ( .A1(n789), .A2(n788), .ZN(n880) );
  INV_X1 U878 ( .A(G1991), .ZN(n858) );
  NOR2_X1 U879 ( .A1(n880), .A2(n858), .ZN(n798) );
  NAND2_X1 U880 ( .A1(G141), .A2(n885), .ZN(n791) );
  NAND2_X1 U881 ( .A1(G117), .A2(n561), .ZN(n790) );
  NAND2_X1 U882 ( .A1(n791), .A2(n790), .ZN(n794) );
  NAND2_X1 U883 ( .A1(n886), .A2(G105), .ZN(n792) );
  XOR2_X1 U884 ( .A(KEYINPUT38), .B(n792), .Z(n793) );
  NOR2_X1 U885 ( .A1(n794), .A2(n793), .ZN(n796) );
  NAND2_X1 U886 ( .A1(n890), .A2(G129), .ZN(n795) );
  NAND2_X1 U887 ( .A1(n796), .A2(n795), .ZN(n877) );
  AND2_X1 U888 ( .A1(G1996), .A2(n877), .ZN(n797) );
  NOR2_X1 U889 ( .A1(n798), .A2(n797), .ZN(n988) );
  INV_X1 U890 ( .A(n799), .ZN(n800) );
  NOR2_X1 U891 ( .A1(n801), .A2(n800), .ZN(n828) );
  INV_X1 U892 ( .A(n828), .ZN(n802) );
  NOR2_X1 U893 ( .A1(n988), .A2(n802), .ZN(n819) );
  INV_X1 U894 ( .A(n819), .ZN(n812) );
  NAND2_X1 U895 ( .A1(G140), .A2(n885), .ZN(n804) );
  NAND2_X1 U896 ( .A1(G104), .A2(n886), .ZN(n803) );
  NAND2_X1 U897 ( .A1(n804), .A2(n803), .ZN(n805) );
  XNOR2_X1 U898 ( .A(KEYINPUT34), .B(n805), .ZN(n810) );
  NAND2_X1 U899 ( .A1(G116), .A2(n561), .ZN(n807) );
  NAND2_X1 U900 ( .A1(G128), .A2(n890), .ZN(n806) );
  NAND2_X1 U901 ( .A1(n807), .A2(n806), .ZN(n808) );
  XOR2_X1 U902 ( .A(KEYINPUT35), .B(n808), .Z(n809) );
  NOR2_X1 U903 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U904 ( .A(KEYINPUT36), .B(n811), .ZN(n896) );
  XNOR2_X1 U905 ( .A(G2067), .B(KEYINPUT37), .ZN(n825) );
  NOR2_X1 U906 ( .A1(n896), .A2(n825), .ZN(n986) );
  NAND2_X1 U907 ( .A1(n828), .A2(n986), .ZN(n823) );
  NAND2_X1 U908 ( .A1(n812), .A2(n823), .ZN(n813) );
  XOR2_X1 U909 ( .A(KEYINPUT93), .B(n813), .Z(n814) );
  XNOR2_X1 U910 ( .A(G1986), .B(G290), .ZN(n931) );
  NAND2_X1 U911 ( .A1(n815), .A2(n515), .ZN(n831) );
  XOR2_X1 U912 ( .A(KEYINPUT39), .B(KEYINPUT107), .Z(n822) );
  NOR2_X1 U913 ( .A1(n877), .A2(G1996), .ZN(n816) );
  XNOR2_X1 U914 ( .A(n816), .B(KEYINPUT106), .ZN(n982) );
  NOR2_X1 U915 ( .A1(G1986), .A2(G290), .ZN(n817) );
  AND2_X1 U916 ( .A1(n858), .A2(n880), .ZN(n990) );
  NOR2_X1 U917 ( .A1(n817), .A2(n990), .ZN(n818) );
  NOR2_X1 U918 ( .A1(n819), .A2(n818), .ZN(n820) );
  NOR2_X1 U919 ( .A1(n982), .A2(n820), .ZN(n821) );
  XNOR2_X1 U920 ( .A(n822), .B(n821), .ZN(n824) );
  NAND2_X1 U921 ( .A1(n824), .A2(n823), .ZN(n826) );
  NAND2_X1 U922 ( .A1(n896), .A2(n825), .ZN(n991) );
  NAND2_X1 U923 ( .A1(n826), .A2(n991), .ZN(n827) );
  XNOR2_X1 U924 ( .A(KEYINPUT108), .B(n827), .ZN(n829) );
  NAND2_X1 U925 ( .A1(n829), .A2(n828), .ZN(n830) );
  NAND2_X1 U926 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U927 ( .A(n832), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n833), .ZN(G217) );
  AND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U930 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U931 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U932 ( .A1(n836), .A2(n835), .ZN(n837) );
  XOR2_X1 U933 ( .A(KEYINPUT111), .B(n837), .Z(G188) );
  XOR2_X1 U934 ( .A(G108), .B(KEYINPUT118), .Z(G238) );
  INV_X1 U936 ( .A(G120), .ZN(G236) );
  INV_X1 U937 ( .A(G96), .ZN(G221) );
  NOR2_X1 U938 ( .A1(n839), .A2(n838), .ZN(G325) );
  INV_X1 U939 ( .A(G325), .ZN(G261) );
  XOR2_X1 U940 ( .A(KEYINPUT112), .B(n840), .Z(G319) );
  XOR2_X1 U941 ( .A(G2100), .B(G2096), .Z(n842) );
  XNOR2_X1 U942 ( .A(KEYINPUT42), .B(G2678), .ZN(n841) );
  XNOR2_X1 U943 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U944 ( .A(KEYINPUT43), .B(G2090), .Z(n844) );
  XNOR2_X1 U945 ( .A(G2067), .B(G2072), .ZN(n843) );
  XNOR2_X1 U946 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U947 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U948 ( .A(G2078), .B(G2084), .ZN(n847) );
  XNOR2_X1 U949 ( .A(n848), .B(n847), .ZN(G227) );
  XOR2_X1 U950 ( .A(G1961), .B(G1966), .Z(n850) );
  XNOR2_X1 U951 ( .A(G1996), .B(G1976), .ZN(n849) );
  XNOR2_X1 U952 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U953 ( .A(G1956), .B(G1971), .Z(n852) );
  XNOR2_X1 U954 ( .A(G1986), .B(G1981), .ZN(n851) );
  XNOR2_X1 U955 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U956 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U957 ( .A(G2474), .B(KEYINPUT113), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n856), .B(n855), .ZN(n857) );
  XNOR2_X1 U959 ( .A(KEYINPUT41), .B(n857), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n859), .B(n858), .ZN(G229) );
  NAND2_X1 U961 ( .A1(G124), .A2(n890), .ZN(n860) );
  XNOR2_X1 U962 ( .A(n860), .B(KEYINPUT44), .ZN(n862) );
  NAND2_X1 U963 ( .A1(n561), .A2(G112), .ZN(n861) );
  NAND2_X1 U964 ( .A1(n862), .A2(n861), .ZN(n866) );
  NAND2_X1 U965 ( .A1(G136), .A2(n885), .ZN(n864) );
  NAND2_X1 U966 ( .A1(G100), .A2(n886), .ZN(n863) );
  NAND2_X1 U967 ( .A1(n864), .A2(n863), .ZN(n865) );
  NOR2_X1 U968 ( .A1(n866), .A2(n865), .ZN(G162) );
  NAND2_X1 U969 ( .A1(G118), .A2(n561), .ZN(n868) );
  NAND2_X1 U970 ( .A1(G130), .A2(n890), .ZN(n867) );
  NAND2_X1 U971 ( .A1(n868), .A2(n867), .ZN(n873) );
  NAND2_X1 U972 ( .A1(G142), .A2(n885), .ZN(n870) );
  NAND2_X1 U973 ( .A1(G106), .A2(n886), .ZN(n869) );
  NAND2_X1 U974 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U975 ( .A(KEYINPUT45), .B(n871), .Z(n872) );
  NOR2_X1 U976 ( .A1(n873), .A2(n872), .ZN(n884) );
  XOR2_X1 U977 ( .A(KEYINPUT48), .B(KEYINPUT114), .Z(n875) );
  XNOR2_X1 U978 ( .A(KEYINPUT116), .B(KEYINPUT46), .ZN(n874) );
  XNOR2_X1 U979 ( .A(n875), .B(n874), .ZN(n876) );
  XOR2_X1 U980 ( .A(n876), .B(G162), .Z(n879) );
  XOR2_X1 U981 ( .A(G164), .B(n877), .Z(n878) );
  XNOR2_X1 U982 ( .A(n879), .B(n878), .ZN(n881) );
  XOR2_X1 U983 ( .A(n881), .B(n880), .Z(n882) );
  XNOR2_X1 U984 ( .A(n882), .B(n987), .ZN(n883) );
  XNOR2_X1 U985 ( .A(n884), .B(n883), .ZN(n898) );
  NAND2_X1 U986 ( .A1(G139), .A2(n885), .ZN(n888) );
  NAND2_X1 U987 ( .A1(G103), .A2(n886), .ZN(n887) );
  NAND2_X1 U988 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U989 ( .A(KEYINPUT115), .B(n889), .Z(n895) );
  NAND2_X1 U990 ( .A1(G115), .A2(n561), .ZN(n892) );
  NAND2_X1 U991 ( .A1(G127), .A2(n890), .ZN(n891) );
  NAND2_X1 U992 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U993 ( .A(KEYINPUT47), .B(n893), .Z(n894) );
  NOR2_X1 U994 ( .A1(n895), .A2(n894), .ZN(n976) );
  XNOR2_X1 U995 ( .A(n896), .B(n976), .ZN(n897) );
  XNOR2_X1 U996 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U997 ( .A(n899), .B(G160), .ZN(n900) );
  NOR2_X1 U998 ( .A1(G37), .A2(n900), .ZN(G395) );
  XOR2_X1 U999 ( .A(KEYINPUT117), .B(n901), .Z(n903) );
  XNOR2_X1 U1000 ( .A(G171), .B(n924), .ZN(n902) );
  XNOR2_X1 U1001 ( .A(n903), .B(n902), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(G286), .B(n934), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n906), .ZN(G397) );
  XNOR2_X1 U1005 ( .A(G2446), .B(G2443), .ZN(n916) );
  XOR2_X1 U1006 ( .A(G2430), .B(KEYINPUT110), .Z(n908) );
  XNOR2_X1 U1007 ( .A(G2454), .B(G2435), .ZN(n907) );
  XNOR2_X1 U1008 ( .A(n908), .B(n907), .ZN(n912) );
  XOR2_X1 U1009 ( .A(G2438), .B(G2427), .Z(n910) );
  XNOR2_X1 U1010 ( .A(G1341), .B(G1348), .ZN(n909) );
  XNOR2_X1 U1011 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1012 ( .A(n912), .B(n911), .Z(n914) );
  XNOR2_X1 U1013 ( .A(KEYINPUT109), .B(G2451), .ZN(n913) );
  XNOR2_X1 U1014 ( .A(n914), .B(n913), .ZN(n915) );
  XNOR2_X1 U1015 ( .A(n916), .B(n915), .ZN(n917) );
  NAND2_X1 U1016 ( .A1(n917), .A2(G14), .ZN(n923) );
  NAND2_X1 U1017 ( .A1(n923), .A2(G319), .ZN(n920) );
  NOR2_X1 U1018 ( .A1(G227), .A2(G229), .ZN(n918) );
  XNOR2_X1 U1019 ( .A(KEYINPUT49), .B(n918), .ZN(n919) );
  NOR2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n922) );
  NOR2_X1 U1021 ( .A1(G395), .A2(G397), .ZN(n921) );
  NAND2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(G225) );
  INV_X1 U1023 ( .A(G225), .ZN(G308) );
  INV_X1 U1024 ( .A(G69), .ZN(G235) );
  INV_X1 U1025 ( .A(n923), .ZN(G401) );
  XOR2_X1 U1026 ( .A(G16), .B(KEYINPUT56), .Z(n950) );
  XNOR2_X1 U1027 ( .A(n924), .B(G1348), .ZN(n927) );
  XNOR2_X1 U1028 ( .A(G171), .B(G1961), .ZN(n925) );
  XNOR2_X1 U1029 ( .A(n925), .B(KEYINPUT124), .ZN(n926) );
  NAND2_X1 U1030 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1031 ( .A(n928), .B(KEYINPUT125), .ZN(n940) );
  XNOR2_X1 U1032 ( .A(n929), .B(G1956), .ZN(n933) );
  AND2_X1 U1033 ( .A1(G303), .A2(G1971), .ZN(n930) );
  NOR2_X1 U1034 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1035 ( .A1(n933), .A2(n932), .ZN(n938) );
  XNOR2_X1 U1036 ( .A(n934), .B(G1341), .ZN(n936) );
  NAND2_X1 U1037 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n947) );
  XNOR2_X1 U1040 ( .A(G1966), .B(G168), .ZN(n942) );
  NAND2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1042 ( .A(KEYINPUT57), .B(n943), .ZN(n945) );
  NAND2_X1 U1043 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1044 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1045 ( .A(n948), .B(KEYINPUT126), .ZN(n949) );
  NOR2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n975) );
  XOR2_X1 U1047 ( .A(KEYINPUT122), .B(G29), .Z(n971) );
  XNOR2_X1 U1048 ( .A(G1991), .B(G25), .ZN(n952) );
  XNOR2_X1 U1049 ( .A(G33), .B(G2072), .ZN(n951) );
  NOR2_X1 U1050 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1051 ( .A1(G28), .A2(n953), .ZN(n956) );
  XOR2_X1 U1052 ( .A(KEYINPUT121), .B(G2067), .Z(n954) );
  XNOR2_X1 U1053 ( .A(G26), .B(n954), .ZN(n955) );
  NOR2_X1 U1054 ( .A1(n956), .A2(n955), .ZN(n962) );
  XOR2_X1 U1055 ( .A(n957), .B(G27), .Z(n960) );
  XNOR2_X1 U1056 ( .A(G32), .B(n958), .ZN(n959) );
  NOR2_X1 U1057 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1059 ( .A(n963), .B(KEYINPUT53), .ZN(n966) );
  XOR2_X1 U1060 ( .A(G2084), .B(G34), .Z(n964) );
  XNOR2_X1 U1061 ( .A(KEYINPUT54), .B(n964), .ZN(n965) );
  NAND2_X1 U1062 ( .A1(n966), .A2(n965), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(G35), .B(G2090), .ZN(n967) );
  NOR2_X1 U1064 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1065 ( .A(KEYINPUT55), .B(n969), .ZN(n970) );
  NAND2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1067 ( .A1(G11), .A2(n972), .ZN(n973) );
  XOR2_X1 U1068 ( .A(KEYINPUT123), .B(n973), .Z(n974) );
  NOR2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n1004) );
  XNOR2_X1 U1070 ( .A(G2072), .B(n976), .ZN(n979) );
  XNOR2_X1 U1071 ( .A(G164), .B(G2078), .ZN(n977) );
  XNOR2_X1 U1072 ( .A(n977), .B(KEYINPUT120), .ZN(n978) );
  NAND2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1074 ( .A(n980), .B(KEYINPUT50), .ZN(n998) );
  XOR2_X1 U1075 ( .A(G2090), .B(G162), .Z(n981) );
  NOR2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  XOR2_X1 U1077 ( .A(KEYINPUT51), .B(n983), .Z(n984) );
  XNOR2_X1 U1078 ( .A(n984), .B(KEYINPUT119), .ZN(n985) );
  NOR2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n996) );
  NAND2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n992) );
  NAND2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n994) );
  XOR2_X1 U1083 ( .A(G160), .B(G2084), .Z(n993) );
  NOR2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1086 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1087 ( .A(KEYINPUT52), .B(n999), .ZN(n1001) );
  INV_X1 U1088 ( .A(KEYINPUT55), .ZN(n1000) );
  NAND2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1090 ( .A1(n1002), .A2(G29), .ZN(n1003) );
  NAND2_X1 U1091 ( .A1(n1004), .A2(n1003), .ZN(n1030) );
  XNOR2_X1 U1092 ( .A(G19), .B(n1005), .ZN(n1009) );
  XNOR2_X1 U1093 ( .A(G1981), .B(G6), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(G1956), .B(G20), .ZN(n1006) );
  NOR2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1012) );
  XOR2_X1 U1097 ( .A(KEYINPUT59), .B(G1348), .Z(n1010) );
  XNOR2_X1 U1098 ( .A(G4), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(KEYINPUT60), .B(n1013), .ZN(n1024) );
  XNOR2_X1 U1101 ( .A(KEYINPUT127), .B(G5), .ZN(n1015) );
  XNOR2_X1 U1102 ( .A(n1015), .B(n1014), .ZN(n1022) );
  XNOR2_X1 U1103 ( .A(G1976), .B(G23), .ZN(n1017) );
  XNOR2_X1 U1104 ( .A(G1971), .B(G22), .ZN(n1016) );
  NOR2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1019) );
  XOR2_X1 U1106 ( .A(G1986), .B(G24), .Z(n1018) );
  NAND2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1108 ( .A(KEYINPUT58), .B(n1020), .ZN(n1021) );
  NOR2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1026) );
  XNOR2_X1 U1111 ( .A(G21), .B(G1966), .ZN(n1025) );
  NOR2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1113 ( .A(KEYINPUT61), .B(n1027), .Z(n1028) );
  NOR2_X1 U1114 ( .A1(G16), .A2(n1028), .ZN(n1029) );
  NOR2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1116 ( .A(n1031), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1117 ( .A(G311), .ZN(G150) );
  INV_X1 U1118 ( .A(G171), .ZN(G301) );
endmodule

