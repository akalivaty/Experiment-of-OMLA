

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755;

  AND2_X1 U372 ( .A1(n399), .A2(n599), .ZN(n379) );
  BUF_X1 U373 ( .A(n537), .Z(n554) );
  INV_X1 U374 ( .A(G953), .ZN(n744) );
  NOR2_X1 U375 ( .A1(n514), .A2(n530), .ZN(n707) );
  XNOR2_X2 U376 ( .A(n452), .B(n451), .ZN(n513) );
  OR2_X2 U377 ( .A1(n672), .A2(G902), .ZN(n452) );
  NOR2_X2 U378 ( .A1(n631), .A2(n520), .ZN(n712) );
  NOR2_X1 U379 ( .A1(n631), .A2(n632), .ZN(n588) );
  INV_X1 U380 ( .A(n542), .ZN(n705) );
  NOR2_X1 U381 ( .A1(n522), .A2(n521), .ZN(n523) );
  NAND2_X1 U382 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U383 ( .A1(n620), .A2(n728), .ZN(n671) );
  NAND2_X1 U384 ( .A1(n712), .A2(n549), .ZN(n411) );
  NAND2_X1 U385 ( .A1(n395), .A2(n393), .ZN(n603) );
  AND2_X1 U386 ( .A1(n397), .A2(n356), .ZN(n395) );
  XNOR2_X1 U387 ( .A(n523), .B(KEYINPUT40), .ZN(n754) );
  AND2_X1 U388 ( .A1(n532), .A2(n509), .ZN(n510) );
  NOR2_X1 U389 ( .A1(n652), .A2(n589), .ZN(n591) );
  AND2_X1 U390 ( .A1(n483), .A2(n482), .ZN(n532) );
  NOR2_X1 U391 ( .A1(n602), .A2(n525), .ZN(n526) );
  INV_X1 U392 ( .A(n579), .ZN(n349) );
  XNOR2_X1 U393 ( .A(n602), .B(KEYINPUT6), .ZN(n607) );
  XNOR2_X1 U394 ( .A(n390), .B(n359), .ZN(n565) );
  NAND2_X1 U395 ( .A1(n537), .A2(n643), .ZN(n390) );
  INV_X2 U396 ( .A(n513), .ZN(n350) );
  XNOR2_X1 U397 ( .A(n502), .B(n741), .ZN(n490) );
  XNOR2_X1 U398 ( .A(n740), .B(n733), .ZN(n502) );
  XNOR2_X1 U399 ( .A(G128), .B(KEYINPUT65), .ZN(n413) );
  XNOR2_X1 U400 ( .A(G110), .B(G107), .ZN(n484) );
  NOR2_X1 U401 ( .A1(n531), .A2(n530), .ZN(n578) );
  XNOR2_X1 U402 ( .A(n352), .B(n417), .ZN(n739) );
  XNOR2_X1 U403 ( .A(KEYINPUT70), .B(KEYINPUT10), .ZN(n417) );
  INV_X1 U404 ( .A(n350), .ZN(n602) );
  XNOR2_X1 U405 ( .A(n490), .B(n491), .ZN(n716) );
  NAND2_X1 U406 ( .A1(n685), .A2(n753), .ZN(n399) );
  XOR2_X1 U407 ( .A(KEYINPUT14), .B(KEYINPUT95), .Z(n476) );
  OR2_X1 U408 ( .A1(n370), .A2(n367), .ZN(n525) );
  INV_X1 U409 ( .A(KEYINPUT72), .ZN(n371) );
  XNOR2_X1 U410 ( .A(n429), .B(n388), .ZN(n531) );
  XNOR2_X1 U411 ( .A(n430), .B(n389), .ZN(n388) );
  XNOR2_X1 U412 ( .A(n434), .B(n433), .ZN(n435) );
  INV_X1 U413 ( .A(KEYINPUT7), .ZN(n433) );
  XNOR2_X1 U414 ( .A(G134), .B(G116), .ZN(n434) );
  XNOR2_X1 U415 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n438) );
  XNOR2_X1 U416 ( .A(n416), .B(G143), .ZN(n387) );
  XNOR2_X1 U417 ( .A(n739), .B(n418), .ZN(n469) );
  XNOR2_X1 U418 ( .A(n364), .B(n502), .ZN(n687) );
  XNOR2_X1 U419 ( .A(n734), .B(n501), .ZN(n364) );
  XNOR2_X1 U420 ( .A(n377), .B(n358), .ZN(n652) );
  NAND2_X1 U421 ( .A1(n588), .A2(n607), .ZN(n377) );
  OR2_X1 U422 ( .A1(n631), .A2(KEYINPUT113), .ZN(n396) );
  XNOR2_X1 U423 ( .A(n443), .B(G478), .ZN(n530) );
  NAND2_X1 U424 ( .A1(n723), .A2(n361), .ZN(n403) );
  NOR2_X1 U425 ( .A1(n402), .A2(n727), .ZN(n401) );
  NOR2_X1 U426 ( .A1(n357), .A2(G469), .ZN(n402) );
  INV_X1 U427 ( .A(G475), .ZN(n389) );
  INV_X1 U428 ( .A(n714), .ZN(n412) );
  NOR2_X1 U429 ( .A1(n712), .A2(n409), .ZN(n408) );
  NAND2_X1 U430 ( .A1(n412), .A2(KEYINPUT48), .ZN(n409) );
  XNOR2_X1 U431 ( .A(n414), .B(n444), .ZN(n740) );
  XNOR2_X1 U432 ( .A(n363), .B(n366), .ZN(n414) );
  INV_X1 U433 ( .A(KEYINPUT4), .ZN(n366) );
  XNOR2_X1 U434 ( .A(KEYINPUT64), .B(G146), .ZN(n363) );
  XNOR2_X1 U435 ( .A(KEYINPUT71), .B(G131), .ZN(n445) );
  AND2_X1 U436 ( .A1(n372), .A2(n629), .ZN(n515) );
  XNOR2_X1 U437 ( .A(G137), .B(G128), .ZN(n459) );
  XNOR2_X1 U438 ( .A(KEYINPUT23), .B(KEYINPUT99), .ZN(n461) );
  XNOR2_X1 U439 ( .A(n385), .B(KEYINPUT115), .ZN(n516) );
  NAND2_X1 U440 ( .A1(n607), .A2(n355), .ZN(n385) );
  OR2_X1 U441 ( .A1(n539), .A2(n561), .ZN(n542) );
  XNOR2_X1 U442 ( .A(n471), .B(n470), .ZN(n368) );
  INV_X1 U443 ( .A(n531), .ZN(n514) );
  NAND2_X1 U444 ( .A1(n349), .A2(n353), .ZN(n582) );
  XNOR2_X1 U445 ( .A(n497), .B(n496), .ZN(n734) );
  XNOR2_X1 U446 ( .A(n495), .B(n494), .ZN(n497) );
  XNOR2_X1 U447 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U448 ( .A(n469), .B(n387), .ZN(n428) );
  AND2_X1 U449 ( .A1(n660), .A2(n360), .ZN(n374) );
  XNOR2_X1 U450 ( .A(n570), .B(n569), .ZN(n710) );
  XNOR2_X1 U451 ( .A(KEYINPUT31), .B(KEYINPUT104), .ZN(n569) );
  NOR2_X1 U452 ( .A1(n404), .A2(n400), .ZN(n717) );
  NOR2_X1 U453 ( .A1(n723), .A2(n357), .ZN(n404) );
  NAND2_X1 U454 ( .A1(n403), .A2(n401), .ZN(n400) );
  AND2_X1 U455 ( .A1(n631), .A2(KEYINPUT113), .ZN(n351) );
  XOR2_X1 U456 ( .A(G125), .B(G140), .Z(n352) );
  XNOR2_X1 U457 ( .A(n413), .B(G143), .ZN(n444) );
  XNOR2_X1 U458 ( .A(n369), .B(n368), .ZN(n604) );
  INV_X1 U459 ( .A(n604), .ZN(n367) );
  AND2_X1 U460 ( .A1(n578), .A2(n629), .ZN(n353) );
  OR2_X1 U461 ( .A1(n564), .A2(n563), .ZN(n354) );
  AND2_X1 U462 ( .A1(n386), .A2(n707), .ZN(n355) );
  AND2_X1 U463 ( .A1(n396), .A2(n602), .ZN(n356) );
  XOR2_X1 U464 ( .A(n716), .B(n715), .Z(n357) );
  XOR2_X1 U465 ( .A(KEYINPUT33), .B(KEYINPUT74), .Z(n358) );
  XOR2_X1 U466 ( .A(n538), .B(KEYINPUT68), .Z(n359) );
  OR2_X1 U467 ( .A1(n642), .A2(n652), .ZN(n360) );
  AND2_X1 U468 ( .A1(n357), .A2(G469), .ZN(n361) );
  NAND2_X1 U469 ( .A1(n362), .A2(n616), .ZN(n398) );
  NAND2_X1 U470 ( .A1(n379), .A2(n378), .ZN(n362) );
  NAND2_X1 U471 ( .A1(n394), .A2(n600), .ZN(n393) );
  NAND2_X1 U472 ( .A1(n398), .A2(n617), .ZN(n619) );
  NOR2_X1 U473 ( .A1(n754), .A2(n755), .ZN(n529) );
  NAND2_X1 U474 ( .A1(n365), .A2(n571), .ZN(n539) );
  XNOR2_X1 U475 ( .A(n526), .B(KEYINPUT28), .ZN(n365) );
  NOR2_X1 U476 ( .A1(n679), .A2(G902), .ZN(n369) );
  XNOR2_X1 U477 ( .A(n515), .B(n371), .ZN(n370) );
  XNOR2_X1 U478 ( .A(n481), .B(KEYINPUT83), .ZN(n372) );
  XNOR2_X1 U479 ( .A(n373), .B(n662), .ZN(G75) );
  NAND2_X1 U480 ( .A1(n375), .A2(n374), .ZN(n373) );
  XNOR2_X1 U481 ( .A(n627), .B(n376), .ZN(n375) );
  INV_X1 U482 ( .A(KEYINPUT86), .ZN(n376) );
  XNOR2_X2 U483 ( .A(n512), .B(KEYINPUT1), .ZN(n631) );
  NAND2_X1 U484 ( .A1(n751), .A2(KEYINPUT91), .ZN(n378) );
  NAND2_X1 U485 ( .A1(n382), .A2(n380), .ZN(n557) );
  NAND2_X1 U486 ( .A1(n381), .A2(n408), .ZN(n380) );
  AND2_X1 U487 ( .A1(n548), .A2(n547), .ZN(n381) );
  NOR2_X2 U488 ( .A1(n545), .A2(n546), .ZN(n547) );
  NAND2_X1 U489 ( .A1(n383), .A2(n412), .ZN(n382) );
  NAND2_X1 U490 ( .A1(n384), .A2(n411), .ZN(n383) );
  NAND2_X1 U491 ( .A1(n410), .A2(n549), .ZN(n384) );
  INV_X1 U492 ( .A(n707), .ZN(n521) );
  INV_X1 U493 ( .A(n525), .ZN(n386) );
  INV_X1 U494 ( .A(n565), .ZN(n561) );
  XNOR2_X2 U495 ( .A(n507), .B(n506), .ZN(n537) );
  XNOR2_X2 U496 ( .A(n392), .B(n391), .ZN(n495) );
  XNOR2_X2 U497 ( .A(KEYINPUT3), .B(G119), .ZN(n391) );
  XNOR2_X2 U498 ( .A(G116), .B(G113), .ZN(n392) );
  AND2_X1 U499 ( .A1(n610), .A2(n631), .ZN(n601) );
  INV_X1 U500 ( .A(n610), .ZN(n394) );
  NAND2_X1 U501 ( .A1(n610), .A2(n351), .ZN(n397) );
  XNOR2_X2 U502 ( .A(n582), .B(n581), .ZN(n610) );
  INV_X1 U503 ( .A(n399), .ZN(n614) );
  AND2_X4 U504 ( .A1(n671), .A2(n670), .ZN(n723) );
  NAND2_X1 U505 ( .A1(n350), .A2(n643), .ZN(n407) );
  NAND2_X1 U506 ( .A1(n350), .A2(n405), .ZN(n457) );
  AND2_X1 U507 ( .A1(n406), .A2(n643), .ZN(n405) );
  INV_X1 U508 ( .A(n455), .ZN(n406) );
  NAND2_X1 U509 ( .A1(n407), .A2(n455), .ZN(n456) );
  NAND2_X1 U510 ( .A1(n548), .A2(n547), .ZN(n410) );
  NOR2_X2 U511 ( .A1(n690), .A2(n727), .ZN(n693) );
  NOR2_X2 U512 ( .A1(n721), .A2(n727), .ZN(n722) );
  XNOR2_X2 U513 ( .A(n568), .B(n567), .ZN(n579) );
  AND2_X1 U514 ( .A1(n743), .A2(n664), .ZN(n415) );
  XOR2_X1 U515 ( .A(n420), .B(n419), .Z(n416) );
  INV_X1 U516 ( .A(KEYINPUT80), .ZN(n485) );
  XNOR2_X1 U517 ( .A(n486), .B(n485), .ZN(n487) );
  INV_X1 U518 ( .A(KEYINPUT48), .ZN(n549) );
  XNOR2_X1 U519 ( .A(n496), .B(n487), .ZN(n488) );
  INV_X1 U520 ( .A(KEYINPUT88), .ZN(n558) );
  XNOR2_X1 U521 ( .A(n559), .B(n558), .ZN(n620) );
  INV_X1 U522 ( .A(KEYINPUT113), .ZN(n600) );
  INV_X1 U523 ( .A(KEYINPUT124), .ZN(n661) );
  INV_X1 U524 ( .A(KEYINPUT63), .ZN(n677) );
  INV_X1 U525 ( .A(KEYINPUT127), .ZN(n682) );
  INV_X1 U526 ( .A(G146), .ZN(n418) );
  XOR2_X1 U527 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n420) );
  XNOR2_X1 U528 ( .A(G104), .B(G122), .ZN(n419) );
  XNOR2_X1 U529 ( .A(G113), .B(n445), .ZN(n422) );
  NOR2_X1 U530 ( .A1(G953), .A2(G237), .ZN(n447) );
  NAND2_X1 U531 ( .A1(G214), .A2(n447), .ZN(n421) );
  XNOR2_X1 U532 ( .A(n422), .B(n421), .ZN(n426) );
  XOR2_X1 U533 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n424) );
  XNOR2_X1 U534 ( .A(KEYINPUT107), .B(KEYINPUT106), .ZN(n423) );
  XNOR2_X1 U535 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U536 ( .A(n426), .B(n425), .Z(n427) );
  XNOR2_X1 U537 ( .A(n428), .B(n427), .ZN(n718) );
  NOR2_X1 U538 ( .A1(G902), .A2(n718), .ZN(n429) );
  INV_X1 U539 ( .A(KEYINPUT13), .ZN(n430) );
  XOR2_X1 U540 ( .A(KEYINPUT9), .B(KEYINPUT110), .Z(n432) );
  XNOR2_X1 U541 ( .A(G107), .B(G122), .ZN(n431) );
  XNOR2_X1 U542 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U543 ( .A(n444), .B(n437), .Z(n441) );
  NAND2_X1 U544 ( .A1(n744), .A2(G234), .ZN(n439) );
  XNOR2_X1 U545 ( .A(n439), .B(n438), .ZN(n465) );
  NAND2_X1 U546 ( .A1(G217), .A2(n465), .ZN(n440) );
  XNOR2_X1 U547 ( .A(n441), .B(n440), .ZN(n725) );
  NOR2_X1 U548 ( .A1(G902), .A2(n725), .ZN(n442) );
  XNOR2_X1 U549 ( .A(n442), .B(KEYINPUT111), .ZN(n443) );
  AND2_X1 U550 ( .A1(n514), .A2(n530), .ZN(n709) );
  INV_X1 U551 ( .A(n709), .ZN(n511) );
  XOR2_X1 U552 ( .A(KEYINPUT118), .B(KEYINPUT30), .Z(n455) );
  INV_X1 U553 ( .A(G101), .ZN(n733) );
  XNOR2_X1 U554 ( .A(G137), .B(G134), .ZN(n446) );
  XNOR2_X1 U555 ( .A(n446), .B(n445), .ZN(n741) );
  NAND2_X1 U556 ( .A1(n447), .A2(G210), .ZN(n448) );
  XNOR2_X1 U557 ( .A(n448), .B(KEYINPUT5), .ZN(n449) );
  XNOR2_X1 U558 ( .A(n495), .B(n449), .ZN(n450) );
  XNOR2_X1 U559 ( .A(n490), .B(n450), .ZN(n672) );
  XNOR2_X1 U560 ( .A(KEYINPUT75), .B(G472), .ZN(n451) );
  INV_X1 U561 ( .A(G902), .ZN(n454) );
  INV_X1 U562 ( .A(G237), .ZN(n453) );
  NAND2_X1 U563 ( .A1(n454), .A2(n453), .ZN(n503) );
  NAND2_X1 U564 ( .A1(n503), .A2(G214), .ZN(n643) );
  NAND2_X1 U565 ( .A1(n457), .A2(n456), .ZN(n483) );
  XNOR2_X1 U566 ( .A(KEYINPUT15), .B(G902), .ZN(n666) );
  NAND2_X1 U567 ( .A1(G234), .A2(n666), .ZN(n458) );
  XNOR2_X1 U568 ( .A(KEYINPUT20), .B(n458), .ZN(n472) );
  AND2_X1 U569 ( .A1(n472), .A2(G217), .ZN(n471) );
  XNOR2_X1 U570 ( .A(KEYINPUT100), .B(KEYINPUT25), .ZN(n470) );
  XOR2_X1 U571 ( .A(G110), .B(G119), .Z(n460) );
  XNOR2_X1 U572 ( .A(n460), .B(n459), .ZN(n464) );
  XOR2_X1 U573 ( .A(KEYINPUT24), .B(KEYINPUT98), .Z(n462) );
  XNOR2_X1 U574 ( .A(n462), .B(n461), .ZN(n463) );
  XOR2_X1 U575 ( .A(n464), .B(n463), .Z(n467) );
  NAND2_X1 U576 ( .A1(G221), .A2(n465), .ZN(n466) );
  XNOR2_X1 U577 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U578 ( .A(n469), .B(n468), .ZN(n679) );
  NAND2_X1 U579 ( .A1(n472), .A2(G221), .ZN(n474) );
  XNOR2_X1 U580 ( .A(KEYINPUT101), .B(KEYINPUT21), .ZN(n473) );
  XNOR2_X1 U581 ( .A(n474), .B(n473), .ZN(n629) );
  NAND2_X1 U582 ( .A1(G237), .A2(G234), .ZN(n475) );
  XNOR2_X1 U583 ( .A(n476), .B(n475), .ZN(n477) );
  NAND2_X1 U584 ( .A1(G952), .A2(n477), .ZN(n658) );
  NOR2_X1 U585 ( .A1(n658), .A2(G953), .ZN(n564) );
  NAND2_X1 U586 ( .A1(G902), .A2(n477), .ZN(n562) );
  NOR2_X1 U587 ( .A1(G900), .A2(n562), .ZN(n478) );
  NAND2_X1 U588 ( .A1(G953), .A2(n478), .ZN(n479) );
  XOR2_X1 U589 ( .A(KEYINPUT114), .B(n479), .Z(n480) );
  NOR2_X1 U590 ( .A1(n564), .A2(n480), .ZN(n481) );
  AND2_X1 U591 ( .A1(n367), .A2(n515), .ZN(n482) );
  XNOR2_X1 U592 ( .A(n484), .B(G104), .ZN(n496) );
  NAND2_X1 U593 ( .A1(G227), .A2(n744), .ZN(n486) );
  XOR2_X1 U594 ( .A(n488), .B(KEYINPUT97), .Z(n489) );
  XNOR2_X1 U595 ( .A(n489), .B(G140), .ZN(n491) );
  NOR2_X1 U596 ( .A1(G902), .A2(n716), .ZN(n493) );
  XOR2_X1 U597 ( .A(KEYINPUT73), .B(G469), .Z(n492) );
  XNOR2_X1 U598 ( .A(n493), .B(n492), .ZN(n512) );
  INV_X1 U599 ( .A(n512), .ZN(n571) );
  XNOR2_X1 U600 ( .A(KEYINPUT16), .B(G122), .ZN(n494) );
  NAND2_X1 U601 ( .A1(n744), .A2(G224), .ZN(n498) );
  XNOR2_X1 U602 ( .A(n498), .B(G125), .ZN(n500) );
  XNOR2_X1 U603 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n499) );
  XNOR2_X1 U604 ( .A(n500), .B(n499), .ZN(n501) );
  NAND2_X1 U605 ( .A1(n687), .A2(n666), .ZN(n507) );
  NAND2_X1 U606 ( .A1(n503), .A2(G210), .ZN(n505) );
  INV_X1 U607 ( .A(KEYINPUT94), .ZN(n504) );
  XNOR2_X1 U608 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U609 ( .A(n554), .B(KEYINPUT38), .ZN(n508) );
  INV_X1 U610 ( .A(n508), .ZN(n644) );
  AND2_X1 U611 ( .A1(n571), .A2(n644), .ZN(n509) );
  XNOR2_X1 U612 ( .A(n510), .B(KEYINPUT39), .ZN(n522) );
  NOR2_X1 U613 ( .A1(n511), .A2(n522), .ZN(n714) );
  NAND2_X1 U614 ( .A1(n516), .A2(n643), .ZN(n550) );
  INV_X1 U615 ( .A(n554), .ZN(n517) );
  NOR2_X1 U616 ( .A1(n550), .A2(n517), .ZN(n519) );
  XOR2_X1 U617 ( .A(KEYINPUT36), .B(KEYINPUT92), .Z(n518) );
  XNOR2_X1 U618 ( .A(n519), .B(n518), .ZN(n520) );
  NAND2_X1 U619 ( .A1(n644), .A2(n643), .ZN(n647) );
  INV_X1 U620 ( .A(n578), .ZN(n646) );
  NOR2_X1 U621 ( .A1(n647), .A2(n646), .ZN(n524) );
  XNOR2_X1 U622 ( .A(n524), .B(KEYINPUT41), .ZN(n642) );
  NOR2_X1 U623 ( .A1(n642), .A2(n539), .ZN(n527) );
  XNOR2_X1 U624 ( .A(n527), .B(KEYINPUT42), .ZN(n755) );
  XNOR2_X1 U625 ( .A(KEYINPUT46), .B(KEYINPUT90), .ZN(n528) );
  XNOR2_X1 U626 ( .A(n529), .B(n528), .ZN(n548) );
  NAND2_X1 U627 ( .A1(n531), .A2(n530), .ZN(n592) );
  NAND2_X1 U628 ( .A1(n532), .A2(n571), .ZN(n533) );
  NOR2_X1 U629 ( .A1(n592), .A2(n533), .ZN(n534) );
  NAND2_X1 U630 ( .A1(n554), .A2(n534), .ZN(n684) );
  NOR2_X1 U631 ( .A1(n707), .A2(n709), .ZN(n648) );
  NAND2_X1 U632 ( .A1(n648), .A2(KEYINPUT47), .ZN(n535) );
  NAND2_X1 U633 ( .A1(n684), .A2(n535), .ZN(n536) );
  XOR2_X1 U634 ( .A(KEYINPUT84), .B(n536), .Z(n541) );
  XNOR2_X1 U635 ( .A(KEYINPUT79), .B(KEYINPUT19), .ZN(n538) );
  NAND2_X1 U636 ( .A1(n542), .A2(KEYINPUT47), .ZN(n540) );
  NAND2_X1 U637 ( .A1(n541), .A2(n540), .ZN(n546) );
  NOR2_X1 U638 ( .A1(n648), .A2(KEYINPUT47), .ZN(n543) );
  NAND2_X1 U639 ( .A1(n705), .A2(n543), .ZN(n544) );
  XOR2_X1 U640 ( .A(KEYINPUT78), .B(n544), .Z(n545) );
  XNOR2_X1 U641 ( .A(KEYINPUT116), .B(n550), .ZN(n552) );
  INV_X1 U642 ( .A(n631), .ZN(n551) );
  NOR2_X1 U643 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U644 ( .A(n553), .B(KEYINPUT43), .ZN(n555) );
  NOR2_X1 U645 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U646 ( .A(n556), .B(KEYINPUT117), .ZN(n752) );
  AND2_X2 U647 ( .A1(n557), .A2(n752), .ZN(n743) );
  NAND2_X1 U648 ( .A1(n743), .A2(KEYINPUT2), .ZN(n559) );
  NAND2_X1 U649 ( .A1(n367), .A2(n629), .ZN(n632) );
  NAND2_X1 U650 ( .A1(n588), .A2(n350), .ZN(n560) );
  XNOR2_X1 U651 ( .A(n560), .B(KEYINPUT103), .ZN(n639) );
  OR2_X1 U652 ( .A1(n744), .A2(G898), .ZN(n735) );
  NOR2_X1 U653 ( .A1(n562), .A2(n735), .ZN(n563) );
  NAND2_X1 U654 ( .A1(n565), .A2(n354), .ZN(n568) );
  INV_X1 U655 ( .A(KEYINPUT93), .ZN(n566) );
  XNOR2_X1 U656 ( .A(n566), .B(KEYINPUT0), .ZN(n567) );
  NAND2_X1 U657 ( .A1(n639), .A2(n349), .ZN(n570) );
  XNOR2_X1 U658 ( .A(n579), .B(KEYINPUT96), .ZN(n589) );
  NOR2_X1 U659 ( .A1(n350), .A2(n632), .ZN(n572) );
  NAND2_X1 U660 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U661 ( .A1(n589), .A2(n573), .ZN(n574) );
  XNOR2_X1 U662 ( .A(n574), .B(KEYINPUT102), .ZN(n698) );
  NOR2_X1 U663 ( .A1(n710), .A2(n698), .ZN(n575) );
  XNOR2_X1 U664 ( .A(KEYINPUT105), .B(n575), .ZN(n577) );
  INV_X1 U665 ( .A(n648), .ZN(n576) );
  NAND2_X1 U666 ( .A1(n577), .A2(n576), .ZN(n587) );
  XNOR2_X1 U667 ( .A(KEYINPUT77), .B(KEYINPUT22), .ZN(n580) );
  XNOR2_X1 U668 ( .A(n580), .B(KEYINPUT76), .ZN(n581) );
  INV_X1 U669 ( .A(KEYINPUT112), .ZN(n583) );
  XNOR2_X1 U670 ( .A(n604), .B(n583), .ZN(n628) );
  INV_X1 U671 ( .A(n628), .ZN(n584) );
  NOR2_X1 U672 ( .A1(n607), .A2(n584), .ZN(n585) );
  AND2_X1 U673 ( .A1(n601), .A2(n585), .ZN(n694) );
  INV_X1 U674 ( .A(n694), .ZN(n586) );
  NAND2_X1 U675 ( .A1(n587), .A2(n586), .ZN(n598) );
  XOR2_X1 U676 ( .A(KEYINPUT34), .B(KEYINPUT81), .Z(n590) );
  XNOR2_X1 U677 ( .A(n591), .B(n590), .ZN(n594) );
  INV_X1 U678 ( .A(n592), .ZN(n593) );
  NAND2_X1 U679 ( .A1(n594), .A2(n593), .ZN(n596) );
  INV_X1 U680 ( .A(KEYINPUT35), .ZN(n595) );
  XNOR2_X2 U681 ( .A(n596), .B(n595), .ZN(n751) );
  INV_X1 U682 ( .A(KEYINPUT44), .ZN(n599) );
  NOR2_X1 U683 ( .A1(n751), .A2(n599), .ZN(n597) );
  NOR2_X1 U684 ( .A1(n598), .A2(n597), .ZN(n617) );
  XNOR2_X1 U685 ( .A(n603), .B(KEYINPUT67), .ZN(n605) );
  NAND2_X1 U686 ( .A1(n605), .A2(n604), .ZN(n685) );
  OR2_X1 U687 ( .A1(n628), .A2(n631), .ZN(n606) );
  NOR2_X1 U688 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U689 ( .A(KEYINPUT82), .B(n608), .ZN(n609) );
  NAND2_X1 U690 ( .A1(n610), .A2(n609), .ZN(n612) );
  XNOR2_X1 U691 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n611) );
  XNOR2_X1 U692 ( .A(n612), .B(n611), .ZN(n753) );
  NOR2_X1 U693 ( .A1(KEYINPUT91), .A2(KEYINPUT44), .ZN(n613) );
  NAND2_X1 U694 ( .A1(n751), .A2(n613), .ZN(n615) );
  NAND2_X1 U695 ( .A1(n615), .A2(n614), .ZN(n616) );
  INV_X1 U696 ( .A(KEYINPUT45), .ZN(n618) );
  XNOR2_X2 U697 ( .A(n619), .B(n618), .ZN(n663) );
  INV_X1 U698 ( .A(n663), .ZN(n728) );
  INV_X1 U699 ( .A(n671), .ZN(n626) );
  INV_X1 U700 ( .A(KEYINPUT2), .ZN(n621) );
  NAND2_X1 U701 ( .A1(n663), .A2(n621), .ZN(n624) );
  NOR2_X1 U702 ( .A1(n743), .A2(KEYINPUT2), .ZN(n622) );
  XNOR2_X1 U703 ( .A(n622), .B(KEYINPUT85), .ZN(n623) );
  NAND2_X1 U704 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U705 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U706 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U707 ( .A(KEYINPUT49), .B(n630), .ZN(n636) );
  NAND2_X1 U708 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U709 ( .A(n633), .B(KEYINPUT122), .ZN(n634) );
  XNOR2_X1 U710 ( .A(KEYINPUT50), .B(n634), .ZN(n635) );
  NAND2_X1 U711 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U712 ( .A1(n350), .A2(n637), .ZN(n638) );
  NOR2_X1 U713 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U714 ( .A(KEYINPUT51), .B(n640), .Z(n641) );
  NOR2_X1 U715 ( .A1(n642), .A2(n641), .ZN(n654) );
  NOR2_X1 U716 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U717 ( .A1(n646), .A2(n645), .ZN(n650) );
  NOR2_X1 U718 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U719 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U720 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U721 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U722 ( .A(n655), .B(KEYINPUT123), .Z(n656) );
  XNOR2_X1 U723 ( .A(KEYINPUT52), .B(n656), .ZN(n657) );
  NOR2_X1 U724 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U725 ( .A1(G953), .A2(n659), .ZN(n660) );
  XNOR2_X1 U726 ( .A(n661), .B(KEYINPUT53), .ZN(n662) );
  INV_X1 U727 ( .A(n663), .ZN(n665) );
  INV_X1 U728 ( .A(n666), .ZN(n664) );
  NAND2_X1 U729 ( .A1(n665), .A2(n415), .ZN(n669) );
  XNOR2_X1 U730 ( .A(n666), .B(KEYINPUT87), .ZN(n667) );
  NAND2_X1 U731 ( .A1(n667), .A2(KEYINPUT2), .ZN(n668) );
  NAND2_X1 U732 ( .A1(n723), .A2(G472), .ZN(n674) );
  XNOR2_X1 U733 ( .A(n672), .B(KEYINPUT62), .ZN(n673) );
  XNOR2_X1 U734 ( .A(n674), .B(n673), .ZN(n676) );
  INV_X1 U735 ( .A(G952), .ZN(n675) );
  AND2_X1 U736 ( .A1(n675), .A2(G953), .ZN(n727) );
  NOR2_X2 U737 ( .A1(n676), .A2(n727), .ZN(n678) );
  XNOR2_X1 U738 ( .A(n678), .B(n677), .ZN(G57) );
  NAND2_X1 U739 ( .A1(n723), .A2(G217), .ZN(n680) );
  XNOR2_X1 U740 ( .A(n680), .B(n679), .ZN(n681) );
  NOR2_X2 U741 ( .A1(n681), .A2(n727), .ZN(n683) );
  XNOR2_X1 U742 ( .A(n683), .B(n682), .ZN(G66) );
  XNOR2_X1 U743 ( .A(n684), .B(G143), .ZN(G45) );
  XNOR2_X1 U744 ( .A(n685), .B(G110), .ZN(G12) );
  NAND2_X1 U745 ( .A1(n723), .A2(G210), .ZN(n689) );
  XNOR2_X1 U746 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n686) );
  XNOR2_X1 U747 ( .A(n687), .B(n686), .ZN(n688) );
  XNOR2_X1 U748 ( .A(n689), .B(n688), .ZN(n690) );
  XNOR2_X1 U749 ( .A(KEYINPUT125), .B(KEYINPUT56), .ZN(n691) );
  XNOR2_X1 U750 ( .A(n691), .B(KEYINPUT89), .ZN(n692) );
  XNOR2_X1 U751 ( .A(n693), .B(n692), .ZN(G51) );
  XNOR2_X1 U752 ( .A(G101), .B(n694), .ZN(n695) );
  XNOR2_X1 U753 ( .A(n695), .B(KEYINPUT119), .ZN(G3) );
  NAND2_X1 U754 ( .A1(n698), .A2(n707), .ZN(n696) );
  XNOR2_X1 U755 ( .A(n696), .B(KEYINPUT120), .ZN(n697) );
  XNOR2_X1 U756 ( .A(G104), .B(n697), .ZN(G6) );
  XOR2_X1 U757 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n700) );
  NAND2_X1 U758 ( .A1(n709), .A2(n698), .ZN(n699) );
  XNOR2_X1 U759 ( .A(n700), .B(n699), .ZN(n701) );
  XNOR2_X1 U760 ( .A(G107), .B(n701), .ZN(G9) );
  XOR2_X1 U761 ( .A(KEYINPUT29), .B(KEYINPUT121), .Z(n703) );
  NAND2_X1 U762 ( .A1(n705), .A2(n709), .ZN(n702) );
  XNOR2_X1 U763 ( .A(n703), .B(n702), .ZN(n704) );
  XOR2_X1 U764 ( .A(G128), .B(n704), .Z(G30) );
  NAND2_X1 U765 ( .A1(n705), .A2(n707), .ZN(n706) );
  XNOR2_X1 U766 ( .A(n706), .B(G146), .ZN(G48) );
  NAND2_X1 U767 ( .A1(n710), .A2(n707), .ZN(n708) );
  XNOR2_X1 U768 ( .A(n708), .B(G113), .ZN(G15) );
  NAND2_X1 U769 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U770 ( .A(n711), .B(G116), .ZN(G18) );
  XNOR2_X1 U771 ( .A(G125), .B(n712), .ZN(n713) );
  XNOR2_X1 U772 ( .A(n713), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U773 ( .A(G134), .B(n714), .Z(G36) );
  XOR2_X1 U774 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n715) );
  XNOR2_X1 U775 ( .A(KEYINPUT126), .B(n717), .ZN(G54) );
  NAND2_X1 U776 ( .A1(n723), .A2(G475), .ZN(n720) );
  XOR2_X1 U777 ( .A(n718), .B(KEYINPUT59), .Z(n719) );
  XNOR2_X1 U778 ( .A(n720), .B(n719), .ZN(n721) );
  XNOR2_X1 U779 ( .A(n722), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U780 ( .A1(n723), .A2(G478), .ZN(n724) );
  XNOR2_X1 U781 ( .A(n725), .B(n724), .ZN(n726) );
  NOR2_X1 U782 ( .A1(n727), .A2(n726), .ZN(G63) );
  NAND2_X1 U783 ( .A1(n728), .A2(n744), .ZN(n732) );
  NAND2_X1 U784 ( .A1(G953), .A2(G224), .ZN(n729) );
  XNOR2_X1 U785 ( .A(KEYINPUT61), .B(n729), .ZN(n730) );
  NAND2_X1 U786 ( .A1(n730), .A2(G898), .ZN(n731) );
  NAND2_X1 U787 ( .A1(n732), .A2(n731), .ZN(n738) );
  XNOR2_X1 U788 ( .A(n734), .B(n733), .ZN(n736) );
  NAND2_X1 U789 ( .A1(n736), .A2(n735), .ZN(n737) );
  XOR2_X1 U790 ( .A(n738), .B(n737), .Z(G69) );
  XNOR2_X1 U791 ( .A(n740), .B(n739), .ZN(n742) );
  XOR2_X1 U792 ( .A(n742), .B(n741), .Z(n746) );
  XOR2_X1 U793 ( .A(n746), .B(n743), .Z(n745) );
  NAND2_X1 U794 ( .A1(n745), .A2(n744), .ZN(n750) );
  XNOR2_X1 U795 ( .A(G227), .B(n746), .ZN(n747) );
  NAND2_X1 U796 ( .A1(n747), .A2(G900), .ZN(n748) );
  NAND2_X1 U797 ( .A1(n748), .A2(G953), .ZN(n749) );
  NAND2_X1 U798 ( .A1(n750), .A2(n749), .ZN(G72) );
  XNOR2_X1 U799 ( .A(G122), .B(n751), .ZN(G24) );
  XNOR2_X1 U800 ( .A(n752), .B(G140), .ZN(G42) );
  XNOR2_X1 U801 ( .A(G119), .B(n753), .ZN(G21) );
  XOR2_X1 U802 ( .A(n754), .B(G131), .Z(G33) );
  XOR2_X1 U803 ( .A(n755), .B(G137), .Z(G39) );
endmodule

