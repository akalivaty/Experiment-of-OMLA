//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 1 0 1 1 1 1 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 1 1 1 0 0 0 1 0 0 0 0 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:59 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n562, new_n564, new_n565,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n629, new_n630,
    new_n631, new_n634, new_n635, new_n637, new_n638, new_n639, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1243, new_n1244, new_n1245;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI21_X1  g030(.A(KEYINPUT66), .B1(new_n451), .B2(G2106), .ZN(new_n456));
  AOI21_X1  g031(.A(new_n456), .B1(G567), .B2(new_n453), .ZN(new_n457));
  NAND3_X1  g032(.A1(new_n451), .A2(KEYINPUT66), .A3(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT67), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n470));
  AND3_X1   g045(.A1(new_n467), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n470), .B1(new_n467), .B2(new_n469), .ZN(new_n472));
  OAI21_X1  g047(.A(G125), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n465), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n467), .A2(new_n469), .ZN(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT67), .B(G2105), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G137), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n466), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G101), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n475), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT69), .ZN(G160));
  OAI221_X1 g059(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n465), .C2(G112), .ZN(new_n485));
  OAI21_X1  g060(.A(KEYINPUT70), .B1(new_n476), .B2(G2105), .ZN(new_n486));
  XNOR2_X1  g061(.A(KEYINPUT3), .B(G2104), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT70), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n487), .A2(new_n488), .A3(new_n461), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G136), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n485), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(KEYINPUT71), .B1(new_n476), .B2(new_n465), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT71), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n487), .A2(new_n477), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n493), .B1(G124), .B2(new_n497), .ZN(G162));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n465), .B(new_n500), .C1(new_n471), .C2(new_n472), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n465), .A2(new_n487), .A3(G138), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(G114), .A2(G2104), .ZN(new_n505));
  INV_X1    g080(.A(G126), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n505), .B1(new_n476), .B2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G2105), .B1(G102), .B2(new_n480), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n513), .A2(KEYINPUT5), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(KEYINPUT6), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G651), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n515), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  INV_X1    g099(.A(G50), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n519), .A2(new_n521), .A3(G543), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n523), .A2(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n518), .A2(new_n527), .ZN(G166));
  INV_X1    g103(.A(KEYINPUT72), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n529), .B1(new_n512), .B2(new_n514), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n513), .A2(KEYINPUT5), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n511), .A2(G543), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n531), .A2(new_n532), .A3(KEYINPUT72), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n534), .A2(G63), .A3(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n531), .A2(new_n532), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n519), .A2(new_n521), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n526), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n538), .A2(G89), .B1(new_n539), .B2(G51), .ZN(new_n540));
  XOR2_X1   g115(.A(KEYINPUT73), .B(KEYINPUT7), .Z(new_n541));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n541), .B(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n535), .A2(new_n540), .A3(new_n543), .ZN(G286));
  INV_X1    g119(.A(G286), .ZN(G168));
  AOI22_X1  g120(.A1(new_n534), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n546), .A2(new_n517), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n538), .A2(G90), .B1(new_n539), .B2(G52), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n547), .A2(new_n549), .ZN(G171));
  AOI22_X1  g125(.A1(new_n538), .A2(G81), .B1(new_n539), .B2(G43), .ZN(new_n551));
  AND3_X1   g126(.A1(new_n531), .A2(new_n532), .A3(KEYINPUT72), .ZN(new_n552));
  AOI21_X1  g127(.A(KEYINPUT72), .B1(new_n531), .B2(new_n532), .ZN(new_n553));
  OAI21_X1  g128(.A(G56), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(G68), .A2(G543), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n554), .A2(KEYINPUT74), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G651), .ZN(new_n557));
  AOI21_X1  g132(.A(KEYINPUT74), .B1(new_n554), .B2(new_n555), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n551), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  AND3_X1   g136(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G36), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n562), .A2(new_n565), .ZN(G188));
  INV_X1    g141(.A(KEYINPUT75), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n539), .A2(new_n567), .A3(G53), .ZN(new_n568));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT75), .B1(new_n526), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(KEYINPUT9), .A3(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT9), .ZN(new_n572));
  OAI211_X1 g147(.A(KEYINPUT75), .B(new_n572), .C1(new_n526), .C2(new_n569), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n538), .A2(G91), .ZN(new_n574));
  NAND2_X1  g149(.A1(G78), .A2(G543), .ZN(new_n575));
  XOR2_X1   g150(.A(new_n575), .B(KEYINPUT76), .Z(new_n576));
  AND3_X1   g151(.A1(new_n531), .A2(new_n532), .A3(G65), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n571), .A2(new_n573), .A3(new_n574), .A4(new_n578), .ZN(G299));
  INV_X1    g154(.A(G171), .ZN(G301));
  INV_X1    g155(.A(G166), .ZN(G303));
  AOI22_X1  g156(.A1(new_n538), .A2(G87), .B1(new_n539), .B2(G49), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT77), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n583), .B(G651), .C1(new_n534), .C2(G74), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(G74), .A2(G651), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(new_n587));
  AOI211_X1 g162(.A(new_n583), .B(new_n587), .C1(new_n534), .C2(G651), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n582), .B1(new_n585), .B2(new_n588), .ZN(G288));
  NAND2_X1  g164(.A1(new_n515), .A2(G61), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(KEYINPUT78), .B1(G73), .B2(G543), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT78), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n515), .A2(new_n592), .A3(G61), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n517), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(G86), .ZN(new_n595));
  INV_X1    g170(.A(G48), .ZN(new_n596));
  OAI22_X1  g171(.A1(new_n523), .A2(new_n595), .B1(new_n596), .B2(new_n526), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(G305));
  INV_X1    g174(.A(G60), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n600), .B1(new_n530), .B2(new_n533), .ZN(new_n601));
  NAND2_X1  g176(.A1(G72), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(G651), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  XOR2_X1   g179(.A(KEYINPUT79), .B(G47), .Z(new_n605));
  NAND2_X1  g180(.A1(new_n539), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n515), .A2(new_n522), .A3(G85), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n606), .A2(new_n607), .A3(KEYINPUT80), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g184(.A(KEYINPUT80), .B1(new_n606), .B2(new_n607), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n604), .B1(new_n609), .B2(new_n610), .ZN(G290));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  INV_X1    g187(.A(G92), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n523), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n538), .A2(KEYINPUT10), .A3(G92), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(G79), .ZN(new_n617));
  OR3_X1    g192(.A1(new_n617), .A2(new_n513), .A3(KEYINPUT81), .ZN(new_n618));
  OAI21_X1  g193(.A(KEYINPUT81), .B1(new_n617), .B2(new_n513), .ZN(new_n619));
  INV_X1    g194(.A(G66), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n618), .B(new_n619), .C1(new_n620), .C2(new_n536), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n621), .A2(G651), .B1(new_n539), .B2(G54), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n616), .A2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(G868), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G171), .B2(new_n624), .ZN(G284));
  OAI21_X1  g201(.A(new_n625), .B1(G171), .B2(new_n624), .ZN(G321));
  NAND2_X1  g202(.A1(G286), .A2(G868), .ZN(new_n628));
  INV_X1    g203(.A(new_n571), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n578), .A2(new_n574), .A3(new_n573), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n628), .B1(new_n631), .B2(G868), .ZN(G297));
  OAI21_X1  g207(.A(new_n628), .B1(new_n631), .B2(G868), .ZN(G280));
  INV_X1    g208(.A(new_n623), .ZN(new_n634));
  INV_X1    g209(.A(G559), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n634), .B1(new_n635), .B2(G860), .ZN(G148));
  NAND2_X1  g211(.A1(new_n559), .A2(new_n624), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n623), .A2(G559), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n637), .B1(new_n624), .B2(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT82), .ZN(G323));
  XNOR2_X1  g215(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g216(.A1(new_n476), .A2(KEYINPUT68), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n487), .A2(new_n470), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(new_n480), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT12), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT13), .Z(new_n647));
  OR2_X1    g222(.A1(new_n647), .A2(G2100), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(G2100), .ZN(new_n649));
  OAI221_X1 g224(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n465), .C2(G111), .ZN(new_n650));
  INV_X1    g225(.A(G135), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n650), .B1(new_n491), .B2(new_n651), .ZN(new_n652));
  AND2_X1   g227(.A1(new_n497), .A2(G123), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2096), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n648), .A2(new_n649), .A3(new_n655), .ZN(G156));
  XOR2_X1   g231(.A(G2443), .B(G2446), .Z(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2451), .B(G2454), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT14), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT15), .B(G2435), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2438), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2427), .B(G2430), .ZN(new_n666));
  INV_X1    g241(.A(KEYINPUT83), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n663), .B1(new_n665), .B2(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT84), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n670), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n665), .A2(new_n668), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n662), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  AOI211_X1 g251(.A(new_n674), .B(new_n661), .C1(new_n671), .C2(new_n672), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n658), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n672), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n669), .A2(new_n670), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n675), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(new_n661), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n673), .A2(new_n675), .A3(new_n662), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n682), .A2(new_n657), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1341), .B(G1348), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n678), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n686), .A2(G14), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n678), .A2(new_n684), .ZN(new_n688));
  INV_X1    g263(.A(new_n685), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n687), .A2(new_n690), .ZN(G401));
  XOR2_X1   g266(.A(G2084), .B(G2090), .Z(new_n692));
  XNOR2_X1  g267(.A(G2067), .B(G2678), .ZN(new_n693));
  XNOR2_X1  g268(.A(G2072), .B(G2078), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT18), .Z(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT86), .B(KEYINPUT17), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n694), .B(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n693), .ZN(new_n699));
  INV_X1    g274(.A(new_n694), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n692), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n699), .A2(new_n692), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n698), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n699), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n696), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(G2096), .B(G2100), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(G227));
  XOR2_X1   g282(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT88), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G1981), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(G1971), .B(G1976), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT19), .ZN(new_n713));
  XNOR2_X1  g288(.A(G1956), .B(G2474), .ZN(new_n714));
  XNOR2_X1  g289(.A(G1961), .B(G1966), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  OR3_X1    g291(.A1(new_n713), .A2(KEYINPUT87), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(KEYINPUT87), .B1(new_n713), .B2(new_n716), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n717), .A2(KEYINPUT20), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n714), .A2(new_n715), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  MUX2_X1   g296(.A(new_n720), .B(new_n721), .S(new_n713), .Z(new_n722));
  NAND2_X1  g297(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(KEYINPUT20), .B1(new_n717), .B2(new_n718), .ZN(new_n724));
  OR3_X1    g299(.A1(new_n723), .A2(G1991), .A3(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(G1991), .B1(new_n723), .B2(new_n724), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n725), .A2(G1996), .A3(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(G1996), .B1(new_n725), .B2(new_n726), .ZN(new_n729));
  NOR3_X1   g304(.A1(new_n728), .A2(new_n729), .A3(G1986), .ZN(new_n730));
  INV_X1    g305(.A(G1986), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n725), .A2(new_n726), .ZN(new_n732));
  INV_X1    g307(.A(G1996), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n731), .B1(new_n734), .B2(new_n727), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n711), .B1(new_n730), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g311(.A(G1986), .B1(new_n728), .B2(new_n729), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n734), .A2(new_n731), .A3(new_n727), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n737), .A2(new_n738), .A3(new_n710), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n736), .A2(new_n739), .ZN(G229));
  NOR2_X1   g315(.A1(G16), .A2(G23), .ZN(new_n741));
  INV_X1    g316(.A(new_n582), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n534), .A2(G651), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n743), .A2(KEYINPUT77), .A3(new_n586), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n742), .B1(new_n744), .B2(new_n584), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n741), .B1(new_n745), .B2(G16), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT33), .B(G1976), .Z(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(G16), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G22), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G166), .B2(new_n749), .ZN(new_n751));
  INV_X1    g326(.A(G1971), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n749), .A2(G6), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n598), .B2(new_n749), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT32), .B(G1981), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n753), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  AOI211_X1 g332(.A(new_n748), .B(new_n757), .C1(new_n755), .C2(new_n756), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT91), .B(KEYINPUT34), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  INV_X1    g336(.A(G29), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(G25), .ZN(new_n763));
  OAI21_X1  g338(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n764));
  INV_X1    g339(.A(G107), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n764), .B1(new_n477), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n497), .B2(G119), .ZN(new_n767));
  AND3_X1   g342(.A1(new_n490), .A2(KEYINPUT89), .A3(G131), .ZN(new_n768));
  AOI21_X1  g343(.A(KEYINPUT89), .B1(new_n490), .B2(G131), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n763), .B1(new_n771), .B2(new_n762), .ZN(new_n772));
  XOR2_X1   g347(.A(KEYINPUT35), .B(G1991), .Z(new_n773));
  XOR2_X1   g348(.A(new_n772), .B(new_n773), .Z(new_n774));
  INV_X1    g349(.A(G24), .ZN(new_n775));
  OAI21_X1  g350(.A(KEYINPUT90), .B1(new_n775), .B2(G16), .ZN(new_n776));
  OR3_X1    g351(.A1(new_n775), .A2(KEYINPUT90), .A3(G16), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n606), .A2(new_n607), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT80), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n534), .A2(G60), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(new_n602), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n780), .A2(new_n608), .B1(new_n782), .B2(G651), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n776), .B(new_n777), .C1(new_n783), .C2(new_n749), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G1986), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n774), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n760), .A2(new_n761), .A3(new_n786), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT36), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n762), .A2(G33), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n644), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n790), .A2(new_n465), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT94), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT25), .Z(new_n794));
  INV_X1    g369(.A(G139), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(new_n491), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n789), .B1(new_n797), .B2(new_n762), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(G2072), .Z(new_n799));
  NOR2_X1   g374(.A1(G164), .A2(new_n762), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G27), .B2(new_n762), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(G168), .A2(G16), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G16), .B2(G21), .ZN(new_n804));
  INV_X1    g379(.A(G1966), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n802), .A2(G2078), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n805), .B2(new_n804), .ZN(new_n807));
  NOR2_X1   g382(.A1(G4), .A2(G16), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT92), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n623), .B2(new_n749), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G1348), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT31), .B(G11), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT99), .ZN(new_n813));
  INV_X1    g388(.A(G28), .ZN(new_n814));
  OR3_X1    g389(.A1(new_n813), .A2(new_n814), .A3(KEYINPUT30), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n813), .B1(new_n814), .B2(KEYINPUT30), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT100), .ZN(new_n817));
  AOI21_X1  g392(.A(G29), .B1(new_n814), .B2(KEYINPUT30), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n815), .B(new_n816), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n818), .A2(new_n817), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n812), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(new_n654), .B2(G29), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n811), .B(new_n822), .C1(new_n802), .C2(G2078), .ZN(new_n823));
  NOR2_X1   g398(.A1(G5), .A2(G16), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(G171), .B2(G16), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G1961), .ZN(new_n826));
  NOR3_X1   g401(.A1(new_n807), .A2(new_n823), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n749), .A2(G19), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n560), .B2(new_n749), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(G1341), .ZN(new_n830));
  INV_X1    g405(.A(G1956), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n749), .A2(G20), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(G299), .A2(G16), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n833), .B1(new_n834), .B2(KEYINPUT23), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(KEYINPUT23), .B2(new_n833), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n830), .B1(new_n831), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n799), .A2(new_n827), .A3(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT26), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(KEYINPUT96), .B1(new_n480), .B2(G105), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n461), .A2(G2104), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT96), .ZN(new_n844));
  INV_X1    g419(.A(G105), .ZN(new_n845));
  NOR3_X1   g420(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n841), .B1(new_n842), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n847), .B1(G141), .B2(new_n490), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n497), .A2(G129), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT97), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n850), .B1(new_n848), .B2(new_n849), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(G29), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT98), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n856), .B1(G29), .B2(G32), .ZN(new_n857));
  XNOR2_X1  g432(.A(KEYINPUT27), .B(G1996), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n836), .A2(new_n831), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n762), .A2(G35), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(G162), .B2(new_n762), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT29), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n863), .A2(G2090), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT101), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n860), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n866), .B1(new_n865), .B2(new_n864), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT28), .ZN(new_n868));
  AND2_X1   g443(.A1(new_n762), .A2(G26), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n490), .A2(G140), .ZN(new_n870));
  OAI221_X1 g445(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n465), .C2(G116), .ZN(new_n871));
  AND2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n497), .A2(G128), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI211_X1 g449(.A(new_n868), .B(new_n869), .C1(new_n874), .C2(G29), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n875), .B1(new_n868), .B2(new_n869), .ZN(new_n876));
  XNOR2_X1  g451(.A(KEYINPUT93), .B(G2067), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n863), .A2(G2090), .ZN(new_n879));
  INV_X1    g454(.A(G34), .ZN(new_n880));
  AOI21_X1  g455(.A(G29), .B1(new_n880), .B2(KEYINPUT24), .ZN(new_n881));
  OAI22_X1  g456(.A1(new_n881), .A2(KEYINPUT95), .B1(KEYINPUT24), .B2(new_n880), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n882), .B1(KEYINPUT95), .B2(new_n881), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n883), .B1(G160), .B2(G29), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(G2084), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n884), .A2(G2084), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n878), .A2(new_n879), .A3(new_n885), .A4(new_n886), .ZN(new_n887));
  NOR4_X1   g462(.A1(new_n838), .A2(new_n859), .A3(new_n867), .A4(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n788), .A2(new_n888), .ZN(G150));
  INV_X1    g464(.A(G150), .ZN(G311));
  INV_X1    g465(.A(G67), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n891), .B1(new_n530), .B2(new_n533), .ZN(new_n892));
  NAND2_X1  g467(.A1(G80), .A2(G543), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(G651), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  AOI22_X1  g470(.A1(new_n538), .A2(G93), .B1(new_n539), .B2(G55), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(G860), .ZN(new_n898));
  XOR2_X1   g473(.A(new_n898), .B(KEYINPUT37), .Z(new_n899));
  NAND2_X1  g474(.A1(new_n634), .A2(G559), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT39), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT104), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(KEYINPUT38), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n895), .A2(KEYINPUT102), .A3(new_n896), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT103), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n895), .A2(KEYINPUT102), .A3(new_n906), .A4(new_n896), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT102), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n897), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n559), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n905), .A2(new_n559), .A3(new_n907), .A4(new_n910), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n903), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(G860), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(new_n903), .B2(new_n914), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n899), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n918), .B(new_n919), .ZN(G145));
  OAI21_X1  g495(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n921));
  INV_X1    g496(.A(G118), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n921), .B1(new_n477), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n923), .B1(new_n490), .B2(G142), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n497), .A2(G130), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n771), .A2(new_n646), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n771), .A2(new_n646), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n770), .B(new_n646), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n931), .A2(new_n925), .A3(new_n924), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n874), .A2(new_n509), .ZN(new_n934));
  NAND3_X1  g509(.A1(G164), .A2(new_n873), .A3(new_n872), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n854), .ZN(new_n937));
  INV_X1    g512(.A(new_n853), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(new_n851), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n939), .A2(new_n934), .A3(new_n935), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n797), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n797), .A2(new_n937), .A3(new_n940), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n933), .A2(new_n943), .A3(KEYINPUT106), .A4(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n654), .ZN(new_n946));
  XNOR2_X1  g521(.A(G160), .B(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(G162), .ZN(new_n948));
  INV_X1    g523(.A(G162), .ZN(new_n949));
  AND2_X1   g524(.A1(G160), .A2(new_n654), .ZN(new_n950));
  NOR2_X1   g525(.A1(G160), .A2(new_n654), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n948), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n930), .A2(new_n932), .A3(KEYINPUT106), .ZN(new_n954));
  INV_X1    g529(.A(new_n944), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n797), .B1(new_n937), .B2(new_n940), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n945), .A2(new_n953), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n933), .B1(new_n955), .B2(new_n956), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n930), .A2(new_n932), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n943), .A2(new_n960), .A3(new_n944), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n948), .A2(new_n952), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n959), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G37), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n958), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  XOR2_X1   g540(.A(new_n965), .B(KEYINPUT40), .Z(G395));
  NAND2_X1  g541(.A1(new_n897), .A2(new_n624), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n914), .B(new_n638), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n631), .A2(new_n623), .ZN(new_n969));
  NAND3_X1  g544(.A1(G299), .A2(new_n616), .A3(new_n622), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n969), .A2(new_n970), .A3(KEYINPUT41), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT41), .B1(new_n969), .B2(new_n970), .ZN(new_n972));
  OAI21_X1  g547(.A(KEYINPUT107), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT107), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n969), .A2(new_n970), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT41), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n973), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n968), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n975), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n979), .B1(new_n980), .B2(new_n968), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n598), .A2(G303), .ZN(new_n982));
  OAI21_X1  g557(.A(G166), .B1(new_n594), .B2(new_n597), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(G288), .A2(new_n783), .ZN(new_n985));
  NAND2_X1  g560(.A1(G290), .A2(new_n745), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n985), .A2(KEYINPUT108), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT108), .B1(new_n985), .B2(new_n986), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n984), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n985), .A2(KEYINPUT108), .A3(new_n986), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n982), .A2(new_n983), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n993), .B(KEYINPUT42), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n981), .B(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n967), .B1(new_n995), .B2(new_n624), .ZN(G295));
  OAI21_X1  g571(.A(new_n967), .B1(new_n995), .B2(new_n624), .ZN(G331));
  OAI21_X1  g572(.A(G168), .B1(new_n547), .B2(new_n549), .ZN(new_n998));
  OAI211_X1 g573(.A(G286), .B(new_n548), .C1(new_n517), .C2(new_n546), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  AND4_X1   g576(.A1(new_n559), .A2(new_n905), .A3(new_n907), .A4(new_n910), .ZN(new_n1002));
  AOI22_X1  g577(.A1(new_n907), .A2(new_n905), .B1(new_n559), .B2(new_n910), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1001), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n912), .A2(new_n913), .A3(new_n1000), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1004), .A2(KEYINPUT110), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT110), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n912), .A2(new_n1007), .A3(new_n913), .A4(new_n1000), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n1006), .A2(new_n978), .A3(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1004), .A2(KEYINPUT111), .A3(new_n1005), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT111), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n914), .A2(new_n1011), .A3(new_n1001), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n980), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1009), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(G37), .B1(new_n1014), .B2(new_n993), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT43), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT108), .ZN(new_n1017));
  NOR2_X1   g592(.A1(G288), .A2(new_n783), .ZN(new_n1018));
  NOR2_X1   g593(.A1(G290), .A2(new_n745), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n991), .B1(new_n1020), .B2(new_n990), .ZN(new_n1021));
  INV_X1    g596(.A(new_n992), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n1021), .A2(new_n1022), .A3(KEYINPUT112), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1024), .B1(new_n989), .B2(new_n992), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1026), .B1(new_n1009), .B2(new_n1013), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1015), .A2(new_n1016), .A3(new_n1027), .ZN(new_n1028));
  OR2_X1    g603(.A1(new_n971), .A2(new_n972), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n1010), .A2(new_n1029), .A3(new_n1012), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n980), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1026), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n1015), .A2(new_n1032), .ZN(new_n1033));
  OAI211_X1 g608(.A(KEYINPUT44), .B(new_n1028), .C1(new_n1033), .C2(new_n1016), .ZN(new_n1034));
  XNOR2_X1  g609(.A(KEYINPUT109), .B(KEYINPUT44), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1016), .B1(new_n1015), .B2(new_n1027), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1006), .A2(new_n978), .A3(new_n1008), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n993), .B(new_n1037), .C1(new_n1038), .C2(new_n980), .ZN(new_n1039));
  AND4_X1   g614(.A1(new_n1016), .A2(new_n1032), .A3(new_n964), .A4(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1035), .B1(new_n1036), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1034), .A2(new_n1041), .ZN(G397));
  XNOR2_X1  g617(.A(KEYINPUT113), .B(G1384), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT45), .B1(new_n509), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G40), .ZN(new_n1045));
  NOR3_X1   g620(.A1(new_n475), .A2(new_n482), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1047), .B(KEYINPUT114), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1047), .A2(G1996), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT46), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1049), .B1(KEYINPUT125), .B2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1050), .A2(KEYINPUT125), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1052), .B1(new_n1047), .B2(G1996), .ZN(new_n1053));
  AOI22_X1  g628(.A1(new_n1048), .A2(new_n939), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n874), .A2(G2067), .ZN(new_n1055));
  INV_X1    g630(.A(G2067), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n872), .A2(new_n1056), .A3(new_n873), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n1048), .A2(new_n1058), .B1(KEYINPUT125), .B2(new_n1050), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1054), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT126), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT126), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1054), .A2(new_n1059), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g639(.A(new_n1064), .B(KEYINPUT47), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1048), .A2(new_n1058), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1049), .B1(new_n1048), .B2(new_n939), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n854), .A2(G1996), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1066), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  XOR2_X1   g644(.A(new_n770), .B(new_n773), .Z(new_n1070));
  AOI21_X1  g645(.A(new_n1069), .B1(new_n1048), .B2(new_n1070), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1047), .A2(G1986), .A3(G290), .ZN(new_n1072));
  XOR2_X1   g647(.A(new_n1072), .B(KEYINPUT48), .Z(new_n1073));
  NAND2_X1  g648(.A1(new_n771), .A2(new_n773), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1057), .B1(new_n1069), .B2(new_n1074), .ZN(new_n1075));
  AOI22_X1  g650(.A1(new_n1071), .A2(new_n1073), .B1(new_n1075), .B2(new_n1048), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n1065), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G8), .ZN(new_n1078));
  INV_X1    g653(.A(G1384), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n465), .A2(new_n500), .ZN(new_n1080));
  AOI22_X1  g655(.A1(new_n644), .A2(new_n1080), .B1(KEYINPUT4), .B2(new_n502), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n480), .A2(G102), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n487), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1082), .B1(new_n1083), .B2(new_n461), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1079), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT45), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n509), .A2(KEYINPUT45), .A3(new_n1079), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1087), .A2(new_n1088), .A3(new_n1046), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n805), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1085), .A2(KEYINPUT50), .ZN(new_n1091));
  INV_X1    g666(.A(G2084), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT50), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n509), .A2(new_n1093), .A3(new_n1079), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1091), .A2(new_n1092), .A3(new_n1094), .A4(new_n1046), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1078), .B1(new_n1090), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(G168), .ZN(new_n1097));
  XNOR2_X1  g672(.A(new_n1097), .B(KEYINPUT117), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1091), .A2(new_n1046), .A3(new_n1094), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT115), .B(G2090), .Z(new_n1101));
  OR2_X1    g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n478), .A2(G137), .B1(G101), .B2(new_n480), .ZN(new_n1103));
  INV_X1    g678(.A(new_n474), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1104), .B1(new_n644), .B2(G125), .ZN(new_n1105));
  OAI211_X1 g680(.A(G40), .B(new_n1103), .C1(new_n1105), .C2(new_n465), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1106), .B1(new_n1086), .B2(new_n1085), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n509), .A2(KEYINPUT45), .A3(new_n1043), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(new_n752), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1078), .B1(new_n1102), .B2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(G166), .A2(new_n1078), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1112), .B(KEYINPUT55), .ZN(new_n1113));
  OR2_X1    g688(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  XOR2_X1   g689(.A(KEYINPUT116), .B(G1981), .Z(new_n1115));
  NAND2_X1  g690(.A1(new_n598), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(G1981), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1116), .B1(new_n1117), .B2(new_n598), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT49), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1106), .A2(new_n1085), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1121), .A2(new_n1078), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1116), .B(KEYINPUT49), .C1(new_n1117), .C2(new_n598), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1120), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(G1976), .ZN(new_n1125));
  AOI21_X1  g700(.A(KEYINPUT52), .B1(G288), .B2(new_n1125), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1122), .B(new_n1126), .C1(new_n1125), .C2(G288), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1122), .B1(new_n1125), .B2(G288), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT52), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1124), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1114), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT63), .B1(new_n1099), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1132), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT63), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1134), .A2(new_n1135), .A3(new_n1098), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1124), .A2(new_n1125), .A3(new_n745), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(new_n1116), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1131), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1138), .A2(new_n1122), .B1(new_n1139), .B2(new_n1130), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1133), .A2(new_n1136), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(G1966), .B1(new_n1107), .B2(new_n1088), .ZN(new_n1142));
  AND4_X1   g717(.A1(new_n1092), .A2(new_n1091), .A3(new_n1046), .A4(new_n1094), .ZN(new_n1143));
  OAI21_X1  g718(.A(G8), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(G286), .A2(G8), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1145), .B(KEYINPUT121), .ZN(new_n1146));
  AOI21_X1  g721(.A(KEYINPUT51), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1146), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1148), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1149), .B1(new_n1096), .B2(new_n1148), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1147), .B1(KEYINPUT51), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT62), .ZN(new_n1152));
  OAI21_X1  g727(.A(KEYINPUT124), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(G2078), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1087), .A2(new_n1154), .A3(new_n1108), .A4(new_n1046), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT53), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT122), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(G1961), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1100), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1155), .A2(KEYINPUT122), .A3(new_n1156), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1107), .A2(KEYINPUT53), .A3(new_n1154), .A4(new_n1088), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1159), .A2(new_n1161), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(G171), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1165), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1150), .A2(KEYINPUT51), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1147), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT124), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1169), .A2(new_n1170), .A3(KEYINPUT62), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1153), .A2(new_n1166), .A3(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT61), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT118), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1174), .A2(KEYINPUT57), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT57), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1176), .A2(KEYINPUT118), .ZN(new_n1177));
  OR3_X1    g752(.A1(G299), .A2(new_n1175), .A3(new_n1177), .ZN(new_n1178));
  NAND3_X1  g753(.A1(G299), .A2(new_n1174), .A3(KEYINPUT57), .ZN(new_n1179));
  AND2_X1   g754(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g755(.A(KEYINPUT56), .B(G2072), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1087), .A2(new_n1046), .A3(new_n1108), .A4(new_n1181), .ZN(new_n1182));
  AOI22_X1  g757(.A1(KEYINPUT119), .A2(new_n1182), .B1(new_n1100), .B2(new_n831), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT119), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1107), .A2(new_n1184), .A3(new_n1108), .A4(new_n1181), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1180), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1182), .A2(KEYINPUT119), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1100), .A2(new_n831), .ZN(new_n1188));
  AND4_X1   g763(.A1(new_n1180), .A2(new_n1187), .A3(new_n1185), .A4(new_n1188), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1173), .B1(new_n1186), .B2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1187), .A2(new_n1185), .A3(new_n1188), .ZN(new_n1191));
  INV_X1    g766(.A(new_n1180), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1183), .A2(new_n1180), .A3(new_n1185), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1193), .A2(new_n1194), .A3(KEYINPUT61), .ZN(new_n1195));
  INV_X1    g770(.A(G1348), .ZN(new_n1196));
  AOI22_X1  g771(.A1(new_n1100), .A2(new_n1196), .B1(new_n1056), .B2(new_n1121), .ZN(new_n1197));
  OR2_X1    g772(.A1(new_n1197), .A2(KEYINPUT60), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1100), .A2(new_n1196), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1121), .A2(new_n1056), .ZN(new_n1200));
  AND4_X1   g775(.A1(KEYINPUT60), .A2(new_n1199), .A3(new_n623), .A4(new_n1200), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n623), .B1(new_n1197), .B2(KEYINPUT60), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1198), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g778(.A(KEYINPUT120), .B(G1996), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1107), .A2(new_n1108), .A3(new_n1204), .ZN(new_n1205));
  XOR2_X1   g780(.A(KEYINPUT58), .B(G1341), .Z(new_n1206));
  OAI21_X1  g781(.A(new_n1206), .B1(new_n1106), .B2(new_n1085), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1205), .A2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g783(.A(KEYINPUT59), .B1(new_n1208), .B2(new_n560), .ZN(new_n1209));
  INV_X1    g784(.A(KEYINPUT59), .ZN(new_n1210));
  AOI211_X1 g785(.A(new_n1210), .B(new_n559), .C1(new_n1205), .C2(new_n1207), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n1209), .A2(new_n1211), .ZN(new_n1212));
  NAND4_X1  g787(.A1(new_n1190), .A2(new_n1195), .A3(new_n1203), .A4(new_n1212), .ZN(new_n1213));
  NOR2_X1   g788(.A1(new_n1197), .A2(new_n623), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1186), .B1(new_n1194), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1213), .A2(new_n1215), .ZN(new_n1216));
  AND2_X1   g791(.A1(new_n1162), .A2(new_n1161), .ZN(new_n1217));
  NOR3_X1   g792(.A1(new_n1044), .A2(new_n1156), .A3(G2078), .ZN(new_n1218));
  NAND3_X1  g793(.A1(new_n1218), .A2(new_n1046), .A3(new_n1108), .ZN(new_n1219));
  NAND4_X1  g794(.A1(new_n1217), .A2(G301), .A3(new_n1159), .A4(new_n1219), .ZN(new_n1220));
  AOI21_X1  g795(.A(KEYINPUT54), .B1(new_n1165), .B2(new_n1220), .ZN(new_n1221));
  NOR2_X1   g796(.A1(new_n1221), .A2(new_n1151), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1216), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g798(.A(KEYINPUT54), .ZN(new_n1224));
  NAND4_X1  g799(.A1(new_n1159), .A2(new_n1161), .A3(new_n1162), .A4(new_n1219), .ZN(new_n1225));
  AOI21_X1  g800(.A(new_n1224), .B1(new_n1225), .B2(G171), .ZN(new_n1226));
  INV_X1    g801(.A(KEYINPUT123), .ZN(new_n1227));
  NAND4_X1  g802(.A1(new_n1217), .A2(G301), .A3(new_n1159), .A4(new_n1163), .ZN(new_n1228));
  AND3_X1   g803(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  AOI21_X1  g804(.A(new_n1227), .B1(new_n1226), .B2(new_n1228), .ZN(new_n1230));
  NOR2_X1   g805(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  OAI21_X1  g806(.A(new_n1172), .B1(new_n1223), .B2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g807(.A(new_n1141), .B1(new_n1232), .B2(new_n1134), .ZN(new_n1233));
  XNOR2_X1  g808(.A(G290), .B(new_n731), .ZN(new_n1234));
  OAI21_X1  g809(.A(new_n1071), .B1(new_n1047), .B2(new_n1234), .ZN(new_n1235));
  OAI21_X1  g810(.A(new_n1077), .B1(new_n1233), .B2(new_n1235), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g811(.A1(new_n459), .A2(G227), .ZN(new_n1238));
  AOI21_X1  g812(.A(new_n1238), .B1(new_n687), .B2(new_n690), .ZN(new_n1239));
  NAND3_X1  g813(.A1(new_n736), .A2(new_n1239), .A3(new_n739), .ZN(new_n1240));
  NOR2_X1   g814(.A1(new_n965), .A2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g815(.A(new_n1241), .B1(new_n1036), .B2(new_n1040), .ZN(G225));
  INV_X1    g816(.A(KEYINPUT127), .ZN(new_n1243));
  NAND2_X1  g817(.A1(G225), .A2(new_n1243), .ZN(new_n1244));
  OAI211_X1 g818(.A(new_n1241), .B(KEYINPUT127), .C1(new_n1036), .C2(new_n1040), .ZN(new_n1245));
  NAND2_X1  g819(.A1(new_n1244), .A2(new_n1245), .ZN(G308));
endmodule


