

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595;

  XNOR2_X1 U324 ( .A(n457), .B(KEYINPUT41), .ZN(n458) );
  NOR2_X1 U325 ( .A1(n495), .A2(n483), .ZN(n575) );
  XNOR2_X1 U326 ( .A(n350), .B(n349), .ZN(n551) );
  XOR2_X1 U327 ( .A(G36GAT), .B(G50GAT), .Z(n292) );
  XOR2_X1 U328 ( .A(n426), .B(n425), .Z(n293) );
  XOR2_X1 U329 ( .A(n439), .B(n438), .Z(n294) );
  XNOR2_X1 U330 ( .A(KEYINPUT46), .B(KEYINPUT107), .ZN(n459) );
  XNOR2_X1 U331 ( .A(n460), .B(n459), .ZN(n461) );
  INV_X1 U332 ( .A(KEYINPUT109), .ZN(n465) );
  XNOR2_X1 U333 ( .A(n465), .B(KEYINPUT47), .ZN(n466) );
  INV_X1 U334 ( .A(n551), .ZN(n367) );
  INV_X1 U335 ( .A(KEYINPUT24), .ZN(n341) );
  NAND2_X1 U336 ( .A1(n367), .A2(n366), .ZN(n388) );
  INV_X1 U337 ( .A(KEYINPUT97), .ZN(n399) );
  XNOR2_X1 U338 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U339 ( .A(n441), .B(n292), .ZN(n442) );
  XNOR2_X1 U340 ( .A(n344), .B(n343), .ZN(n348) );
  XNOR2_X1 U341 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U342 ( .A(n443), .B(n442), .ZN(n451) );
  XNOR2_X1 U343 ( .A(n435), .B(n434), .ZN(n437) );
  XNOR2_X1 U344 ( .A(n586), .B(n458), .ZN(n486) );
  INV_X1 U345 ( .A(KEYINPUT28), .ZN(n349) );
  XOR2_X1 U346 ( .A(KEYINPUT124), .B(n582), .Z(n592) );
  XNOR2_X1 U347 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n484) );
  XNOR2_X1 U348 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n455) );
  XNOR2_X1 U349 ( .A(n485), .B(n484), .ZN(G1351GAT) );
  XNOR2_X1 U350 ( .A(n456), .B(n455), .ZN(G1330GAT) );
  XOR2_X1 U351 ( .A(G99GAT), .B(G190GAT), .Z(n296) );
  XOR2_X1 U352 ( .A(KEYINPUT0), .B(G127GAT), .Z(n376) );
  XOR2_X1 U353 ( .A(G120GAT), .B(G71GAT), .Z(n425) );
  XNOR2_X1 U354 ( .A(n376), .B(n425), .ZN(n295) );
  XNOR2_X1 U355 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U356 ( .A(n297), .B(G134GAT), .Z(n302) );
  XOR2_X1 U357 ( .A(KEYINPUT20), .B(KEYINPUT82), .Z(n299) );
  XNOR2_X1 U358 ( .A(G113GAT), .B(KEYINPUT81), .ZN(n298) );
  XNOR2_X1 U359 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U360 ( .A(G43GAT), .B(n300), .ZN(n301) );
  XNOR2_X1 U361 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U362 ( .A(G176GAT), .B(KEYINPUT84), .Z(n304) );
  NAND2_X1 U363 ( .A1(G227GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U364 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U365 ( .A(n306), .B(n305), .Z(n312) );
  XNOR2_X1 U366 ( .A(KEYINPUT83), .B(KEYINPUT18), .ZN(n307) );
  XNOR2_X1 U367 ( .A(n307), .B(KEYINPUT17), .ZN(n308) );
  XOR2_X1 U368 ( .A(n308), .B(KEYINPUT19), .Z(n310) );
  XNOR2_X1 U369 ( .A(G169GAT), .B(G183GAT), .ZN(n309) );
  XNOR2_X1 U370 ( .A(n310), .B(n309), .ZN(n361) );
  XNOR2_X1 U371 ( .A(G15GAT), .B(n361), .ZN(n311) );
  XOR2_X2 U372 ( .A(n312), .B(n311), .Z(n549) );
  XOR2_X1 U373 ( .A(G155GAT), .B(G211GAT), .Z(n314) );
  XNOR2_X1 U374 ( .A(G22GAT), .B(G78GAT), .ZN(n313) );
  XNOR2_X1 U375 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U376 ( .A(G71GAT), .B(G127GAT), .Z(n316) );
  XNOR2_X1 U377 ( .A(G15GAT), .B(G183GAT), .ZN(n315) );
  XNOR2_X1 U378 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U379 ( .A(n318), .B(n317), .Z(n323) );
  XOR2_X1 U380 ( .A(G57GAT), .B(KEYINPUT13), .Z(n431) );
  XOR2_X1 U381 ( .A(G8GAT), .B(KEYINPUT76), .Z(n351) );
  XOR2_X1 U382 ( .A(n351), .B(G64GAT), .Z(n320) );
  NAND2_X1 U383 ( .A1(G231GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U384 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U385 ( .A(n431), .B(n321), .ZN(n322) );
  XNOR2_X1 U386 ( .A(n323), .B(n322), .ZN(n331) );
  XOR2_X1 U387 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n325) );
  XNOR2_X1 U388 ( .A(KEYINPUT78), .B(KEYINPUT77), .ZN(n324) );
  XNOR2_X1 U389 ( .A(n325), .B(n324), .ZN(n329) );
  XOR2_X1 U390 ( .A(KEYINPUT80), .B(KEYINPUT14), .Z(n327) );
  XNOR2_X1 U391 ( .A(G1GAT), .B(KEYINPUT79), .ZN(n326) );
  XNOR2_X1 U392 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U393 ( .A(n329), .B(n328), .Z(n330) );
  XOR2_X1 U394 ( .A(n331), .B(n330), .Z(n510) );
  INV_X1 U395 ( .A(n510), .ZN(n589) );
  XOR2_X1 U396 ( .A(KEYINPUT21), .B(G218GAT), .Z(n333) );
  XNOR2_X1 U397 ( .A(KEYINPUT85), .B(G211GAT), .ZN(n332) );
  XNOR2_X1 U398 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U399 ( .A(G197GAT), .B(n334), .ZN(n362) );
  XOR2_X1 U400 ( .A(G141GAT), .B(G22GAT), .Z(n438) );
  XOR2_X1 U401 ( .A(G50GAT), .B(G162GAT), .Z(n419) );
  XNOR2_X1 U402 ( .A(n438), .B(n419), .ZN(n336) );
  XOR2_X1 U403 ( .A(KEYINPUT86), .B(KEYINPUT22), .Z(n335) );
  XNOR2_X1 U404 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U405 ( .A(n362), .B(n337), .ZN(n339) );
  NAND2_X1 U406 ( .A1(G228GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U407 ( .A(n339), .B(n338), .ZN(n344) );
  XNOR2_X1 U408 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n340) );
  XNOR2_X1 U409 ( .A(n340), .B(KEYINPUT2), .ZN(n383) );
  XNOR2_X1 U410 ( .A(n383), .B(KEYINPUT23), .ZN(n342) );
  XOR2_X1 U411 ( .A(G148GAT), .B(G106GAT), .Z(n346) );
  XNOR2_X1 U412 ( .A(G204GAT), .B(G78GAT), .ZN(n345) );
  XNOR2_X1 U413 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U414 ( .A(KEYINPUT70), .B(n347), .ZN(n436) );
  XNOR2_X1 U415 ( .A(n348), .B(n436), .ZN(n480) );
  XOR2_X1 U416 ( .A(n480), .B(KEYINPUT67), .Z(n350) );
  XOR2_X1 U417 ( .A(G176GAT), .B(G64GAT), .Z(n430) );
  XOR2_X1 U418 ( .A(n430), .B(n351), .Z(n353) );
  XNOR2_X1 U419 ( .A(G204GAT), .B(G92GAT), .ZN(n352) );
  XNOR2_X1 U420 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U421 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n355) );
  NAND2_X1 U422 ( .A1(G226GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U423 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U424 ( .A(n357), .B(n356), .Z(n359) );
  XOR2_X1 U425 ( .A(G36GAT), .B(G190GAT), .Z(n411) );
  XNOR2_X1 U426 ( .A(n411), .B(KEYINPUT90), .ZN(n358) );
  XNOR2_X1 U427 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U428 ( .A(n361), .B(n360), .ZN(n364) );
  INV_X1 U429 ( .A(n362), .ZN(n363) );
  XOR2_X1 U430 ( .A(n364), .B(n363), .Z(n476) );
  INV_X1 U431 ( .A(n476), .ZN(n547) );
  XOR2_X1 U432 ( .A(KEYINPUT27), .B(KEYINPUT93), .Z(n365) );
  XOR2_X1 U433 ( .A(n547), .B(n365), .Z(n492) );
  NOR2_X1 U434 ( .A1(n492), .A2(n549), .ZN(n366) );
  XOR2_X1 U435 ( .A(KEYINPUT89), .B(KEYINPUT6), .Z(n369) );
  XNOR2_X1 U436 ( .A(KEYINPUT87), .B(KEYINPUT1), .ZN(n368) );
  XNOR2_X1 U437 ( .A(n369), .B(n368), .ZN(n387) );
  XOR2_X1 U438 ( .A(G85GAT), .B(G162GAT), .Z(n371) );
  XNOR2_X1 U439 ( .A(G29GAT), .B(G148GAT), .ZN(n370) );
  XNOR2_X1 U440 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U441 ( .A(KEYINPUT88), .B(G57GAT), .Z(n373) );
  XNOR2_X1 U442 ( .A(G141GAT), .B(G120GAT), .ZN(n372) );
  XNOR2_X1 U443 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U444 ( .A(n375), .B(n374), .Z(n381) );
  XOR2_X1 U445 ( .A(G113GAT), .B(G1GAT), .Z(n441) );
  XOR2_X1 U446 ( .A(G134GAT), .B(KEYINPUT75), .Z(n410) );
  XOR2_X1 U447 ( .A(n410), .B(n376), .Z(n378) );
  NAND2_X1 U448 ( .A1(G225GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U449 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U450 ( .A(n441), .B(n379), .ZN(n380) );
  XNOR2_X1 U451 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U452 ( .A(n382), .B(KEYINPUT5), .Z(n385) );
  XNOR2_X1 U453 ( .A(n383), .B(KEYINPUT4), .ZN(n384) );
  XNOR2_X1 U454 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U455 ( .A(n387), .B(n386), .ZN(n544) );
  NAND2_X1 U456 ( .A1(n388), .A2(n544), .ZN(n398) );
  NAND2_X1 U457 ( .A1(n547), .A2(n549), .ZN(n389) );
  NAND2_X1 U458 ( .A1(n480), .A2(n389), .ZN(n390) );
  XOR2_X1 U459 ( .A(KEYINPUT25), .B(n390), .Z(n396) );
  NOR2_X1 U460 ( .A1(n480), .A2(n549), .ZN(n392) );
  XNOR2_X1 U461 ( .A(KEYINPUT95), .B(KEYINPUT26), .ZN(n391) );
  XNOR2_X1 U462 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U463 ( .A(KEYINPUT94), .B(n393), .ZN(n560) );
  NOR2_X1 U464 ( .A1(n492), .A2(n560), .ZN(n394) );
  NOR2_X1 U465 ( .A1(n544), .A2(n394), .ZN(n395) );
  NAND2_X1 U466 ( .A1(n396), .A2(n395), .ZN(n397) );
  NAND2_X1 U467 ( .A1(n398), .A2(n397), .ZN(n512) );
  NOR2_X1 U468 ( .A1(n589), .A2(n512), .ZN(n400) );
  XNOR2_X1 U469 ( .A(n400), .B(n399), .ZN(n422) );
  XOR2_X1 U470 ( .A(KEYINPUT73), .B(KEYINPUT11), .Z(n402) );
  NAND2_X1 U471 ( .A1(G232GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U472 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U473 ( .A(n403), .B(KEYINPUT9), .Z(n409) );
  XOR2_X1 U474 ( .A(G29GAT), .B(G43GAT), .Z(n405) );
  XNOR2_X1 U475 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n404) );
  XNOR2_X1 U476 ( .A(n405), .B(n404), .ZN(n439) );
  XOR2_X1 U477 ( .A(G92GAT), .B(KEYINPUT71), .Z(n407) );
  XNOR2_X1 U478 ( .A(G99GAT), .B(G85GAT), .ZN(n406) );
  XNOR2_X1 U479 ( .A(n407), .B(n406), .ZN(n426) );
  XNOR2_X1 U480 ( .A(n439), .B(n426), .ZN(n408) );
  XNOR2_X1 U481 ( .A(n409), .B(n408), .ZN(n415) );
  XOR2_X1 U482 ( .A(n411), .B(n410), .Z(n413) );
  XNOR2_X1 U483 ( .A(G106GAT), .B(G218GAT), .ZN(n412) );
  XNOR2_X1 U484 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U485 ( .A(n415), .B(n414), .Z(n421) );
  XOR2_X1 U486 ( .A(KEYINPUT10), .B(KEYINPUT66), .Z(n417) );
  XNOR2_X1 U487 ( .A(KEYINPUT74), .B(KEYINPUT65), .ZN(n416) );
  XNOR2_X1 U488 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U489 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U490 ( .A(n421), .B(n420), .ZN(n571) );
  XNOR2_X1 U491 ( .A(n571), .B(KEYINPUT36), .ZN(n591) );
  NAND2_X1 U492 ( .A1(n422), .A2(n591), .ZN(n424) );
  XOR2_X1 U493 ( .A(KEYINPUT98), .B(KEYINPUT37), .Z(n423) );
  XNOR2_X1 U494 ( .A(n424), .B(n423), .ZN(n543) );
  NAND2_X1 U495 ( .A1(G230GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U496 ( .A(n293), .B(n427), .ZN(n435) );
  XOR2_X1 U497 ( .A(KEYINPUT72), .B(KEYINPUT31), .Z(n429) );
  XNOR2_X1 U498 ( .A(KEYINPUT33), .B(KEYINPUT32), .ZN(n428) );
  XOR2_X1 U499 ( .A(n429), .B(n428), .Z(n433) );
  XNOR2_X1 U500 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U501 ( .A(n437), .B(n436), .Z(n586) );
  NAND2_X1 U502 ( .A1(G229GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U503 ( .A(n294), .B(n440), .ZN(n443) );
  XOR2_X1 U504 ( .A(G8GAT), .B(G15GAT), .Z(n445) );
  XNOR2_X1 U505 ( .A(G169GAT), .B(G197GAT), .ZN(n444) );
  XNOR2_X1 U506 ( .A(n445), .B(n444), .ZN(n449) );
  XOR2_X1 U507 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n447) );
  XNOR2_X1 U508 ( .A(KEYINPUT29), .B(KEYINPUT69), .ZN(n446) );
  XNOR2_X1 U509 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U510 ( .A(n449), .B(n448), .Z(n450) );
  XOR2_X1 U511 ( .A(n451), .B(n450), .Z(n531) );
  OR2_X1 U512 ( .A1(n586), .A2(n531), .ZN(n515) );
  NOR2_X1 U513 ( .A1(n543), .A2(n515), .ZN(n453) );
  XNOR2_X1 U514 ( .A(KEYINPUT100), .B(KEYINPUT38), .ZN(n452) );
  XNOR2_X1 U515 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X1 U516 ( .A(KEYINPUT99), .B(n454), .Z(n528) );
  NAND2_X1 U517 ( .A1(n549), .A2(n528), .ZN(n456) );
  INV_X1 U518 ( .A(n549), .ZN(n495) );
  XOR2_X1 U519 ( .A(KEYINPUT122), .B(KEYINPUT55), .Z(n482) );
  INV_X1 U520 ( .A(KEYINPUT48), .ZN(n475) );
  INV_X1 U521 ( .A(KEYINPUT108), .ZN(n463) );
  INV_X1 U522 ( .A(n531), .ZN(n583) );
  INV_X1 U523 ( .A(KEYINPUT64), .ZN(n457) );
  NAND2_X1 U524 ( .A1(n583), .A2(n486), .ZN(n460) );
  NOR2_X1 U525 ( .A1(n461), .A2(n589), .ZN(n462) );
  XNOR2_X1 U526 ( .A(n463), .B(n462), .ZN(n464) );
  NOR2_X1 U527 ( .A1(n571), .A2(n464), .ZN(n467) );
  XNOR2_X1 U528 ( .A(n467), .B(n466), .ZN(n473) );
  XOR2_X1 U529 ( .A(KEYINPUT45), .B(KEYINPUT110), .Z(n469) );
  NAND2_X1 U530 ( .A1(n591), .A2(n589), .ZN(n468) );
  XNOR2_X1 U531 ( .A(n469), .B(n468), .ZN(n471) );
  NOR2_X1 U532 ( .A1(n583), .A2(n586), .ZN(n470) );
  NAND2_X1 U533 ( .A1(n471), .A2(n470), .ZN(n472) );
  NAND2_X1 U534 ( .A1(n473), .A2(n472), .ZN(n474) );
  XNOR2_X1 U535 ( .A(n475), .B(n474), .ZN(n491) );
  NOR2_X1 U536 ( .A1(n491), .A2(n476), .ZN(n478) );
  INV_X1 U537 ( .A(KEYINPUT54), .ZN(n477) );
  XNOR2_X1 U538 ( .A(n478), .B(n477), .ZN(n479) );
  NOR2_X1 U539 ( .A1(n479), .A2(n544), .ZN(n581) );
  NAND2_X1 U540 ( .A1(n581), .A2(n480), .ZN(n481) );
  XNOR2_X1 U541 ( .A(n482), .B(n481), .ZN(n483) );
  NAND2_X1 U542 ( .A1(n575), .A2(n571), .ZN(n485) );
  NAND2_X1 U543 ( .A1(n575), .A2(n486), .ZN(n490) );
  XOR2_X1 U544 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n488) );
  XOR2_X1 U545 ( .A(G176GAT), .B(KEYINPUT123), .Z(n487) );
  XNOR2_X1 U546 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U547 ( .A(n490), .B(n489), .ZN(G1349GAT) );
  XOR2_X1 U548 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n499) );
  NOR2_X1 U549 ( .A1(n492), .A2(n491), .ZN(n493) );
  NAND2_X1 U550 ( .A1(n493), .A2(n544), .ZN(n494) );
  XNOR2_X1 U551 ( .A(KEYINPUT111), .B(n494), .ZN(n561) );
  NOR2_X1 U552 ( .A1(n551), .A2(n495), .ZN(n496) );
  AND2_X1 U553 ( .A1(n561), .A2(n496), .ZN(n497) );
  XNOR2_X1 U554 ( .A(n497), .B(KEYINPUT112), .ZN(n556) );
  NAND2_X1 U555 ( .A1(n556), .A2(n589), .ZN(n498) );
  XNOR2_X1 U556 ( .A(n499), .B(n498), .ZN(n501) );
  INV_X1 U557 ( .A(G127GAT), .ZN(n500) );
  XNOR2_X1 U558 ( .A(n501), .B(n500), .ZN(G1342GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n503) );
  NAND2_X1 U560 ( .A1(n486), .A2(n556), .ZN(n502) );
  XNOR2_X1 U561 ( .A(n503), .B(n502), .ZN(n505) );
  INV_X1 U562 ( .A(G120GAT), .ZN(n504) );
  XNOR2_X1 U563 ( .A(n505), .B(n504), .ZN(G1341GAT) );
  INV_X1 U564 ( .A(G134GAT), .ZN(n509) );
  XOR2_X1 U565 ( .A(KEYINPUT51), .B(KEYINPUT117), .Z(n507) );
  NAND2_X1 U566 ( .A1(n571), .A2(n556), .ZN(n506) );
  XNOR2_X1 U567 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U568 ( .A(n509), .B(n508), .ZN(G1343GAT) );
  XNOR2_X1 U569 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n517) );
  NOR2_X1 U570 ( .A1(n571), .A2(n510), .ZN(n511) );
  XNOR2_X1 U571 ( .A(KEYINPUT16), .B(n511), .ZN(n514) );
  INV_X1 U572 ( .A(n512), .ZN(n513) );
  NAND2_X1 U573 ( .A1(n514), .A2(n513), .ZN(n532) );
  NOR2_X1 U574 ( .A1(n515), .A2(n532), .ZN(n522) );
  NAND2_X1 U575 ( .A1(n522), .A2(n544), .ZN(n516) );
  XNOR2_X1 U576 ( .A(n517), .B(n516), .ZN(G1324GAT) );
  NAND2_X1 U577 ( .A1(n522), .A2(n547), .ZN(n518) );
  XNOR2_X1 U578 ( .A(n518), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT96), .B(KEYINPUT35), .Z(n520) );
  NAND2_X1 U580 ( .A1(n522), .A2(n549), .ZN(n519) );
  XNOR2_X1 U581 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U582 ( .A(G15GAT), .B(n521), .ZN(G1326GAT) );
  NAND2_X1 U583 ( .A1(n522), .A2(n551), .ZN(n523) );
  XNOR2_X1 U584 ( .A(n523), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U585 ( .A1(n544), .A2(n528), .ZN(n526) );
  XNOR2_X1 U586 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n524) );
  XNOR2_X1 U587 ( .A(n524), .B(KEYINPUT101), .ZN(n525) );
  XNOR2_X1 U588 ( .A(n526), .B(n525), .ZN(G1328GAT) );
  NAND2_X1 U589 ( .A1(n528), .A2(n547), .ZN(n527) );
  XNOR2_X1 U590 ( .A(n527), .B(G36GAT), .ZN(G1329GAT) );
  XNOR2_X1 U591 ( .A(G50GAT), .B(KEYINPUT102), .ZN(n530) );
  NAND2_X1 U592 ( .A1(n551), .A2(n528), .ZN(n529) );
  XNOR2_X1 U593 ( .A(n530), .B(n529), .ZN(G1331GAT) );
  NAND2_X1 U594 ( .A1(n531), .A2(n486), .ZN(n542) );
  NOR2_X1 U595 ( .A1(n532), .A2(n542), .ZN(n533) );
  XNOR2_X1 U596 ( .A(n533), .B(KEYINPUT104), .ZN(n539) );
  NAND2_X1 U597 ( .A1(n539), .A2(n544), .ZN(n536) );
  XOR2_X1 U598 ( .A(G57GAT), .B(KEYINPUT103), .Z(n534) );
  XNOR2_X1 U599 ( .A(KEYINPUT42), .B(n534), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n536), .B(n535), .ZN(G1332GAT) );
  NAND2_X1 U601 ( .A1(n539), .A2(n547), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n537), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U603 ( .A1(n539), .A2(n549), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n538), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U605 ( .A(G78GAT), .B(KEYINPUT43), .Z(n541) );
  NAND2_X1 U606 ( .A1(n551), .A2(n539), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(G1335GAT) );
  XOR2_X1 U608 ( .A(G85GAT), .B(KEYINPUT105), .Z(n546) );
  NOR2_X1 U609 ( .A1(n543), .A2(n542), .ZN(n552) );
  NAND2_X1 U610 ( .A1(n552), .A2(n544), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n546), .B(n545), .ZN(G1336GAT) );
  NAND2_X1 U612 ( .A1(n552), .A2(n547), .ZN(n548) );
  XNOR2_X1 U613 ( .A(n548), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U614 ( .A1(n549), .A2(n552), .ZN(n550) );
  XNOR2_X1 U615 ( .A(n550), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT44), .B(KEYINPUT106), .Z(n554) );
  NAND2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U619 ( .A(G106GAT), .B(n555), .Z(G1339GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n558) );
  NAND2_X1 U621 ( .A1(n556), .A2(n583), .ZN(n557) );
  XNOR2_X1 U622 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U623 ( .A(G113GAT), .B(n559), .ZN(G1340GAT) );
  INV_X1 U624 ( .A(n560), .ZN(n580) );
  AND2_X1 U625 ( .A1(n580), .A2(n561), .ZN(n572) );
  NAND2_X1 U626 ( .A1(n572), .A2(n583), .ZN(n562) );
  XNOR2_X1 U627 ( .A(KEYINPUT118), .B(n562), .ZN(n563) );
  XNOR2_X1 U628 ( .A(G141GAT), .B(n563), .ZN(G1344GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT119), .B(KEYINPUT53), .Z(n565) );
  NAND2_X1 U630 ( .A1(n572), .A2(n486), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(n567) );
  XOR2_X1 U632 ( .A(G148GAT), .B(KEYINPUT52), .Z(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(G1345GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n569) );
  NAND2_X1 U635 ( .A1(n572), .A2(n589), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U637 ( .A(G155GAT), .B(n570), .ZN(G1346GAT) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n573), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U640 ( .A1(n583), .A2(n575), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n574), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U642 ( .A1(n589), .A2(n575), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n576), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n578) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n577) );
  XNOR2_X1 U646 ( .A(n578), .B(n577), .ZN(n579) );
  XOR2_X1 U647 ( .A(KEYINPUT59), .B(n579), .Z(n585) );
  NAND2_X1 U648 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U649 ( .A1(n592), .A2(n583), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1352GAT) );
  XOR2_X1 U651 ( .A(G204GAT), .B(KEYINPUT61), .Z(n588) );
  NAND2_X1 U652 ( .A1(n592), .A2(n586), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(G1353GAT) );
  NAND2_X1 U654 ( .A1(n592), .A2(n589), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n590), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U656 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n594) );
  NAND2_X1 U657 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U658 ( .A(n594), .B(n593), .ZN(n595) );
  XNOR2_X1 U659 ( .A(n595), .B(G218GAT), .ZN(G1355GAT) );
endmodule

