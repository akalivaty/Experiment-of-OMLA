//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 1 1 0 0 0 0 1 1 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 0 0 0 0 1 0 1 1 0 1 1 1 0 1 0 0 0 0 0 1 0 1 1 0 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n539, new_n541, new_n542, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n555, new_n556, new_n558, new_n559, new_n560, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n601, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT64), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  OR2_X1    g027(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT65), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  AOI22_X1  g030(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n452), .ZN(G319));
  INV_X1    g031(.A(G2105), .ZN(new_n457));
  INV_X1    g032(.A(G2104), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(KEYINPUT3), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n459), .A2(new_n461), .A3(G125), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n457), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n459), .A2(new_n461), .A3(G137), .ZN(new_n465));
  NAND2_X1  g040(.A1(G101), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n464), .A2(new_n467), .ZN(G160));
  NAND2_X1  g043(.A1(new_n459), .A2(new_n461), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G136), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n469), .A2(new_n457), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G124), .ZN(new_n473));
  OAI21_X1  g048(.A(G2104), .B1(new_n457), .B2(G112), .ZN(new_n474));
  NOR2_X1   g049(.A1(G100), .A2(G2105), .ZN(new_n475));
  XOR2_X1   g050(.A(new_n475), .B(KEYINPUT66), .Z(new_n476));
  OAI211_X1 g051(.A(new_n471), .B(new_n473), .C1(new_n474), .C2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G162));
  NAND2_X1  g053(.A1(G114), .A2(G2104), .ZN(new_n479));
  INV_X1    g054(.A(G126), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n479), .B1(new_n469), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n458), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G102), .ZN(new_n484));
  NAND4_X1  g059(.A1(new_n459), .A2(new_n461), .A3(G138), .A4(new_n457), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g062(.A(KEYINPUT3), .B(G2104), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n488), .A2(KEYINPUT4), .A3(G138), .A4(new_n457), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n482), .A2(new_n484), .A3(new_n487), .A4(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G164));
  AND2_X1   g066(.A1(KEYINPUT6), .A2(G651), .ZN(new_n492));
  NOR2_X1   g067(.A1(KEYINPUT6), .A2(G651), .ZN(new_n493));
  OAI211_X1 g068(.A(G50), .B(G543), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G543), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT5), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT5), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G543), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n496), .B(new_n498), .C1(new_n492), .C2(new_n493), .ZN(new_n499));
  INV_X1    g074(.A(G88), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n494), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT67), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n496), .A2(new_n498), .ZN(new_n503));
  INV_X1    g078(.A(G62), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(G75), .A2(G543), .ZN(new_n506));
  XOR2_X1   g081(.A(new_n506), .B(KEYINPUT68), .Z(new_n507));
  NAND4_X1  g082(.A1(new_n496), .A2(new_n498), .A3(KEYINPUT67), .A4(G62), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n505), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n501), .B1(new_n509), .B2(G651), .ZN(G166));
  AND2_X1   g085(.A1(new_n496), .A2(new_n498), .ZN(new_n511));
  OR2_X1    g086(.A1(new_n492), .A2(new_n493), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n512), .A2(G89), .ZN(new_n513));
  AND2_X1   g088(.A1(G63), .A2(G651), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n511), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n492), .A2(new_n493), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n516), .A2(new_n495), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G51), .ZN(new_n518));
  XOR2_X1   g093(.A(KEYINPUT69), .B(KEYINPUT7), .Z(new_n519));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n519), .B(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n515), .A2(new_n518), .A3(new_n521), .ZN(G286));
  INV_X1    g097(.A(G286), .ZN(G168));
  AOI22_X1  g098(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n524));
  INV_X1    g099(.A(G651), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n512), .A2(G543), .ZN(new_n527));
  INV_X1    g102(.A(G52), .ZN(new_n528));
  INV_X1    g103(.A(G90), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n527), .A2(new_n528), .B1(new_n529), .B2(new_n499), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n526), .A2(new_n530), .ZN(G171));
  AOI22_X1  g106(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n525), .ZN(new_n533));
  INV_X1    g108(.A(G43), .ZN(new_n534));
  INV_X1    g109(.A(G81), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n527), .A2(new_n534), .B1(new_n535), .B2(new_n499), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G860), .ZN(G153));
  AND3_X1   g113(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G36), .ZN(G176));
  NAND2_X1  g115(.A1(G1), .A2(G3), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT8), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n539), .A2(new_n542), .ZN(G188));
  INV_X1    g118(.A(KEYINPUT9), .ZN(new_n544));
  INV_X1    g119(.A(G53), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n527), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n517), .A2(KEYINPUT9), .A3(G53), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n499), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G91), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n511), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n551), .B2(new_n525), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n548), .A2(new_n552), .ZN(G299));
  INV_X1    g128(.A(G171), .ZN(G301));
  NAND2_X1  g129(.A1(new_n509), .A2(G651), .ZN(new_n555));
  INV_X1    g130(.A(new_n501), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(G303));
  NAND2_X1  g132(.A1(new_n549), .A2(G87), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n517), .A2(G49), .ZN(new_n559));
  OAI21_X1  g134(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(G288));
  INV_X1    g136(.A(G48), .ZN(new_n562));
  INV_X1    g137(.A(G86), .ZN(new_n563));
  OAI22_X1  g138(.A1(new_n527), .A2(new_n562), .B1(new_n563), .B2(new_n499), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n511), .A2(G61), .ZN(new_n565));
  NAND2_X1  g140(.A1(G73), .A2(G543), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n525), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  XOR2_X1   g143(.A(new_n568), .B(KEYINPUT70), .Z(G305));
  NAND2_X1  g144(.A1(G72), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G60), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n503), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G651), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT71), .ZN(new_n574));
  INV_X1    g149(.A(G47), .ZN(new_n575));
  INV_X1    g150(.A(G85), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n527), .A2(new_n575), .B1(new_n576), .B2(new_n499), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n574), .A2(new_n578), .ZN(G290));
  INV_X1    g154(.A(G868), .ZN(new_n580));
  OAI21_X1  g155(.A(KEYINPUT72), .B1(G171), .B2(new_n580), .ZN(new_n581));
  OR3_X1    g156(.A1(G171), .A2(KEYINPUT72), .A3(new_n580), .ZN(new_n582));
  NAND2_X1  g157(.A1(G79), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G66), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n503), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(G651), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n512), .A2(G54), .A3(G543), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(KEYINPUT73), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT73), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n586), .A2(new_n590), .A3(new_n587), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n549), .A2(G92), .ZN(new_n593));
  XOR2_X1   g168(.A(new_n593), .B(KEYINPUT10), .Z(new_n594));
  AND3_X1   g169(.A1(new_n592), .A2(new_n594), .A3(KEYINPUT74), .ZN(new_n595));
  AOI21_X1  g170(.A(KEYINPUT74), .B1(new_n592), .B2(new_n594), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI211_X1 g172(.A(new_n581), .B(new_n582), .C1(new_n597), .C2(G868), .ZN(G284));
  OAI211_X1 g173(.A(new_n581), .B(new_n582), .C1(new_n597), .C2(G868), .ZN(G321));
  NAND2_X1  g174(.A1(G286), .A2(G868), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n548), .A2(new_n552), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(G868), .ZN(G297));
  OAI21_X1  g177(.A(new_n600), .B1(new_n601), .B2(G868), .ZN(G280));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n597), .B1(new_n604), .B2(G860), .ZN(G148));
  INV_X1    g180(.A(new_n537), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(new_n580), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n592), .A2(new_n594), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT74), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n592), .A2(new_n594), .A3(KEYINPUT74), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n612), .A2(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n607), .B1(new_n613), .B2(new_n580), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n488), .A2(new_n483), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT12), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT13), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2100), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n470), .A2(G135), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n472), .A2(G123), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n622), .A2(KEYINPUT76), .ZN(new_n623));
  OAI21_X1  g198(.A(KEYINPUT75), .B1(new_n457), .B2(G111), .ZN(new_n624));
  OR3_X1    g199(.A1(new_n457), .A2(KEYINPUT75), .A3(G111), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n622), .A2(KEYINPUT76), .ZN(new_n626));
  NAND4_X1  g201(.A1(new_n623), .A2(new_n624), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n620), .A2(new_n621), .A3(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(KEYINPUT77), .B(G2096), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n619), .A2(new_n630), .ZN(G156));
  XNOR2_X1  g206(.A(G2443), .B(G2446), .ZN(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2430), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2435), .ZN(new_n635));
  XOR2_X1   g210(.A(G2427), .B(G2438), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(KEYINPUT14), .ZN(new_n638));
  XOR2_X1   g213(.A(G2451), .B(G2454), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n638), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G1341), .B(G1348), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n641), .A2(new_n642), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n633), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n647), .A2(new_n632), .A3(new_n643), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n646), .A2(new_n648), .A3(G14), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(G401));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2067), .B(G2678), .Z(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(new_n655), .A3(KEYINPUT17), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT18), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2072), .B(G2078), .Z(new_n659));
  AOI21_X1  g234(.A(new_n659), .B1(new_n654), .B2(KEYINPUT18), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n658), .B(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2096), .B(G2100), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT78), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n661), .B(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(G227));
  XOR2_X1   g240(.A(G1971), .B(G1976), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  XOR2_X1   g242(.A(G1956), .B(G2474), .Z(new_n668));
  XOR2_X1   g243(.A(G1961), .B(G1966), .Z(new_n669));
  AOI21_X1  g244(.A(KEYINPUT79), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AND3_X1   g245(.A1(new_n668), .A2(new_n669), .A3(KEYINPUT79), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n667), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT20), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n668), .A2(new_n669), .ZN(new_n674));
  AOI22_X1  g249(.A1(new_n672), .A2(new_n673), .B1(new_n667), .B2(new_n674), .ZN(new_n675));
  AND2_X1   g250(.A1(new_n668), .A2(new_n669), .ZN(new_n676));
  OR3_X1    g251(.A1(new_n667), .A2(new_n676), .A3(new_n674), .ZN(new_n677));
  OAI211_X1 g252(.A(new_n675), .B(new_n677), .C1(new_n673), .C2(new_n672), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(G1986), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n678), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n678), .B(new_n679), .ZN(new_n684));
  INV_X1    g259(.A(new_n682), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT22), .B(G1981), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n683), .A2(new_n686), .A3(new_n688), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(G229));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G4), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(new_n597), .B2(new_n694), .ZN(new_n696));
  INV_X1    g271(.A(G1348), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G33), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n457), .A2(G103), .A3(G2104), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT25), .Z(new_n702));
  NAND2_X1  g277(.A1(new_n470), .A2(G139), .ZN(new_n703));
  AOI22_X1  g278(.A1(new_n488), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n702), .B(new_n703), .C1(new_n457), .C2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n700), .B1(new_n706), .B2(new_n699), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT92), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n708), .A2(G2072), .ZN(new_n709));
  NAND2_X1  g284(.A1(G160), .A2(G29), .ZN(new_n710));
  AND2_X1   g285(.A1(KEYINPUT24), .A2(G34), .ZN(new_n711));
  NOR2_X1   g286(.A1(KEYINPUT24), .A2(G34), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n699), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(G2084), .B1(new_n710), .B2(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(G16), .A2(G21), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G168), .B2(G16), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n714), .B1(new_n716), .B2(G1966), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n698), .A2(new_n709), .A3(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n716), .A2(G1966), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n699), .A2(G26), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT28), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n472), .A2(G128), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n470), .A2(G140), .ZN(new_n723));
  OR2_X1    g298(.A1(G104), .A2(G2105), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n724), .B(G2104), .C1(G116), .C2(new_n457), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n722), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT89), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g303(.A1(new_n722), .A2(new_n723), .A3(KEYINPUT89), .A4(new_n725), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AND3_X1   g305(.A1(new_n730), .A2(KEYINPUT90), .A3(G29), .ZN(new_n731));
  AOI21_X1  g306(.A(KEYINPUT90), .B1(new_n730), .B2(G29), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n721), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT91), .B(G2067), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NOR3_X1   g310(.A1(new_n718), .A2(new_n719), .A3(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(G5), .A2(G16), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G171), .B2(G16), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n738), .A2(G1961), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n694), .A2(G19), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n537), .B2(new_n694), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT87), .B(G1341), .Z(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT88), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n741), .B(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G35), .ZN(new_n745));
  OAI21_X1  g320(.A(KEYINPUT94), .B1(new_n745), .B2(G29), .ZN(new_n746));
  OR3_X1    g321(.A1(new_n745), .A2(KEYINPUT94), .A3(G29), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n746), .B(new_n747), .C1(G162), .C2(new_n699), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT29), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n749), .A2(G2090), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n699), .A2(G27), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G164), .B2(new_n699), .ZN(new_n752));
  INV_X1    g327(.A(G2078), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT31), .B(G11), .Z(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT93), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT30), .B(G28), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n756), .B1(new_n699), .B2(new_n757), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n754), .B(new_n758), .C1(new_n749), .C2(G2090), .ZN(new_n759));
  AND2_X1   g334(.A1(new_n708), .A2(G2072), .ZN(new_n760));
  NOR3_X1   g335(.A1(new_n750), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  AOI22_X1  g336(.A1(G129), .A2(new_n472), .B1(new_n470), .B2(G141), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n483), .A2(G105), .ZN(new_n763));
  NAND3_X1  g338(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT26), .Z(new_n765));
  NAND3_X1  g340(.A1(new_n762), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(G29), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G29), .B2(G32), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT27), .B(G1996), .Z(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n694), .A2(KEYINPUT23), .A3(G20), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT23), .ZN(new_n774));
  INV_X1    g349(.A(G20), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(G16), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n773), .B(new_n776), .C1(new_n601), .C2(new_n694), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(G1956), .Z(new_n778));
  NAND2_X1  g353(.A1(new_n738), .A2(G1961), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n710), .A2(G2084), .A3(new_n713), .ZN(new_n780));
  AND4_X1   g355(.A1(new_n772), .A2(new_n778), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n769), .A2(new_n771), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n628), .A2(new_n699), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n761), .A2(new_n781), .A3(new_n782), .A4(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n736), .A2(new_n739), .A3(new_n744), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(KEYINPUT95), .ZN(new_n788));
  NOR4_X1   g363(.A1(new_n785), .A2(new_n718), .A3(new_n719), .A4(new_n735), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT95), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n789), .A2(new_n790), .A3(new_n739), .A4(new_n744), .ZN(new_n791));
  MUX2_X1   g366(.A(G6), .B(G305), .S(G16), .Z(new_n792));
  XOR2_X1   g367(.A(KEYINPUT32), .B(G1981), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT85), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n792), .B(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(G16), .A2(G23), .ZN(new_n796));
  INV_X1    g371(.A(G288), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(G16), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT33), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G1976), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n694), .A2(G22), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G166), .B2(new_n694), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT86), .B(G1971), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n795), .A2(new_n800), .A3(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT34), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n795), .A2(new_n800), .A3(KEYINPUT34), .A4(new_n804), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(G16), .A2(G24), .ZN(new_n810));
  XNOR2_X1  g385(.A(G290), .B(KEYINPUT83), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(G16), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT84), .B(G1986), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n699), .A2(G25), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n470), .A2(G131), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT80), .ZN(new_n817));
  OAI21_X1  g392(.A(G2104), .B1(new_n457), .B2(G107), .ZN(new_n818));
  INV_X1    g393(.A(G95), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n818), .B1(new_n819), .B2(new_n457), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n472), .A2(G119), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(KEYINPUT81), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT81), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n472), .A2(new_n823), .A3(G119), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n820), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT82), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n817), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n826), .B1(new_n817), .B2(new_n825), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n815), .B1(new_n830), .B2(new_n699), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT35), .B(G1991), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n831), .A2(new_n832), .ZN(new_n834));
  NOR3_X1   g409(.A1(new_n814), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n809), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(KEYINPUT36), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT36), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n809), .A2(new_n838), .A3(new_n835), .ZN(new_n839));
  AOI22_X1  g414(.A1(new_n788), .A2(new_n791), .B1(new_n837), .B2(new_n839), .ZN(G311));
  NAND2_X1  g415(.A1(new_n788), .A2(new_n791), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n837), .A2(new_n839), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(G150));
  AOI22_X1  g418(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n844), .A2(new_n525), .ZN(new_n845));
  INV_X1    g420(.A(G55), .ZN(new_n846));
  INV_X1    g421(.A(G93), .ZN(new_n847));
  OAI22_X1  g422(.A1(new_n527), .A2(new_n846), .B1(new_n847), .B2(new_n499), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(G860), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT37), .Z(new_n851));
  NOR2_X1   g426(.A1(new_n612), .A2(new_n604), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT38), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT39), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT96), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n849), .A2(new_n855), .ZN(new_n856));
  OR3_X1    g431(.A1(new_n845), .A2(new_n848), .A3(new_n855), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n856), .A2(new_n537), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n606), .A2(new_n849), .A3(new_n855), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n854), .B(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n851), .B1(new_n861), .B2(G860), .ZN(G145));
  INV_X1    g437(.A(G37), .ZN(new_n863));
  INV_X1    g438(.A(new_n829), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n617), .B(KEYINPUT98), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n866), .A3(new_n827), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n865), .B1(new_n828), .B2(new_n829), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n470), .A2(G142), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n472), .A2(G130), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n870), .A2(KEYINPUT97), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(KEYINPUT97), .ZN(new_n872));
  OR2_X1    g447(.A1(G106), .A2(G2105), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n873), .B(G2104), .C1(G118), .C2(new_n457), .ZN(new_n874));
  AND4_X1   g449(.A1(new_n869), .A2(new_n871), .A3(new_n872), .A4(new_n874), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n867), .A2(new_n868), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n875), .B1(new_n867), .B2(new_n868), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n730), .A2(G164), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n728), .A2(new_n490), .A3(new_n729), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(new_n766), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n766), .B1(new_n879), .B2(new_n880), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n705), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n883), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n885), .A2(new_n706), .A3(new_n881), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n878), .A2(new_n887), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n884), .B(new_n886), .C1(new_n876), .C2(new_n877), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n628), .B(G160), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(G162), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n888), .A2(new_n889), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT99), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n888), .A2(new_n894), .A3(new_n889), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n891), .B1(new_n889), .B2(new_n894), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n863), .B(new_n893), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(KEYINPUT100), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n888), .A2(new_n894), .A3(new_n889), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n899), .B(new_n891), .C1(new_n894), .C2(new_n889), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT100), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n900), .A2(new_n901), .A3(new_n863), .A4(new_n893), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n898), .A2(new_n902), .A3(KEYINPUT40), .ZN(new_n903));
  AOI21_X1  g478(.A(KEYINPUT40), .B1(new_n898), .B2(new_n902), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(G395));
  NAND3_X1  g480(.A1(new_n592), .A2(new_n594), .A3(new_n601), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n601), .B1(new_n592), .B2(new_n594), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT102), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT41), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  OR3_X1    g487(.A1(new_n907), .A2(KEYINPUT41), .A3(new_n908), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT41), .B1(new_n907), .B2(new_n908), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n913), .A2(KEYINPUT102), .A3(new_n914), .ZN(new_n915));
  OR2_X1    g490(.A1(new_n860), .A2(KEYINPUT101), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n860), .A2(KEYINPUT101), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(new_n613), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n613), .B1(new_n916), .B2(new_n917), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n912), .B(new_n915), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n920), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n922), .A2(new_n909), .A3(new_n918), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT42), .ZN(new_n925));
  INV_X1    g500(.A(G290), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n797), .B(G166), .ZN(new_n927));
  OR2_X1    g502(.A1(G305), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(G305), .A2(new_n927), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n928), .A2(new_n926), .A3(new_n929), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT42), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n921), .A2(new_n934), .A3(new_n923), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n925), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n933), .B1(new_n925), .B2(new_n935), .ZN(new_n937));
  OAI21_X1  g512(.A(G868), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n849), .A2(new_n580), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(G295));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n939), .ZN(G331));
  OAI21_X1  g516(.A(G286), .B1(G171), .B2(KEYINPUT103), .ZN(new_n942));
  OR2_X1    g517(.A1(new_n942), .A2(KEYINPUT104), .ZN(new_n943));
  NAND2_X1  g518(.A1(G171), .A2(KEYINPUT103), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(KEYINPUT104), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n944), .B1(new_n943), .B2(new_n945), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n947), .A2(new_n948), .A3(new_n860), .ZN(new_n949));
  INV_X1    g524(.A(new_n860), .ZN(new_n950));
  INV_X1    g525(.A(new_n945), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n942), .A2(KEYINPUT104), .ZN(new_n952));
  OAI211_X1 g527(.A(KEYINPUT103), .B(G171), .C1(new_n951), .C2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n950), .B1(new_n953), .B2(new_n946), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n909), .B1(new_n949), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n860), .B1(new_n947), .B2(new_n948), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n953), .A2(new_n950), .A3(new_n946), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n956), .A2(new_n915), .A3(new_n912), .A4(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n955), .A2(new_n958), .A3(new_n933), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n863), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT105), .ZN(new_n961));
  INV_X1    g536(.A(new_n932), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n961), .B1(new_n962), .B2(new_n930), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n931), .A2(KEYINPUT105), .A3(new_n932), .ZN(new_n964));
  AOI22_X1  g539(.A1(new_n955), .A2(new_n958), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT43), .B1(new_n960), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n913), .A2(new_n914), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n956), .A2(new_n967), .A3(new_n957), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n955), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n963), .A2(new_n964), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n971), .A2(new_n972), .A3(new_n863), .A4(new_n959), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n966), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n972), .B1(new_n960), .B2(new_n965), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n971), .A2(KEYINPUT43), .A3(new_n863), .A4(new_n959), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  MUX2_X1   g552(.A(new_n974), .B(new_n977), .S(KEYINPUT44), .Z(G397));
  INV_X1    g553(.A(G1384), .ZN(new_n979));
  INV_X1    g554(.A(new_n479), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n980), .B1(new_n488), .B2(G126), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n484), .B1(new_n981), .B2(new_n457), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n487), .A2(new_n489), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n979), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n462), .A2(new_n463), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(G2105), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n465), .A2(new_n466), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n457), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n986), .A2(new_n988), .A3(G40), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT106), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(G160), .A2(KEYINPUT106), .A3(G40), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n984), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G8), .ZN(new_n994));
  INV_X1    g569(.A(G1976), .ZN(new_n995));
  NOR2_X1   g570(.A1(G288), .A2(new_n995), .ZN(new_n996));
  NOR3_X1   g571(.A1(new_n993), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n999));
  NAND2_X1  g574(.A1(G288), .A2(new_n995), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n997), .A2(new_n998), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G1981), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n568), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(G1981), .B1(new_n564), .B2(new_n567), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT49), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n993), .A2(new_n994), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1003), .A2(KEYINPUT49), .A3(new_n1004), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n983), .ZN(new_n1011));
  AOI22_X1  g586(.A1(new_n481), .A2(G2105), .B1(G102), .B2(new_n483), .ZN(new_n1012));
  AOI21_X1  g587(.A(G1384), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT106), .B1(G160), .B2(G40), .ZN(new_n1014));
  INV_X1    g589(.A(G40), .ZN(new_n1015));
  NOR4_X1   g590(.A1(new_n464), .A2(new_n467), .A3(new_n990), .A4(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1013), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n996), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1017), .A2(G8), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT110), .B1(new_n1019), .B2(KEYINPUT52), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1017), .A2(new_n999), .A3(G8), .A4(new_n1018), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1000), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1001), .B(new_n1010), .C1(new_n1020), .C2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G2090), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT50), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n984), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n490), .A2(KEYINPUT50), .A3(new_n979), .ZN(new_n1028));
  AOI22_X1  g603(.A1(new_n1027), .A2(new_n1028), .B1(new_n992), .B2(new_n991), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n991), .A2(new_n992), .ZN(new_n1030));
  OAI211_X1 g605(.A(KEYINPUT45), .B(new_n979), .C1(new_n982), .C2(new_n983), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT45), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n984), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1030), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G1971), .ZN(new_n1035));
  AOI22_X1  g610(.A1(new_n1025), .A2(new_n1029), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1037), .B1(G303), .B2(G8), .ZN(new_n1038));
  NOR3_X1   g613(.A1(G166), .A2(KEYINPUT55), .A3(new_n994), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT109), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(G303), .A2(new_n1037), .A3(G8), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT55), .B1(G166), .B2(new_n994), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT109), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1040), .A2(new_n1044), .ZN(new_n1045));
  NOR3_X1   g620(.A1(new_n1036), .A2(new_n1045), .A3(new_n994), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1024), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT112), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1029), .A2(new_n1025), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n994), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1048), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1052), .ZN(new_n1054));
  OAI211_X1 g629(.A(KEYINPUT112), .B(new_n1054), .C1(new_n1036), .C2(new_n994), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G2084), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1029), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G1966), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1034), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1058), .A2(new_n1060), .A3(G168), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(G8), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT51), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT51), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1065), .B1(new_n1066), .B2(G286), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1067), .A2(new_n1062), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1047), .B(new_n1056), .C1(new_n1064), .C2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G2067), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1030), .A2(new_n1070), .A3(new_n1013), .ZN(new_n1071));
  OAI211_X1 g646(.A(KEYINPUT60), .B(new_n1071), .C1(new_n1029), .C2(G1348), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(new_n597), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n1030), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n1077), .A2(new_n697), .B1(new_n1070), .B2(new_n993), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1078), .A2(KEYINPUT117), .A3(KEYINPUT60), .A4(new_n612), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n1072), .B2(new_n597), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1072), .A2(new_n597), .A3(KEYINPUT118), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1075), .A2(new_n1079), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  OR2_X1    g658(.A1(new_n1078), .A2(KEYINPUT60), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT56), .B(G2072), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1030), .A2(new_n1033), .A3(new_n1031), .A4(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1088), .B1(new_n1029), .B2(G1956), .ZN(new_n1089));
  XNOR2_X1  g664(.A(G299), .B(KEYINPUT57), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n601), .B(KEYINPUT57), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1092), .B(new_n1088), .C1(G1956), .C2(new_n1029), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT61), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1086), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1091), .A2(new_n1093), .A3(KEYINPUT116), .A4(KEYINPUT61), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  XNOR2_X1  g673(.A(KEYINPUT58), .B(G1341), .ZN(new_n1099));
  OAI22_X1  g674(.A1(new_n1034), .A2(G1996), .B1(new_n993), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n537), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT59), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1100), .A2(new_n1103), .A3(new_n537), .ZN(new_n1104));
  AOI22_X1  g679(.A1(new_n1094), .A2(new_n1095), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1085), .A2(new_n1098), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1078), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1107), .A2(new_n597), .A3(new_n1093), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1108), .A2(new_n1091), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1069), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(G1961), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1077), .A2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1030), .A2(new_n1033), .A3(new_n753), .A4(new_n1031), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT119), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT53), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1112), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(KEYINPUT120), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT121), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT53), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1113), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1119), .B1(new_n1113), .B2(new_n1120), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT120), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1125), .B(new_n1112), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1118), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(G301), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1015), .B1(new_n988), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1130), .B(new_n1131), .C1(new_n1129), .C2(G160), .ZN(new_n1132));
  AND4_X1   g707(.A1(KEYINPUT53), .A2(new_n1132), .A3(new_n753), .A4(new_n1031), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT45), .B1(new_n490), .B2(new_n979), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1130), .B1(new_n1129), .B2(G160), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1134), .B1(KEYINPUT123), .B2(new_n1135), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n1133), .A2(new_n1136), .B1(new_n1077), .B2(new_n1111), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1137), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(KEYINPUT124), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT124), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1137), .B(new_n1140), .C1(new_n1122), .C2(new_n1121), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1139), .A2(G171), .A3(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1128), .A2(KEYINPUT54), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1127), .A2(G171), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1138), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT54), .B1(new_n1145), .B2(G301), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1143), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1110), .A2(new_n1148), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1010), .A2(new_n995), .A3(new_n797), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n1003), .B(KEYINPUT111), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1008), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1046), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1152), .B1(new_n1024), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT62), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1155), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1063), .B(KEYINPUT62), .C1(new_n1062), .C2(new_n1067), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1144), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1047), .A2(new_n1056), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1154), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1031), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1134), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(G1966), .B1(new_n1162), .B2(new_n1030), .ZN(new_n1163));
  AOI221_X4 g738(.A(G2084), .B1(new_n991), .B2(new_n992), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1164));
  OAI211_X1 g739(.A(G8), .B(G168), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(KEYINPUT113), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT113), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1066), .A2(new_n1167), .A3(G8), .A4(G168), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1047), .A2(new_n1169), .A3(new_n1056), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT63), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(KEYINPUT114), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT114), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1170), .A2(new_n1174), .A3(new_n1171), .ZN(new_n1175));
  OR2_X1    g750(.A1(new_n1051), .A2(KEYINPUT115), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1051), .A2(KEYINPUT115), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1176), .A2(new_n1054), .A3(new_n1177), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1178), .A2(KEYINPUT63), .A3(new_n1047), .A4(new_n1169), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1173), .A2(new_n1175), .A3(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1149), .A2(new_n1160), .A3(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(new_n830), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1182), .A2(new_n832), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n730), .A2(G2067), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n728), .A2(new_n1070), .A3(new_n729), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1186), .B(KEYINPUT108), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1182), .A2(new_n832), .ZN(new_n1188));
  INV_X1    g763(.A(G1996), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n766), .B(new_n1189), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1187), .A2(new_n1188), .A3(new_n1190), .ZN(new_n1191));
  NOR2_X1   g766(.A1(G290), .A2(G1986), .ZN(new_n1192));
  XNOR2_X1  g767(.A(new_n1192), .B(KEYINPUT107), .ZN(new_n1193));
  AND2_X1   g768(.A1(G290), .A2(G1986), .ZN(new_n1194));
  OR4_X1    g769(.A1(new_n1183), .A2(new_n1191), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1033), .B1(new_n992), .B2(new_n991), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1181), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1196), .A2(new_n1189), .ZN(new_n1199));
  XOR2_X1   g774(.A(new_n1199), .B(KEYINPUT46), .Z(new_n1200));
  NAND2_X1  g775(.A1(new_n1187), .A2(new_n767), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1200), .B1(new_n1201), .B2(new_n1196), .ZN(new_n1202));
  XOR2_X1   g777(.A(new_n1202), .B(KEYINPUT47), .Z(new_n1203));
  XNOR2_X1  g778(.A(new_n1183), .B(KEYINPUT125), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1187), .A2(new_n1190), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1185), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1206), .A2(new_n1196), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1196), .B1(new_n1191), .B2(new_n1183), .ZN(new_n1208));
  OR2_X1    g783(.A1(new_n1208), .A2(KEYINPUT126), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1208), .A2(KEYINPUT126), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1193), .A2(new_n1196), .ZN(new_n1211));
  XNOR2_X1  g786(.A(new_n1211), .B(KEYINPUT48), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1209), .A2(new_n1210), .A3(new_n1212), .ZN(new_n1213));
  AND3_X1   g788(.A1(new_n1203), .A2(new_n1207), .A3(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1198), .A2(new_n1214), .ZN(G329));
  assign    G231 = 1'b0;
  AND3_X1   g790(.A1(new_n690), .A2(new_n664), .A3(new_n691), .ZN(new_n1217));
  AND2_X1   g791(.A1(new_n649), .A2(G319), .ZN(new_n1218));
  AOI21_X1  g792(.A(KEYINPUT127), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g793(.A(new_n1219), .B1(new_n966), .B2(new_n973), .ZN(new_n1220));
  NAND2_X1  g794(.A1(new_n898), .A2(new_n902), .ZN(new_n1221));
  NAND3_X1  g795(.A1(new_n1217), .A2(KEYINPUT127), .A3(new_n1218), .ZN(new_n1222));
  AND3_X1   g796(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .ZN(G308));
  NAND3_X1  g797(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .ZN(G225));
endmodule


