//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 0 1 0 1 0 0 1 1 1 1 1 0 0 1 0 1 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 1 1 1 0 1 0 1 0 0 0 0 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970;
  NOR2_X1   g000(.A1(G237), .A2(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G210), .ZN(new_n188));
  INV_X1    g002(.A(G101), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n188), .B(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT28), .ZN(new_n193));
  XOR2_X1   g007(.A(KEYINPUT2), .B(G113), .Z(new_n194));
  XNOR2_X1  g008(.A(G116), .B(G119), .ZN(new_n195));
  AND2_X1   g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n194), .A2(new_n195), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G143), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  AND3_X1   g016(.A1(new_n202), .A2(KEYINPUT65), .A3(G146), .ZN(new_n203));
  AOI21_X1  g017(.A(KEYINPUT65), .B1(new_n202), .B2(G146), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n201), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT0), .ZN(new_n206));
  INV_X1    g020(.A(G128), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT64), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT64), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n211), .B1(KEYINPUT0), .B2(G128), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n205), .A2(new_n209), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n202), .A2(G146), .ZN(new_n215));
  AND2_X1   g029(.A1(new_n201), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(new_n208), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT11), .ZN(new_n219));
  INV_X1    g033(.A(G134), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n219), .B1(new_n220), .B2(G137), .ZN(new_n221));
  INV_X1    g035(.A(G137), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n222), .A2(KEYINPUT11), .A3(G134), .ZN(new_n223));
  INV_X1    g037(.A(G131), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n220), .A2(G137), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n221), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n227));
  XNOR2_X1  g041(.A(new_n226), .B(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n221), .A2(new_n225), .A3(new_n223), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n221), .A2(new_n223), .A3(KEYINPUT67), .A4(new_n225), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(G131), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n218), .B1(new_n228), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT1), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n201), .A2(new_n215), .A3(new_n235), .A4(G128), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n202), .A2(G146), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT65), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n238), .B1(new_n200), .B2(G143), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n202), .A2(KEYINPUT65), .A3(G146), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n237), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n207), .B1(new_n201), .B2(KEYINPUT1), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n236), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n225), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n220), .A2(G137), .ZN(new_n245));
  OAI21_X1  g059(.A(G131), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n226), .A2(new_n227), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n226), .A2(new_n227), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n243), .B(new_n246), .C1(new_n247), .C2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n199), .B1(new_n234), .B2(new_n250), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n229), .A2(new_n230), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n232), .A2(G131), .ZN(new_n253));
  OAI22_X1  g067(.A1(new_n247), .A2(new_n248), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n241), .A2(new_n208), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n255), .A2(new_n213), .B1(new_n208), .B2(new_n216), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(new_n198), .A3(new_n249), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n193), .B1(new_n251), .B2(new_n258), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n258), .A2(new_n193), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n192), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT30), .ZN(new_n262));
  AND3_X1   g076(.A1(new_n257), .A2(new_n262), .A3(new_n249), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n262), .B1(new_n257), .B2(new_n249), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n199), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n192), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n265), .A2(new_n258), .A3(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT31), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n261), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G472), .ZN(new_n270));
  INV_X1    g084(.A(G902), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n265), .A2(KEYINPUT31), .A3(new_n258), .A4(new_n266), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n269), .A2(new_n270), .A3(new_n271), .A4(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT32), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n272), .A2(new_n271), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT32), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n275), .A2(new_n276), .A3(new_n270), .A4(new_n269), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT68), .ZN(new_n279));
  INV_X1    g093(.A(new_n259), .ZN(new_n280));
  INV_X1    g094(.A(new_n260), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n266), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT29), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n265), .A2(new_n258), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n282), .B(new_n283), .C1(new_n284), .C2(new_n266), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n280), .A2(new_n281), .A3(KEYINPUT29), .A4(new_n266), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(new_n271), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G472), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n278), .A2(new_n279), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n279), .B1(new_n278), .B2(new_n288), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g105(.A(G110), .B(G140), .ZN(new_n292));
  INV_X1    g106(.A(G953), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n293), .A2(G227), .ZN(new_n294));
  XOR2_X1   g108(.A(new_n292), .B(new_n294), .Z(new_n295));
  NOR2_X1   g109(.A1(new_n295), .A2(KEYINPUT74), .ZN(new_n296));
  INV_X1    g110(.A(G107), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G104), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT75), .B(G107), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n298), .B1(new_n299), .B2(G104), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G101), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT3), .ZN(new_n302));
  AND2_X1   g116(.A1(KEYINPUT75), .A2(G107), .ZN(new_n303));
  NOR2_X1   g117(.A1(KEYINPUT75), .A2(G107), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n302), .B(G104), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n298), .A2(KEYINPUT3), .ZN(new_n306));
  INV_X1    g120(.A(G104), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G107), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n305), .A2(new_n189), .A3(new_n306), .A4(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n301), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n242), .ZN(new_n311));
  AND3_X1   g125(.A1(new_n201), .A2(new_n215), .A3(G128), .ZN(new_n312));
  AOI22_X1  g126(.A1(new_n205), .A2(new_n311), .B1(new_n312), .B2(new_n235), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT77), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n310), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n236), .B1(new_n216), .B2(new_n242), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n301), .A2(new_n309), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT77), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n243), .B1(new_n309), .B2(new_n301), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n254), .B(new_n315), .C1(new_n318), .C2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT12), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n301), .A2(new_n309), .ZN(new_n323));
  OAI211_X1 g137(.A(KEYINPUT77), .B(new_n317), .C1(new_n323), .C2(new_n243), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n324), .A2(KEYINPUT12), .A3(new_n254), .A4(new_n315), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT10), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n310), .A2(new_n313), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n305), .A2(new_n306), .A3(new_n308), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G101), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(KEYINPUT4), .A3(new_n309), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT4), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n329), .A2(new_n332), .A3(G101), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n331), .A2(new_n256), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n328), .B1(new_n334), .B2(KEYINPUT76), .ZN(new_n335));
  INV_X1    g149(.A(new_n254), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n317), .A2(new_n327), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT76), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n331), .A2(new_n256), .A3(new_n338), .A4(new_n333), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n335), .A2(new_n336), .A3(new_n337), .A4(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n296), .B1(new_n326), .B2(new_n340), .ZN(new_n341));
  AND2_X1   g155(.A1(new_n295), .A2(KEYINPUT74), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n335), .A2(new_n337), .A3(new_n339), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n254), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(new_n295), .A3(new_n340), .ZN(new_n347));
  AOI21_X1  g161(.A(G902), .B1(new_n344), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(new_n350), .A3(G469), .ZN(new_n351));
  INV_X1    g165(.A(G469), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n295), .B1(new_n346), .B2(new_n340), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n326), .A2(new_n340), .A3(new_n295), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n352), .B(new_n271), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  OAI211_X1 g169(.A(KEYINPUT78), .B(new_n355), .C1(new_n348), .C2(new_n352), .ZN(new_n356));
  XOR2_X1   g170(.A(KEYINPUT9), .B(G234), .Z(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(G221), .B1(new_n358), .B2(G902), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n351), .A2(new_n356), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n331), .A2(new_n199), .A3(new_n333), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n195), .A2(KEYINPUT5), .ZN(new_n362));
  INV_X1    g176(.A(G116), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n363), .A2(KEYINPUT5), .A3(G119), .ZN(new_n364));
  INV_X1    g178(.A(G113), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI22_X1  g180(.A1(new_n362), .A2(new_n366), .B1(new_n194), .B2(new_n195), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n323), .A2(KEYINPUT79), .A3(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(new_n301), .A3(new_n309), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT79), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n361), .A2(new_n368), .A3(new_n371), .ZN(new_n372));
  XOR2_X1   g186(.A(G110), .B(G122), .Z(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n373), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n361), .A2(new_n368), .A3(new_n375), .A4(new_n371), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n374), .A2(KEYINPUT6), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT6), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n372), .A2(new_n378), .A3(new_n373), .ZN(new_n379));
  INV_X1    g193(.A(G125), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n243), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n381), .B1(new_n218), .B2(new_n380), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n293), .A2(G224), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n382), .B(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n377), .A2(new_n379), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(KEYINPUT7), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n382), .B(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n310), .A2(new_n367), .ZN(new_n388));
  XOR2_X1   g202(.A(new_n373), .B(KEYINPUT8), .Z(new_n389));
  XNOR2_X1  g203(.A(new_n362), .B(KEYINPUT80), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n196), .B1(new_n390), .B2(new_n366), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n388), .B(new_n389), .C1(new_n391), .C2(new_n310), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n387), .A2(new_n392), .A3(new_n376), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n385), .A2(new_n271), .A3(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(G210), .B1(G237), .B2(G902), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n385), .A2(new_n271), .A3(new_n395), .A4(new_n393), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(G214), .B1(G237), .B2(G902), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(G140), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G125), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n380), .A2(G140), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT70), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n406), .B1(new_n405), .B2(new_n403), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT82), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT82), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n406), .B(new_n409), .C1(new_n405), .C2(new_n403), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n200), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(G125), .B(G140), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT72), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n412), .B(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n414), .A2(G146), .ZN(new_n415));
  INV_X1    g229(.A(G237), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(new_n293), .A3(G214), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n202), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n187), .A2(G143), .A3(G214), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(KEYINPUT18), .A2(G131), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n420), .A2(new_n421), .ZN(new_n423));
  OAI22_X1  g237(.A1(new_n411), .A2(new_n415), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT16), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(new_n402), .A3(G125), .ZN(new_n426));
  NOR3_X1   g240(.A1(new_n405), .A2(new_n380), .A3(G140), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n427), .B1(new_n405), .B2(new_n412), .ZN(new_n428));
  OAI211_X1 g242(.A(G146), .B(new_n426), .C1(new_n428), .C2(new_n425), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT71), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n428), .A2(new_n425), .ZN(new_n431));
  INV_X1    g245(.A(new_n426), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n200), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n407), .A2(KEYINPUT16), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT71), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n434), .A2(new_n435), .A3(G146), .A4(new_n426), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n430), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n420), .A2(KEYINPUT17), .A3(G131), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n420), .A2(G131), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n418), .A2(new_n224), .A3(new_n419), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n438), .B1(new_n441), .B2(KEYINPUT17), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n424), .B1(new_n437), .B2(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(G113), .B(G122), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n444), .B(new_n307), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n445), .B(new_n424), .C1(new_n437), .C2(new_n442), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n271), .ZN(new_n450));
  AND2_X1   g264(.A1(new_n450), .A2(G475), .ZN(new_n451));
  NOR2_X1   g265(.A1(G475), .A2(G902), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n429), .A2(new_n441), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n408), .A2(KEYINPUT19), .A3(new_n410), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT19), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n414), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n453), .B1(new_n457), .B2(new_n200), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n422), .A2(new_n423), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n408), .A2(new_n410), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(G146), .ZN(new_n461));
  INV_X1    g275(.A(new_n415), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n446), .B1(new_n458), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n464), .A2(KEYINPUT83), .A3(new_n448), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(KEYINPUT83), .B1(new_n464), .B2(new_n448), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n452), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(KEYINPUT81), .B(KEYINPUT20), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n464), .A2(new_n448), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT20), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(new_n472), .A3(new_n452), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n451), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n357), .A2(G217), .A3(new_n293), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  XOR2_X1   g290(.A(G116), .B(G122), .Z(new_n477));
  NOR2_X1   g291(.A1(new_n303), .A2(new_n304), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(G116), .B(G122), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n299), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(G128), .B(G143), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n220), .B1(new_n483), .B2(KEYINPUT13), .ZN(new_n484));
  OR3_X1    g298(.A1(new_n207), .A2(KEYINPUT13), .A3(G143), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n483), .A2(new_n220), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n482), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT84), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n484), .A2(new_n485), .B1(new_n220), .B2(new_n483), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT84), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n491), .A3(new_n482), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  XOR2_X1   g307(.A(G128), .B(G143), .Z(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(G134), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n487), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n363), .A2(KEYINPUT14), .A3(G122), .ZN(new_n497));
  OAI211_X1 g311(.A(G107), .B(new_n497), .C1(new_n477), .C2(KEYINPUT14), .ZN(new_n498));
  AND3_X1   g312(.A1(new_n496), .A2(new_n481), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n476), .B1(new_n493), .B2(new_n500), .ZN(new_n501));
  AOI211_X1 g315(.A(new_n475), .B(new_n499), .C1(new_n489), .C2(new_n492), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n271), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(KEYINPUT85), .ZN(new_n504));
  INV_X1    g318(.A(G478), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n505), .A2(KEYINPUT15), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT85), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n507), .B(new_n271), .C1(new_n501), .C2(new_n502), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n504), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  OR2_X1    g323(.A1(new_n503), .A2(new_n506), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n293), .A2(G952), .ZN(new_n513));
  NAND2_X1  g327(.A1(G234), .A2(G237), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XOR2_X1   g329(.A(KEYINPUT21), .B(G898), .Z(new_n516));
  NAND3_X1  g330(.A1(new_n514), .A2(G902), .A3(G953), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n474), .A2(new_n512), .A3(new_n518), .ZN(new_n519));
  NOR3_X1   g333(.A1(new_n360), .A2(new_n401), .A3(new_n519), .ZN(new_n520));
  XOR2_X1   g334(.A(KEYINPUT24), .B(G110), .Z(new_n521));
  XNOR2_X1  g335(.A(G119), .B(G128), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT69), .ZN(new_n524));
  INV_X1    g338(.A(G119), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n524), .B1(new_n525), .B2(G128), .ZN(new_n526));
  OR2_X1    g340(.A1(new_n526), .A2(KEYINPUT23), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(KEYINPUT23), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n527), .B(new_n528), .C1(G119), .C2(new_n207), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(G110), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n437), .A2(new_n523), .A3(new_n530), .ZN(new_n531));
  OAI22_X1  g345(.A1(new_n529), .A2(G110), .B1(new_n522), .B2(new_n521), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n462), .A2(new_n532), .A3(new_n429), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n293), .A2(G221), .A3(G234), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n534), .B(G137), .ZN(new_n535));
  XNOR2_X1  g349(.A(KEYINPUT73), .B(KEYINPUT22), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n535), .B(new_n536), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n531), .A2(new_n533), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n537), .B1(new_n531), .B2(new_n533), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n271), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(KEYINPUT25), .ZN(new_n541));
  INV_X1    g355(.A(G217), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n542), .B1(G234), .B2(new_n271), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT25), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n544), .B(new_n271), .C1(new_n538), .C2(new_n539), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n541), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  OR2_X1    g360(.A1(new_n540), .A2(new_n543), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n291), .A2(new_n520), .A3(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(G101), .ZN(G3));
  AND2_X1   g365(.A1(new_n273), .A2(KEYINPUT86), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n270), .B1(new_n275), .B2(new_n269), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n552), .B(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n360), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n555), .A2(new_n556), .A3(new_n549), .ZN(new_n557));
  XOR2_X1   g371(.A(new_n557), .B(KEYINPUT87), .Z(new_n558));
  NAND3_X1  g372(.A1(new_n397), .A2(KEYINPUT88), .A3(new_n398), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT88), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n394), .A2(new_n560), .A3(new_n396), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n559), .A2(new_n400), .A3(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n452), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT83), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n471), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n564), .B1(new_n566), .B2(new_n465), .ZN(new_n567));
  INV_X1    g381(.A(new_n469), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n473), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n451), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n504), .A2(new_n508), .ZN(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT90), .B(G478), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NOR3_X1   g388(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT33), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT33), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n490), .A2(new_n491), .A3(new_n482), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n491), .B1(new_n490), .B2(new_n482), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n500), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n475), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n493), .A2(new_n500), .A3(new_n476), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n576), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OAI211_X1 g396(.A(G478), .B(new_n271), .C1(new_n575), .C2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT89), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(KEYINPUT33), .B1(new_n501), .B2(new_n502), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n580), .A2(new_n576), .A3(new_n581), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n505), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(KEYINPUT89), .B1(new_n588), .B2(new_n271), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n574), .B1(new_n585), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n571), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n518), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n563), .A2(new_n593), .ZN(new_n594));
  XOR2_X1   g408(.A(KEYINPUT34), .B(G104), .Z(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(G6));
  NAND2_X1  g410(.A1(new_n567), .A2(new_n568), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n470), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n598), .A2(new_n511), .A3(new_n570), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n599), .A2(new_n592), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n563), .A2(new_n600), .ZN(new_n601));
  XOR2_X1   g415(.A(KEYINPUT35), .B(G107), .Z(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G9));
  AND3_X1   g417(.A1(new_n541), .A2(new_n543), .A3(new_n545), .ZN(new_n604));
  INV_X1    g418(.A(new_n543), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n537), .A2(KEYINPUT36), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n531), .A2(new_n533), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n607), .B1(new_n531), .B2(new_n533), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n271), .B(new_n605), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(KEYINPUT91), .ZN(new_n612));
  INV_X1    g426(.A(new_n610), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n608), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT91), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n614), .A2(new_n615), .A3(new_n271), .A4(new_n605), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(KEYINPUT92), .B1(new_n604), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT92), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n546), .A2(new_n619), .A3(new_n612), .A4(new_n616), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n520), .A2(new_n555), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(G110), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT93), .B(KEYINPUT37), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G12));
  NAND2_X1  g439(.A1(new_n618), .A2(new_n620), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n289), .A2(new_n290), .A3(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n562), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n515), .B1(new_n517), .B2(G900), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n351), .A2(new_n356), .A3(new_n359), .A4(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n630), .A2(new_n599), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n627), .A2(new_n628), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G128), .ZN(G30));
  XOR2_X1   g447(.A(new_n629), .B(KEYINPUT39), .Z(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n556), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(new_n636), .B(KEYINPUT40), .Z(new_n637));
  NAND3_X1  g451(.A1(new_n571), .A2(new_n400), .A3(new_n511), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n621), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT95), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n284), .A2(new_n192), .ZN(new_n641));
  AND3_X1   g455(.A1(new_n251), .A2(new_n258), .A3(new_n192), .ZN(new_n642));
  OR3_X1    g456(.A1(new_n641), .A2(KEYINPUT94), .A3(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(KEYINPUT94), .B1(new_n641), .B2(new_n642), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n643), .A2(new_n271), .A3(new_n644), .ZN(new_n645));
  AOI22_X1  g459(.A1(new_n645), .A2(G472), .B1(new_n274), .B2(new_n277), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n399), .B(KEYINPUT38), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n637), .A2(new_n640), .A3(new_n647), .A4(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G143), .ZN(G45));
  NAND2_X1  g464(.A1(new_n583), .A2(new_n584), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n588), .A2(KEYINPUT89), .A3(new_n271), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n653), .A2(new_n574), .B1(new_n569), .B2(new_n570), .ZN(new_n654));
  INV_X1    g468(.A(new_n630), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n627), .A2(new_n654), .A3(new_n628), .A4(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G146), .ZN(G48));
  NOR3_X1   g471(.A1(new_n289), .A2(new_n290), .A3(new_n548), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n271), .B1(new_n353), .B2(new_n354), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(G469), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n660), .A2(new_n355), .A3(new_n359), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n562), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n658), .A2(new_n593), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT41), .B(G113), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G15));
  NAND3_X1  g479(.A1(new_n658), .A2(new_n600), .A3(new_n662), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G116), .ZN(G18));
  INV_X1    g481(.A(new_n519), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n627), .A2(KEYINPUT96), .A3(new_n668), .A4(new_n662), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT96), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n278), .A2(new_n288), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(KEYINPUT68), .ZN(new_n672));
  AOI22_X1  g486(.A1(new_n274), .A2(new_n277), .B1(new_n287), .B2(G472), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n279), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n672), .A2(new_n662), .A3(new_n621), .A4(new_n674), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n670), .B1(new_n675), .B2(new_n519), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n669), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G119), .ZN(G21));
  NAND2_X1  g492(.A1(new_n559), .A2(new_n561), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n638), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n661), .ZN(new_n681));
  INV_X1    g495(.A(new_n273), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n548), .A2(new_n682), .A3(new_n553), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n680), .A2(new_n518), .A3(new_n681), .A4(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G122), .ZN(G24));
  NOR2_X1   g499(.A1(new_n682), .A2(new_n553), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n618), .A2(new_n686), .A3(new_n620), .ZN(new_n687));
  AOI21_X1  g501(.A(KEYINPUT97), .B1(new_n654), .B2(new_n629), .ZN(new_n688));
  AOI22_X1  g502(.A1(new_n651), .A2(new_n652), .B1(new_n572), .B2(new_n573), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT97), .ZN(new_n690));
  INV_X1    g504(.A(new_n629), .ZN(new_n691));
  NOR4_X1   g505(.A1(new_n474), .A2(new_n689), .A3(new_n690), .A4(new_n691), .ZN(new_n692));
  OAI211_X1 g506(.A(new_n687), .B(new_n662), .C1(new_n688), .C2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G125), .ZN(G27));
  NAND3_X1  g508(.A1(new_n571), .A2(new_n590), .A3(new_n629), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n690), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n571), .A2(new_n590), .A3(KEYINPUT97), .A4(new_n629), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n348), .A2(new_n352), .ZN(new_n699));
  INV_X1    g513(.A(new_n355), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n359), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n397), .A2(new_n400), .A3(new_n398), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT42), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n673), .A2(new_n704), .A3(new_n548), .ZN(new_n705));
  AND3_X1   g519(.A1(new_n698), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n291), .A2(new_n549), .A3(new_n698), .A4(new_n703), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n706), .B1(new_n707), .B2(new_n704), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(new_n224), .ZN(G33));
  NAND4_X1  g523(.A1(new_n672), .A2(new_n703), .A3(new_n674), .A4(new_n549), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n710), .A2(new_n599), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n629), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G134), .ZN(G36));
  AOI21_X1  g527(.A(KEYINPUT100), .B1(new_n474), .B2(new_n590), .ZN(new_n714));
  XOR2_X1   g528(.A(new_n714), .B(KEYINPUT43), .Z(new_n715));
  INV_X1    g529(.A(new_n555), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n715), .A2(new_n716), .A3(new_n621), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(KEYINPUT101), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n702), .B1(new_n717), .B2(new_n718), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n344), .A2(new_n347), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT45), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n352), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  OR2_X1    g538(.A1(new_n724), .A2(KEYINPUT98), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(KEYINPUT98), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n725), .B(new_n726), .C1(new_n723), .C2(new_n722), .ZN(new_n727));
  NAND2_X1  g541(.A1(G469), .A2(G902), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n727), .A2(KEYINPUT46), .A3(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT99), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n729), .A2(new_n730), .A3(new_n355), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n730), .B1(new_n729), .B2(new_n355), .ZN(new_n732));
  AOI21_X1  g546(.A(KEYINPUT46), .B1(new_n727), .B2(new_n728), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(new_n359), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n720), .A2(new_n635), .A3(new_n721), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G137), .ZN(G39));
  XNOR2_X1  g552(.A(new_n736), .B(KEYINPUT47), .ZN(new_n739));
  INV_X1    g553(.A(new_n702), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n291), .A2(new_n695), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n739), .A2(new_n548), .A3(new_n740), .A4(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G140), .ZN(G42));
  AND3_X1   g557(.A1(new_n715), .A2(new_n514), .A3(new_n513), .ZN(new_n744));
  INV_X1    g558(.A(new_n400), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n745), .B1(KEYINPUT108), .B2(KEYINPUT50), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n648), .A2(new_n746), .ZN(new_n747));
  AND4_X1   g561(.A1(new_n681), .A2(new_n744), .A3(new_n683), .A4(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g563(.A(KEYINPUT108), .B1(KEYINPUT107), .B2(KEYINPUT50), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n748), .A2(new_n750), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT109), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n661), .A2(new_n702), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n744), .A2(new_n687), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n646), .A2(new_n756), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n758), .A2(new_n548), .A3(new_n515), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(new_n474), .A3(new_n689), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n755), .A2(new_n757), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n754), .B1(new_n752), .B2(new_n753), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n744), .A2(new_n683), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n660), .A2(new_n355), .ZN(new_n765));
  XOR2_X1   g579(.A(new_n765), .B(KEYINPUT106), .Z(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n359), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n740), .B(new_n764), .C1(new_n739), .C2(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(KEYINPUT51), .B1(new_n763), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n757), .A2(new_n760), .ZN(new_n770));
  OAI21_X1  g584(.A(KEYINPUT51), .B1(new_n770), .B2(KEYINPUT110), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n771), .B1(KEYINPUT110), .B2(new_n770), .ZN(new_n772));
  AND4_X1   g586(.A1(new_n768), .A2(new_n752), .A3(new_n753), .A4(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n673), .A2(new_n548), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n744), .A2(new_n774), .A3(new_n756), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT48), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n759), .A2(new_n654), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n777), .A2(new_n513), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n769), .A2(new_n773), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n764), .A2(new_n662), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n672), .A2(new_n674), .A3(new_n621), .A4(new_n628), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n783), .A2(new_n591), .A3(new_n630), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n630), .A2(new_n599), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n693), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n701), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n604), .A2(new_n617), .A3(new_n691), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n647), .A2(new_n680), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(KEYINPUT52), .B1(new_n787), .B2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n656), .A2(new_n632), .A3(new_n693), .A4(new_n790), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  AOI211_X1 g609(.A(new_n451), .B(new_n511), .C1(new_n470), .C2(new_n597), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n630), .A2(new_n702), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n291), .A2(new_n621), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n399), .A2(new_n400), .A3(new_n518), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n474), .A2(new_n511), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n799), .B1(new_n591), .B2(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n555), .A2(new_n801), .A3(new_n556), .A4(new_n549), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n798), .A2(new_n550), .A3(new_n622), .A4(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n708), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n698), .A2(new_n687), .A3(new_n703), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT103), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n698), .A2(KEYINPUT103), .A3(new_n687), .A4(new_n703), .ZN(new_n808));
  AOI22_X1  g622(.A1(new_n807), .A2(new_n808), .B1(new_n711), .B2(new_n629), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n663), .A2(new_n666), .ZN(new_n810));
  INV_X1    g624(.A(new_n684), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n811), .B1(new_n669), .B2(new_n676), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n804), .A2(new_n809), .A3(new_n810), .A4(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n795), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT53), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n816));
  XNOR2_X1  g630(.A(KEYINPUT105), .B(KEYINPUT53), .ZN(new_n817));
  OAI21_X1  g631(.A(KEYINPUT104), .B1(new_n791), .B2(new_n794), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n792), .A2(new_n793), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT104), .ZN(new_n820));
  INV_X1    g634(.A(new_n786), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n821), .A2(KEYINPUT52), .A3(new_n656), .A4(new_n790), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n819), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n813), .B1(new_n818), .B2(new_n823), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n815), .B(new_n816), .C1(new_n817), .C2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n824), .A2(new_n817), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n809), .A2(new_n812), .A3(new_n810), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n707), .A2(new_n704), .ZN(new_n829));
  INV_X1    g643(.A(new_n706), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n550), .A2(new_n622), .A3(new_n802), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n831), .A2(new_n832), .A3(new_n798), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n828), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n819), .A2(new_n822), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT53), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n816), .B1(new_n827), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n826), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n781), .A2(new_n782), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n841), .B1(G952), .B2(G953), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n647), .B1(KEYINPUT49), .B2(new_n765), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n474), .A2(new_n590), .A3(new_n400), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n844), .A2(new_n548), .A3(new_n735), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n845), .A2(KEYINPUT102), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(KEYINPUT102), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n765), .A2(KEYINPUT49), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n648), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n843), .A2(new_n846), .A3(new_n847), .A4(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n842), .A2(new_n850), .ZN(G75));
  INV_X1    g665(.A(KEYINPUT113), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n815), .B1(new_n817), .B2(new_n824), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(G902), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT112), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n853), .A2(KEYINPUT112), .A3(G902), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n852), .B1(new_n858), .B2(new_n395), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT56), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n377), .A2(new_n379), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(new_n384), .ZN(new_n862));
  XNOR2_X1  g676(.A(KEYINPUT111), .B(KEYINPUT55), .ZN(new_n863));
  XOR2_X1   g677(.A(new_n862), .B(new_n863), .Z(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n856), .A2(KEYINPUT113), .A3(new_n396), .A4(new_n857), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n859), .A2(new_n860), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  OR3_X1    g681(.A1(new_n293), .A2(KEYINPUT114), .A3(G952), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT114), .B1(new_n293), .B2(G952), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT115), .ZN(new_n871));
  INV_X1    g685(.A(G210), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n860), .B1(new_n854), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n871), .B1(new_n873), .B2(new_n864), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n867), .A2(new_n874), .ZN(G51));
  AND3_X1   g689(.A1(new_n819), .A2(new_n820), .A3(new_n822), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n820), .B1(new_n819), .B2(new_n822), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n834), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(new_n817), .ZN(new_n879));
  AOI22_X1  g693(.A1(new_n878), .A2(new_n879), .B1(new_n814), .B2(KEYINPUT53), .ZN(new_n880));
  OAI21_X1  g694(.A(KEYINPUT116), .B1(new_n880), .B2(new_n816), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT116), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n818), .A2(new_n823), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n817), .B1(new_n883), .B2(new_n834), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n836), .A2(new_n837), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n882), .B(KEYINPUT54), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n881), .A2(new_n825), .A3(new_n886), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n728), .B(KEYINPUT57), .Z(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n889), .B1(new_n353), .B2(new_n354), .ZN(new_n890));
  OR2_X1    g704(.A1(new_n858), .A2(new_n727), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n870), .B1(new_n890), .B2(new_n891), .ZN(G54));
  AND2_X1   g706(.A1(new_n856), .A2(new_n857), .ZN(new_n893));
  NAND2_X1  g707(.A1(KEYINPUT58), .A2(G475), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT117), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n896), .A2(new_n566), .A3(new_n465), .ZN(new_n897));
  INV_X1    g711(.A(new_n870), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n893), .B(new_n895), .C1(new_n467), .C2(new_n466), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(G60));
  NAND2_X1  g714(.A1(new_n586), .A2(new_n587), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(G478), .A2(G902), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT59), .Z(new_n904));
  NOR2_X1   g718(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n887), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT118), .ZN(new_n907));
  INV_X1    g721(.A(new_n904), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n908), .B1(new_n826), .B2(new_n839), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n871), .B1(new_n909), .B2(new_n902), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT118), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n887), .A2(new_n911), .A3(new_n905), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n907), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(KEYINPUT119), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT119), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n907), .A2(new_n915), .A3(new_n910), .A4(new_n912), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n914), .A2(new_n916), .ZN(G63));
  NAND2_X1  g731(.A1(G217), .A2(G902), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT121), .ZN(new_n919));
  XOR2_X1   g733(.A(KEYINPUT120), .B(KEYINPUT60), .Z(new_n920));
  XNOR2_X1  g734(.A(new_n919), .B(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n853), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n538), .A2(new_n539), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n871), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(KEYINPUT61), .B1(new_n924), .B2(KEYINPUT122), .ZN(new_n925));
  INV_X1    g739(.A(new_n614), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n924), .B1(new_n926), .B2(new_n922), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n925), .B(new_n927), .ZN(G66));
  AOI21_X1  g742(.A(new_n293), .B1(new_n516), .B2(G224), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n812), .A2(new_n810), .A3(new_n832), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n929), .B1(new_n930), .B2(new_n293), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n861), .B1(G898), .B2(new_n293), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n931), .B(new_n932), .Z(G69));
  NOR2_X1   g747(.A1(new_n293), .A2(G900), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT126), .Z(new_n935));
  NAND4_X1  g749(.A1(new_n736), .A2(new_n635), .A3(new_n680), .A4(new_n774), .ZN(new_n936));
  AND4_X1   g750(.A1(new_n831), .A2(new_n936), .A3(new_n712), .A4(new_n787), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n742), .A2(new_n737), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n935), .B1(new_n938), .B2(new_n293), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n263), .A2(new_n264), .ZN(new_n940));
  XNOR2_X1  g754(.A(KEYINPUT123), .B(KEYINPUT124), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(new_n457), .ZN(new_n943));
  OAI21_X1  g757(.A(KEYINPUT125), .B1(new_n939), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n293), .B1(G227), .B2(G900), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n649), .A2(new_n787), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT62), .Z(new_n949));
  INV_X1    g763(.A(new_n636), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n591), .A2(new_n800), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n950), .A2(new_n658), .A3(new_n740), .A4(new_n951), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n742), .A2(new_n737), .A3(new_n949), .A4(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n293), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n943), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n955), .B1(new_n943), .B2(new_n939), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n947), .B(new_n956), .ZN(G72));
  NAND2_X1  g771(.A1(G472), .A2(G902), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT63), .Z(new_n959));
  OAI21_X1  g773(.A(new_n959), .B1(new_n953), .B2(new_n930), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT127), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI211_X1 g776(.A(KEYINPUT127), .B(new_n959), .C1(new_n953), .C2(new_n930), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n962), .A2(new_n641), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n959), .B1(new_n938), .B2(new_n930), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n965), .A2(new_n284), .A3(new_n192), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n827), .A2(new_n838), .ZN(new_n967));
  INV_X1    g781(.A(new_n641), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n284), .A2(new_n192), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n967), .A2(new_n968), .A3(new_n959), .A4(new_n969), .ZN(new_n970));
  AND4_X1   g784(.A1(new_n898), .A2(new_n964), .A3(new_n966), .A4(new_n970), .ZN(G57));
endmodule


