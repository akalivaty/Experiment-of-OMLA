//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 0 0 1 0 0 0 1 1 1 0 1 1 0 0 1 1 0 1 1 1 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:05 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n550,
    new_n551, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n568, new_n569, new_n570, new_n571, new_n573, new_n574,
    new_n576, new_n577, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n623, new_n624, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT66), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  INV_X1    g035(.A(G137), .ZN(new_n461));
  OR2_X1    g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AND2_X1   g039(.A1(G101), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n460), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(G125), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n460), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n466), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI211_X1 g048(.A(KEYINPUT67), .B(new_n460), .C1(new_n469), .C2(new_n470), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n473), .A2(new_n474), .ZN(G160));
  NOR2_X1   g050(.A1(new_n467), .A2(new_n468), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n476), .A2(new_n460), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  OAI21_X1  g055(.A(KEYINPUT68), .B1(G100), .B2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NOR3_X1   g057(.A1(KEYINPUT68), .A2(G100), .A3(G2105), .ZN(new_n483));
  OAI221_X1 g058(.A(G2104), .B1(G112), .B2(new_n460), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n478), .A2(new_n480), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  OAI211_X1 g061(.A(G138), .B(new_n460), .C1(new_n467), .C2(new_n468), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n462), .A2(new_n463), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .A3(G138), .A4(new_n460), .ZN(new_n491));
  NAND2_X1  g066(.A1(G126), .A2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n493), .B1(new_n467), .B2(new_n468), .ZN(new_n494));
  INV_X1    g069(.A(G102), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(new_n460), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n496), .A2(new_n498), .A3(G2104), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n500));
  AND3_X1   g075(.A1(new_n494), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n500), .B1(new_n494), .B2(new_n499), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n489), .B(new_n491), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  NAND2_X1  g079(.A1(G75), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT5), .B1(new_n506), .B2(KEYINPUT70), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n508), .A2(new_n509), .A3(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G62), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n505), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT71), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT6), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n511), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n506), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n521), .A2(G88), .B1(new_n522), .B2(G50), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n515), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n514), .A2(KEYINPUT71), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(G166));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT6), .B(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n529), .A2(G51), .A3(G543), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n507), .A2(new_n510), .A3(G63), .A4(G651), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n528), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n532), .B1(G89), .B2(new_n521), .ZN(G168));
  NAND4_X1  g108(.A1(new_n529), .A2(G90), .A3(new_n507), .A4(new_n510), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n529), .A2(G52), .A3(G543), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n507), .A2(new_n510), .A3(G64), .ZN(new_n537));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n516), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(G171));
  NAND4_X1  g115(.A1(new_n529), .A2(G81), .A3(new_n507), .A4(new_n510), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n529), .A2(G43), .A3(G543), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n507), .A2(new_n510), .A3(G56), .ZN(new_n544));
  NAND2_X1  g119(.A1(G68), .A2(G543), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n516), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  NAND2_X1  g127(.A1(G78), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G65), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n511), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G651), .ZN(new_n556));
  INV_X1    g131(.A(G91), .ZN(new_n557));
  AND2_X1   g132(.A1(new_n507), .A2(new_n510), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(new_n529), .ZN(new_n559));
  AND2_X1   g134(.A1(G53), .A2(G543), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n529), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT72), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AND2_X1   g139(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n561), .A2(new_n564), .ZN(new_n566));
  OAI221_X1 g141(.A(new_n556), .B1(new_n557), .B2(new_n559), .C1(new_n565), .C2(new_n566), .ZN(G299));
  INV_X1    g142(.A(KEYINPUT73), .ZN(new_n568));
  NAND2_X1  g143(.A1(G171), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT73), .B1(new_n536), .B2(new_n539), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(G301));
  INV_X1    g147(.A(new_n532), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n521), .A2(G89), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(G286));
  OR3_X1    g150(.A1(new_n524), .A2(KEYINPUT74), .A3(new_n525), .ZN(new_n576));
  OAI21_X1  g151(.A(KEYINPUT74), .B1(new_n524), .B2(new_n525), .ZN(new_n577));
  AND2_X1   g152(.A1(new_n576), .A2(new_n577), .ZN(G303));
  NAND2_X1  g153(.A1(new_n522), .A2(G49), .ZN(new_n579));
  INV_X1    g154(.A(G87), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n559), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n558), .B2(G74), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n581), .A2(new_n583), .ZN(G288));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G61), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n511), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(G651), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n521), .A2(G86), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n522), .A2(G48), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(G305));
  XOR2_X1   g166(.A(KEYINPUT75), .B(G85), .Z(new_n592));
  AOI22_X1  g167(.A1(new_n521), .A2(new_n592), .B1(new_n522), .B2(G47), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n558), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n516), .B2(new_n594), .ZN(G290));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  INV_X1    g171(.A(G92), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n559), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n521), .A2(KEYINPUT10), .A3(G92), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n507), .A2(new_n510), .A3(G66), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G651), .ZN(new_n604));
  AND3_X1   g179(.A1(new_n529), .A2(G54), .A3(G543), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(KEYINPUT76), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n516), .B1(new_n601), .B2(new_n602), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT76), .ZN(new_n609));
  NOR3_X1   g184(.A1(new_n608), .A2(new_n605), .A3(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n600), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  MUX2_X1   g186(.A(new_n611), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g187(.A(new_n611), .B(G301), .S(G868), .Z(G321));
  INV_X1    g188(.A(KEYINPUT77), .ZN(new_n614));
  INV_X1    g189(.A(G868), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(G168), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g191(.A1(G286), .A2(KEYINPUT77), .A3(G868), .ZN(new_n617));
  OAI22_X1  g192(.A1(new_n565), .A2(new_n566), .B1(new_n559), .B2(new_n557), .ZN(new_n618));
  INV_X1    g193(.A(new_n556), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n616), .B(new_n617), .C1(G868), .C2(new_n620), .ZN(G297));
  OAI211_X1 g196(.A(new_n616), .B(new_n617), .C1(G868), .C2(new_n620), .ZN(G280));
  INV_X1    g197(.A(G860), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n611), .B1(G559), .B2(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT78), .Z(G148));
  OR2_X1    g200(.A1(new_n611), .A2(G559), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G868), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(G868), .B2(new_n547), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g204(.A1(new_n477), .A2(G2104), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n633), .A2(G2100), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(G2100), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n477), .A2(G135), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n479), .A2(G123), .ZN(new_n637));
  NOR2_X1   g212(.A1(G99), .A2(G2105), .ZN(new_n638));
  OAI21_X1  g213(.A(G2104), .B1(new_n460), .B2(G111), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n636), .B(new_n637), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(G2096), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n634), .A2(new_n635), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT80), .ZN(G156));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2443), .B(G2446), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(KEYINPUT15), .B(G2435), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2438), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2427), .B(G2430), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  AND2_X1   g229(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n652), .A2(new_n654), .ZN(new_n656));
  XOR2_X1   g231(.A(KEYINPUT81), .B(KEYINPUT14), .Z(new_n657));
  NOR3_X1   g232(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n650), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n650), .A2(new_n658), .ZN(new_n660));
  AND3_X1   g235(.A1(new_n659), .A2(G14), .A3(new_n660), .ZN(G401));
  XNOR2_X1  g236(.A(G2072), .B(G2078), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT82), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT17), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  NOR2_X1   g243(.A1(new_n665), .A2(new_n662), .ZN(new_n669));
  NOR3_X1   g244(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT83), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n668), .A2(new_n665), .A3(new_n662), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT18), .Z(new_n673));
  NAND3_X1  g248(.A1(new_n664), .A2(new_n666), .A3(new_n668), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n671), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(new_n641), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G2100), .ZN(G227));
  XOR2_X1   g252(.A(G1961), .B(G1966), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT84), .ZN(new_n679));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n681), .A2(KEYINPUT85), .ZN(new_n682));
  XOR2_X1   g257(.A(G1971), .B(G1976), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT19), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(KEYINPUT85), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n682), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT20), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n679), .A2(new_n680), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(new_n681), .B2(new_n684), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n684), .A2(KEYINPUT86), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT87), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n692), .B(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(G1981), .B(G1986), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1991), .B(G1996), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(G229));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G21), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(G168), .B2(new_n700), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT98), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n703), .A2(G1966), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n703), .A2(G1966), .ZN(new_n705));
  INV_X1    g280(.A(G28), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n706), .A2(KEYINPUT30), .ZN(new_n707));
  AOI21_X1  g282(.A(G29), .B1(new_n706), .B2(KEYINPUT30), .ZN(new_n708));
  OR2_X1    g283(.A1(KEYINPUT31), .A2(G11), .ZN(new_n709));
  NAND2_X1  g284(.A1(KEYINPUT31), .A2(G11), .ZN(new_n710));
  AOI22_X1  g285(.A1(new_n707), .A2(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NOR2_X1   g287(.A1(G171), .A2(new_n700), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(G5), .B2(new_n700), .ZN(new_n714));
  INV_X1    g289(.A(G1961), .ZN(new_n715));
  OAI221_X1 g290(.A(new_n711), .B1(new_n712), .B2(new_n640), .C1(new_n714), .C2(new_n715), .ZN(new_n716));
  NOR3_X1   g291(.A1(new_n704), .A2(new_n705), .A3(new_n716), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT99), .Z(new_n718));
  NAND2_X1  g293(.A1(new_n712), .A2(G32), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n479), .A2(G129), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT95), .ZN(new_n721));
  AND3_X1   g296(.A1(new_n460), .A2(G105), .A3(G2104), .ZN(new_n722));
  NAND3_X1  g297(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT26), .ZN(new_n724));
  AOI211_X1 g299(.A(new_n722), .B(new_n724), .C1(G141), .C2(new_n477), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT96), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n719), .B1(new_n727), .B2(new_n712), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT27), .B(G1996), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT24), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n712), .B1(new_n732), .B2(G34), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(KEYINPUT93), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n733), .A2(KEYINPUT93), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(new_n732), .B2(G34), .ZN(new_n736));
  AOI22_X1  g311(.A1(G160), .A2(G29), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT94), .Z(new_n738));
  INV_X1    g313(.A(G2084), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n712), .A2(G27), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G164), .B2(new_n712), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT100), .B(G2078), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n715), .B2(new_n714), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n731), .A2(new_n740), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n728), .A2(new_n730), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n738), .A2(new_n739), .ZN(new_n748));
  NAND2_X1  g323(.A1(G115), .A2(G2104), .ZN(new_n749));
  INV_X1    g324(.A(G127), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n749), .B1(new_n476), .B2(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n460), .B1(new_n751), .B2(KEYINPUT92), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(KEYINPUT92), .B2(new_n751), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT25), .ZN(new_n754));
  NAND2_X1  g329(.A1(G103), .A2(G2104), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n754), .B1(new_n755), .B2(G2105), .ZN(new_n756));
  NAND4_X1  g331(.A1(new_n460), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n477), .A2(G139), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n753), .A2(new_n758), .ZN(new_n759));
  MUX2_X1   g334(.A(G33), .B(new_n759), .S(G29), .Z(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G2072), .ZN(new_n761));
  NOR3_X1   g336(.A1(new_n747), .A2(new_n748), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n746), .B1(new_n762), .B2(KEYINPUT97), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n718), .B(new_n763), .C1(KEYINPUT97), .C2(new_n762), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT101), .ZN(new_n765));
  MUX2_X1   g340(.A(G23), .B(G288), .S(G16), .Z(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT89), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT33), .B(G1976), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(G16), .A2(G22), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G166), .B2(G16), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n772), .A2(G1971), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n767), .B2(new_n769), .ZN(new_n774));
  NOR2_X1   g349(.A1(G6), .A2(G16), .ZN(new_n775));
  INV_X1    g350(.A(G305), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(G16), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT32), .B(G1981), .Z(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n772), .A2(G1971), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n770), .A2(new_n774), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n781), .A2(KEYINPUT34), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(KEYINPUT34), .ZN(new_n783));
  MUX2_X1   g358(.A(G24), .B(G290), .S(G16), .Z(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(G1986), .Z(new_n785));
  INV_X1    g360(.A(KEYINPUT88), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n712), .A2(G25), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n477), .A2(G131), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n479), .A2(G119), .ZN(new_n791));
  OR2_X1    g366(.A1(G95), .A2(G2105), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n792), .B(G2104), .C1(G107), .C2(new_n460), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n790), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n789), .B1(new_n795), .B2(new_n712), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT35), .B(G1991), .Z(new_n797));
  XOR2_X1   g372(.A(new_n796), .B(new_n797), .Z(new_n798));
  NOR3_X1   g373(.A1(new_n787), .A2(new_n788), .A3(new_n798), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n782), .A2(new_n783), .A3(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT36), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n800), .B1(KEYINPUT90), .B2(new_n801), .ZN(new_n802));
  OR3_X1    g377(.A1(new_n800), .A2(KEYINPUT90), .A3(new_n801), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n712), .A2(G35), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G162), .B2(new_n712), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT29), .Z(new_n806));
  INV_X1    g381(.A(G2090), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT102), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n712), .A2(G26), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT91), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT28), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n477), .A2(G140), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n479), .A2(G128), .ZN(new_n814));
  OR2_X1    g389(.A1(G104), .A2(G2105), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n815), .B(G2104), .C1(G116), .C2(new_n460), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n813), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n812), .B1(new_n818), .B2(new_n712), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(G2067), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n700), .A2(G19), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n547), .B2(new_n700), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G1341), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n700), .A2(G20), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT23), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n620), .B2(new_n700), .ZN(new_n827));
  INV_X1    g402(.A(G1956), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n824), .B(new_n829), .C1(new_n807), .C2(new_n806), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n700), .A2(G4), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n604), .A2(new_n606), .A3(KEYINPUT76), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n609), .B1(new_n608), .B2(new_n605), .ZN(new_n833));
  AOI22_X1  g408(.A1(new_n832), .A2(new_n833), .B1(new_n598), .B2(new_n599), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n831), .B1(new_n834), .B2(new_n700), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(G1348), .ZN(new_n836));
  NOR3_X1   g411(.A1(new_n809), .A2(new_n830), .A3(new_n836), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n765), .A2(new_n802), .A3(new_n803), .A4(new_n837), .ZN(G150));
  INV_X1    g413(.A(G150), .ZN(G311));
  NAND4_X1  g414(.A1(new_n529), .A2(G93), .A3(new_n507), .A4(new_n510), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n529), .A2(G55), .A3(G543), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n507), .A2(new_n510), .A3(G67), .ZN(new_n843));
  NAND2_X1  g418(.A1(G80), .A2(G543), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n516), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT104), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(KEYINPUT104), .B1(new_n842), .B2(new_n845), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(G860), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT37), .Z(new_n852));
  NAND2_X1  g427(.A1(new_n834), .A2(G559), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT38), .Z(new_n854));
  INV_X1    g429(.A(new_n547), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n848), .A2(new_n855), .A3(new_n849), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT103), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n855), .B2(new_n846), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n843), .A2(new_n844), .ZN(new_n859));
  OAI211_X1 g434(.A(new_n841), .B(new_n840), .C1(new_n859), .C2(new_n516), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n860), .A2(KEYINPUT103), .A3(new_n547), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n856), .A2(new_n858), .A3(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n854), .B(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  AND2_X1   g439(.A1(new_n864), .A2(KEYINPUT39), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n623), .B1(new_n864), .B2(KEYINPUT39), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n852), .B1(new_n865), .B2(new_n866), .ZN(G145));
  MUX2_X1   g442(.A(new_n727), .B(new_n726), .S(new_n759), .Z(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n632), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n479), .A2(G130), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT105), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n477), .A2(G142), .ZN(new_n872));
  NOR2_X1   g447(.A1(G106), .A2(G2105), .ZN(new_n873));
  OAI21_X1  g448(.A(G2104), .B1(new_n460), .B2(G118), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n871), .B(new_n872), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n794), .ZN(new_n876));
  INV_X1    g451(.A(G2104), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n877), .B1(new_n497), .B2(G2105), .ZN(new_n878));
  AOI22_X1  g453(.A1(new_n490), .A2(new_n493), .B1(new_n878), .B2(new_n496), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n879), .A2(new_n489), .A3(new_n491), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n817), .B(new_n880), .Z(new_n881));
  XOR2_X1   g456(.A(new_n876), .B(new_n881), .Z(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n869), .B(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(G162), .B(new_n640), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(G160), .ZN(new_n886));
  AOI21_X1  g461(.A(G37), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT106), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n887), .B(new_n888), .C1(new_n886), .C2(new_n884), .ZN(new_n889));
  INV_X1    g464(.A(G37), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n869), .B(new_n882), .ZN(new_n891));
  INV_X1    g466(.A(new_n886), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n884), .A2(new_n886), .ZN(new_n894));
  OAI21_X1  g469(.A(KEYINPUT106), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n889), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g472(.A1(new_n850), .A2(new_n615), .ZN(new_n898));
  XNOR2_X1  g473(.A(G305), .B(KEYINPUT108), .ZN(new_n899));
  OR2_X1    g474(.A1(new_n899), .A2(G166), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(G166), .ZN(new_n901));
  XNOR2_X1  g476(.A(G288), .B(G290), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n902), .B1(new_n900), .B2(new_n901), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(KEYINPUT109), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(KEYINPUT42), .ZN(new_n908));
  XOR2_X1   g483(.A(new_n626), .B(new_n862), .Z(new_n909));
  INV_X1    g484(.A(KEYINPUT107), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n910), .B1(new_n834), .B2(G299), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n611), .A2(KEYINPUT107), .A3(new_n620), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n834), .A2(G299), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n909), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(KEYINPUT41), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT41), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n911), .A2(new_n912), .A3(new_n917), .A4(new_n913), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n915), .B1(new_n909), .B2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n908), .B(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n898), .B1(new_n921), .B2(new_n615), .ZN(G295));
  OAI21_X1  g497(.A(new_n898), .B1(new_n921), .B2(new_n615), .ZN(G331));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n534), .A2(new_n535), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n537), .A2(new_n538), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(G651), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n568), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  NOR3_X1   g503(.A1(new_n536), .A2(new_n539), .A3(KEYINPUT73), .ZN(new_n929));
  OAI21_X1  g504(.A(G168), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(G286), .B1(new_n539), .B2(new_n536), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n932), .A2(new_n856), .A3(new_n861), .A4(new_n858), .ZN(new_n933));
  AOI21_X1  g508(.A(G171), .B1(new_n574), .B2(new_n573), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n934), .B1(new_n571), .B2(G168), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n862), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n916), .A2(new_n937), .A3(new_n918), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n914), .A2(new_n933), .A3(new_n936), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n905), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(new_n903), .ZN(new_n942));
  AOI21_X1  g517(.A(G37), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT110), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n939), .A2(new_n944), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n914), .A2(new_n933), .A3(new_n936), .A4(KEYINPUT110), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n906), .A2(new_n938), .A3(new_n945), .A4(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n943), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n924), .B1(new_n948), .B2(KEYINPUT43), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n938), .A2(new_n945), .A3(new_n946), .ZN(new_n950));
  AOI21_X1  g525(.A(G37), .B1(new_n950), .B2(new_n942), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT111), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n947), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AOI211_X1 g528(.A(KEYINPUT111), .B(G37), .C1(new_n950), .C2(new_n942), .ZN(new_n954));
  OR2_X1    g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n949), .B1(new_n955), .B2(KEYINPUT43), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT43), .B1(new_n953), .B2(new_n954), .ZN(new_n957));
  OR2_X1    g532(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT112), .B1(new_n959), .B2(new_n924), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT112), .ZN(new_n961));
  AOI211_X1 g536(.A(new_n961), .B(KEYINPUT44), .C1(new_n957), .C2(new_n958), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n956), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT113), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI211_X1 g540(.A(KEYINPUT113), .B(new_n956), .C1(new_n960), .C2(new_n962), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(G397));
  INV_X1    g542(.A(G1996), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n727), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n817), .B(G2067), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n970), .B1(G1996), .B2(new_n726), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n795), .A2(new_n797), .ZN(new_n973));
  OAI22_X1  g548(.A1(new_n972), .A2(new_n973), .B1(G2067), .B2(new_n817), .ZN(new_n974));
  INV_X1    g549(.A(G1384), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n880), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT45), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n470), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n979), .B1(new_n490), .B2(G125), .ZN(new_n980));
  OAI21_X1  g555(.A(KEYINPUT67), .B1(new_n980), .B2(new_n460), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n471), .A2(new_n472), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n981), .A2(new_n982), .A3(G40), .A4(new_n466), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n978), .A2(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n794), .B(new_n797), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n985), .B(KEYINPUT114), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n969), .A2(new_n971), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n984), .ZN(new_n988));
  NOR2_X1   g563(.A1(G290), .A2(G1986), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n984), .A2(new_n989), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n990), .B(KEYINPUT48), .ZN(new_n991));
  AOI22_X1  g566(.A1(new_n974), .A2(new_n984), .B1(new_n988), .B2(new_n991), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n978), .A2(new_n983), .A3(G1996), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n993), .A2(KEYINPUT46), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(KEYINPUT46), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n984), .B1(new_n970), .B2(new_n726), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n997), .B(KEYINPUT47), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n992), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT127), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n576), .A2(G8), .A3(new_n577), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n1001), .B(KEYINPUT55), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1003), .B1(new_n503), .B2(new_n975), .ZN(new_n1004));
  AND3_X1   g579(.A1(new_n880), .A2(new_n1003), .A3(new_n975), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n1004), .A2(new_n983), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n807), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n977), .A2(G1384), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n983), .B1(new_n880), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n503), .A2(new_n975), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n977), .ZN(new_n1012));
  AOI21_X1  g587(.A(G1971), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(G8), .B1(new_n1008), .B2(new_n1013), .ZN(new_n1014));
  OR2_X1    g589(.A1(new_n1002), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n983), .A2(new_n976), .ZN(new_n1017));
  INV_X1    g592(.A(G8), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G1976), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1019), .B1(new_n1020), .B2(G288), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT52), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT116), .ZN(new_n1023));
  AND2_X1   g598(.A1(G305), .A2(G1981), .ZN(new_n1024));
  NOR2_X1   g599(.A1(G305), .A2(G1981), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1023), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n1026), .A2(KEYINPUT49), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1019), .B1(new_n1026), .B2(KEYINPUT49), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1022), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT52), .B1(G288), .B2(new_n1020), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT115), .B1(new_n1021), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1021), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT115), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1033), .A2(new_n1034), .A3(new_n1030), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1029), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1016), .A2(new_n1036), .ZN(new_n1037));
  OR2_X1    g612(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1038));
  NOR2_X1   g613(.A1(G288), .A2(G1976), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1025), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1019), .ZN(new_n1041));
  OR2_X1    g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1037), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT63), .ZN(new_n1044));
  INV_X1    g619(.A(G40), .ZN(new_n1045));
  NOR3_X1   g620(.A1(new_n473), .A2(new_n1045), .A3(new_n474), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n976), .A2(KEYINPUT50), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1046), .B(new_n1047), .C1(new_n1011), .C2(KEYINPUT50), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1048), .A2(G2090), .ZN(new_n1049));
  OAI21_X1  g624(.A(G8), .B1(new_n1049), .B2(new_n1013), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1002), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1002), .A2(KEYINPUT117), .A3(new_n1050), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1053), .A2(new_n1015), .A3(new_n1054), .A4(new_n1036), .ZN(new_n1055));
  INV_X1    g630(.A(G1966), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1009), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n496), .A2(new_n498), .A3(G2104), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n492), .B1(new_n462), .B2(new_n463), .ZN(new_n1059));
  OAI21_X1  g634(.A(KEYINPUT69), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n494), .A2(new_n499), .A3(new_n500), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n489), .A2(new_n491), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1057), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n978), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n501), .A2(new_n502), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n489), .A2(new_n491), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1065), .B(new_n1009), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(new_n1046), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1056), .B1(new_n1066), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1004), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1005), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1072), .A2(new_n739), .A3(new_n1046), .A4(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1018), .B1(new_n1071), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(G168), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1044), .B1(new_n1055), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1002), .A2(new_n1014), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1076), .A2(new_n1044), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1015), .A2(new_n1036), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1043), .B1(new_n1077), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1082), .B1(new_n1083), .B2(G2078), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT45), .B1(new_n880), .B2(new_n975), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n503), .A2(new_n1009), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1085), .B1(new_n1086), .B2(KEYINPUT118), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n983), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1088));
  INV_X1    g663(.A(G2078), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1087), .A2(new_n1088), .A3(KEYINPUT53), .A4(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1072), .A2(new_n1046), .A3(new_n1073), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n715), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1084), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n571), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT124), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1093), .A2(KEYINPUT124), .A3(new_n571), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT123), .ZN(new_n1100));
  NAND2_X1  g675(.A1(G286), .A2(G8), .ZN(new_n1101));
  XNOR2_X1  g676(.A(new_n1101), .B(KEYINPUT121), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(KEYINPUT122), .B1(new_n1075), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(G1966), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1105));
  NOR4_X1   g680(.A1(new_n1004), .A2(new_n1005), .A3(new_n983), .A4(G2084), .ZN(new_n1106));
  OAI21_X1  g681(.A(G8), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1107), .A2(new_n1108), .A3(new_n1102), .ZN(new_n1109));
  AND3_X1   g684(.A1(new_n1104), .A2(KEYINPUT51), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1102), .B1(new_n1071), .B2(new_n1074), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1112), .B1(new_n1104), .B2(KEYINPUT51), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1100), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1108), .B1(new_n1107), .B2(new_n1102), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT51), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1111), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1104), .A2(new_n1109), .A3(KEYINPUT51), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1117), .A2(KEYINPUT123), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1114), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1099), .B1(new_n1120), .B2(KEYINPUT62), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT62), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1114), .A2(new_n1122), .A3(new_n1119), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n466), .A2(G40), .ZN(new_n1124));
  NOR3_X1   g699(.A1(new_n1085), .A2(new_n471), .A3(new_n1124), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1125), .A2(KEYINPUT125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1125), .A2(KEYINPUT125), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n880), .A2(new_n1009), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1129), .A2(KEYINPUT53), .A3(new_n1089), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1092), .B(new_n1084), .C1(new_n1128), .C2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(G171), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT126), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1133), .B1(new_n1093), .B2(new_n571), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  NOR3_X1   g710(.A1(new_n1093), .A2(new_n1133), .A3(new_n571), .ZN(new_n1136));
  OAI21_X1  g711(.A(KEYINPUT54), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT54), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1138), .B1(new_n1131), .B2(new_n571), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1137), .B1(new_n1098), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(KEYINPUT57), .B1(G299), .B2(KEYINPUT119), .ZN(new_n1141));
  OAI211_X1 g716(.A(KEYINPUT119), .B(KEYINPUT57), .C1(new_n618), .C2(new_n619), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1048), .A2(new_n828), .ZN(new_n1145));
  XNOR2_X1  g720(.A(KEYINPUT56), .B(G2072), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1010), .A2(new_n1012), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1144), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(G1348), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1091), .A2(new_n1149), .ZN(new_n1150));
  OR2_X1    g725(.A1(new_n983), .A2(new_n976), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1151), .A2(G2067), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n611), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1144), .A2(new_n1145), .A3(new_n1147), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1148), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT60), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1150), .A2(new_n1153), .A3(new_n1157), .A4(new_n834), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT59), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1010), .A2(new_n1012), .A3(new_n968), .ZN(new_n1160));
  XOR2_X1   g735(.A(KEYINPUT58), .B(G1341), .Z(new_n1161));
  NAND2_X1  g736(.A1(new_n1151), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1159), .B1(new_n1163), .B2(new_n547), .ZN(new_n1164));
  AOI211_X1 g739(.A(KEYINPUT59), .B(new_n855), .C1(new_n1160), .C2(new_n1162), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1158), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1006), .A2(G1348), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n834), .B1(new_n1167), .B2(new_n1152), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1150), .A2(new_n611), .A3(new_n1153), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1157), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1156), .B1(new_n1166), .B2(new_n1170), .ZN(new_n1171));
  OR2_X1    g746(.A1(new_n1155), .A2(KEYINPUT61), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT61), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(KEYINPUT120), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1156), .A2(new_n1155), .A3(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1171), .A2(new_n1172), .A3(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1176), .B1(new_n1114), .B2(new_n1119), .ZN(new_n1177));
  AOI22_X1  g752(.A1(new_n1121), .A2(new_n1123), .B1(new_n1140), .B2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1081), .B1(new_n1178), .B2(new_n1055), .ZN(new_n1179));
  XNOR2_X1  g754(.A(G290), .B(G1986), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n984), .B1(new_n987), .B2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1000), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1182));
  AND3_X1   g757(.A1(new_n1117), .A2(KEYINPUT123), .A3(new_n1118), .ZN(new_n1183));
  AOI21_X1  g758(.A(KEYINPUT123), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1184));
  OAI21_X1  g759(.A(KEYINPUT62), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1185), .A2(new_n1123), .A3(new_n1098), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1176), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1140), .A2(new_n1120), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1055), .B1(new_n1186), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(new_n1081), .ZN(new_n1190));
  OAI211_X1 g765(.A(new_n1000), .B(new_n1181), .C1(new_n1189), .C2(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n999), .B1(new_n1182), .B2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g768(.A1(G229), .A2(new_n458), .A3(G401), .A4(G227), .ZN(new_n1195));
  NAND3_X1  g769(.A1(new_n1195), .A2(new_n896), .A3(new_n959), .ZN(G225));
  INV_X1    g770(.A(G225), .ZN(G308));
endmodule


