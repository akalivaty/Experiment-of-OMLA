//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1 0 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 1 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993;
  INV_X1    g000(.A(G224), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G953), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT83), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT7), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT84), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT66), .B1(new_n193), .B2(G143), .ZN(new_n194));
  AND2_X1   g008(.A1(KEYINPUT64), .A2(G146), .ZN(new_n195));
  NOR2_X1   g009(.A1(KEYINPUT64), .A2(G146), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n194), .B1(new_n197), .B2(G143), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(new_n193), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT66), .ZN(new_n201));
  NAND2_X1  g015(.A1(KEYINPUT64), .A2(G146), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n200), .A2(new_n201), .A3(G143), .A4(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  OAI211_X1 g018(.A(KEYINPUT0), .B(G128), .C1(new_n198), .C2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT0), .B(G128), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n208), .B1(new_n195), .B2(new_n196), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(G146), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  AOI211_X1 g025(.A(new_n206), .B(new_n207), .C1(new_n209), .C2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n209), .A2(new_n211), .ZN(new_n213));
  INV_X1    g027(.A(new_n207), .ZN(new_n214));
  AOI21_X1  g028(.A(KEYINPUT65), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n205), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G125), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT1), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n218), .B(G128), .C1(new_n198), .C2(new_n204), .ZN(new_n219));
  INV_X1    g033(.A(G125), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n218), .B1(new_n197), .B2(G143), .ZN(new_n221));
  INV_X1    g035(.A(G128), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n213), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n219), .A2(new_n220), .A3(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n192), .B1(new_n217), .B2(new_n224), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n219), .A2(new_n220), .A3(new_n223), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n226), .A2(KEYINPUT84), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n191), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n191), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT64), .B(G146), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n210), .B1(new_n230), .B2(new_n208), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n206), .B1(new_n231), .B2(new_n207), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n213), .A2(KEYINPUT65), .A3(new_n214), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n200), .A2(G143), .A3(new_n202), .ZN(new_n234));
  INV_X1    g048(.A(new_n194), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n222), .B1(new_n236), .B2(new_n203), .ZN(new_n237));
  AOI22_X1  g051(.A1(new_n232), .A2(new_n233), .B1(new_n237), .B2(KEYINPUT0), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n224), .B(new_n229), .C1(new_n238), .C2(new_n220), .ZN(new_n239));
  INV_X1    g053(.A(G104), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n240), .A2(G107), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT78), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n242), .A2(KEYINPUT3), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT3), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n244), .A2(KEYINPUT78), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n241), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G101), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n240), .A2(G107), .ZN(new_n248));
  INV_X1    g062(.A(G107), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G104), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n244), .A2(KEYINPUT78), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n246), .A2(new_n247), .A3(new_n248), .A4(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n250), .A2(new_n248), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G101), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G119), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G116), .ZN(new_n258));
  INV_X1    g072(.A(G116), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G119), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n258), .A2(new_n260), .A3(KEYINPUT69), .ZN(new_n261));
  AOI21_X1  g075(.A(KEYINPUT69), .B1(new_n258), .B2(new_n260), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT5), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(new_n257), .A3(G116), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n265), .A2(G113), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n258), .A2(new_n260), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT2), .B(G113), .ZN(new_n269));
  OR2_X1    g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n256), .A2(new_n267), .A3(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(G110), .B(G122), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n272), .B(KEYINPUT8), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n266), .B1(new_n264), .B2(new_n268), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n274), .A2(new_n270), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n271), .B(new_n273), .C1(new_n256), .C2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n252), .A2(new_n248), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n242), .A2(KEYINPUT3), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n250), .B1(new_n251), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(G101), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n280), .A2(new_n253), .A3(KEYINPUT4), .ZN(new_n281));
  INV_X1    g095(.A(new_n262), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n258), .A2(new_n260), .A3(KEYINPUT69), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(new_n283), .A3(new_n269), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n270), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT4), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n286), .B(G101), .C1(new_n277), .C2(new_n279), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n281), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n267), .A2(new_n253), .A3(new_n255), .A4(new_n270), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(new_n272), .A3(new_n289), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n239), .A2(new_n276), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(G902), .B1(new_n228), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n232), .A2(new_n233), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n220), .B1(new_n293), .B2(new_n205), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT82), .B1(new_n294), .B2(new_n226), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT82), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n296), .B(new_n224), .C1(new_n238), .C2(new_n220), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n295), .A2(new_n190), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n190), .B1(new_n295), .B2(new_n297), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n288), .A2(new_n289), .ZN(new_n301));
  INV_X1    g115(.A(new_n272), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n303), .A2(KEYINPUT81), .A3(KEYINPUT6), .A4(new_n290), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT81), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT6), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n301), .B(new_n302), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n292), .B1(new_n300), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(G210), .B1(G237), .B2(G902), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT85), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n292), .B(new_n310), .C1(new_n300), .C2(new_n308), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  OR2_X1    g129(.A1(new_n314), .A2(new_n313), .ZN(new_n316));
  AND2_X1   g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT9), .B(G234), .ZN(new_n318));
  OAI21_X1  g132(.A(G221), .B1(new_n318), .B2(G902), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G469), .ZN(new_n321));
  INV_X1    g135(.A(G902), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G134), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G137), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT11), .ZN(new_n326));
  INV_X1    g140(.A(G137), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n326), .B1(G134), .B2(new_n327), .ZN(new_n328));
  NOR3_X1   g142(.A1(new_n324), .A2(KEYINPUT11), .A3(G137), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n325), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G131), .ZN(new_n331));
  INV_X1    g145(.A(G131), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n332), .B(new_n325), .C1(new_n328), .C2(new_n329), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n219), .A2(new_n223), .ZN(new_n335));
  INV_X1    g149(.A(new_n256), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(G128), .B1(new_n210), .B2(new_n218), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n236), .A2(new_n203), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n256), .B1(new_n339), .B2(new_n219), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n334), .B1(new_n337), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT12), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI211_X1 g157(.A(KEYINPUT12), .B(new_n334), .C1(new_n337), .C2(new_n340), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT79), .B(KEYINPUT10), .ZN(new_n346));
  OR2_X1    g160(.A1(new_n340), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n334), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n293), .A2(new_n281), .A3(new_n205), .A4(new_n287), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n335), .A2(KEYINPUT10), .A3(new_n336), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n347), .A2(new_n348), .A3(new_n349), .A4(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n345), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(G110), .B(G140), .ZN(new_n353));
  INV_X1    g167(.A(G227), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n354), .A2(G953), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n353), .B(new_n355), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n350), .B(new_n349), .C1(new_n340), .C2(new_n346), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n357), .A2(new_n334), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n358), .A2(new_n356), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n334), .ZN(new_n360));
  AOI22_X1  g174(.A1(new_n352), .A2(new_n356), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n323), .B1(new_n361), .B2(G469), .ZN(new_n362));
  INV_X1    g176(.A(new_n356), .ZN(new_n363));
  OAI211_X1 g177(.A(KEYINPUT80), .B(new_n363), .C1(new_n357), .C2(new_n334), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n345), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(KEYINPUT80), .B1(new_n351), .B2(new_n363), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n351), .A2(new_n360), .ZN(new_n367));
  OAI22_X1  g181(.A1(new_n365), .A2(new_n366), .B1(new_n367), .B2(new_n363), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(new_n321), .A3(new_n322), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n320), .B1(new_n362), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G952), .ZN(new_n371));
  AOI211_X1 g185(.A(G953), .B(new_n371), .C1(G234), .C2(G237), .ZN(new_n372));
  NAND2_X1  g186(.A1(G234), .A2(G237), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(G902), .A3(G953), .ZN(new_n374));
  XOR2_X1   g188(.A(new_n374), .B(KEYINPUT92), .Z(new_n375));
  XNOR2_X1  g189(.A(KEYINPUT21), .B(G898), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n372), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(G214), .B1(G237), .B2(G902), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n317), .A2(new_n370), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT17), .ZN(new_n382));
  INV_X1    g196(.A(G237), .ZN(new_n383));
  INV_X1    g197(.A(G953), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(G214), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT86), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G143), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(KEYINPUT86), .B(G143), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n388), .B1(new_n389), .B2(new_n385), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n332), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT88), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n390), .A2(new_n393), .A3(G131), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n393), .B1(new_n390), .B2(G131), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n382), .B(new_n392), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n390), .A2(G131), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(KEYINPUT88), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n390), .A2(new_n393), .A3(G131), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n398), .A2(KEYINPUT17), .A3(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT89), .ZN(new_n401));
  INV_X1    g215(.A(G140), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G125), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n220), .A2(G140), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n403), .A2(new_n404), .A3(KEYINPUT75), .ZN(new_n405));
  OR3_X1    g219(.A1(new_n402), .A2(KEYINPUT75), .A3(G125), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT16), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT16), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n403), .A2(new_n408), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n407), .A2(new_n193), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n193), .B1(new_n407), .B2(new_n409), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n401), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n407), .A2(new_n409), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G146), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n407), .A2(new_n193), .A3(new_n409), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(KEYINPUT89), .A3(new_n415), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n396), .A2(new_n400), .A3(new_n412), .A4(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(G113), .B(G122), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(new_n240), .ZN(new_n419));
  NAND2_X1  g233(.A1(KEYINPUT87), .A2(KEYINPUT18), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n391), .B1(new_n332), .B2(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(G125), .B(G140), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n197), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n405), .A2(new_n406), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n423), .B1(new_n424), .B2(new_n193), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n421), .B(new_n425), .C1(new_n420), .C2(new_n397), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n417), .A2(new_n419), .A3(new_n426), .ZN(new_n427));
  AOI22_X1  g241(.A1(new_n398), .A2(new_n399), .B1(new_n332), .B2(new_n391), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n422), .A2(KEYINPUT19), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n429), .B1(new_n424), .B2(KEYINPUT19), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n414), .B1(new_n230), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n426), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n419), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n427), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g249(.A1(G475), .A2(G902), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(KEYINPUT90), .B1(new_n427), .B2(new_n434), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n437), .B1(KEYINPUT20), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT20), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n435), .A2(KEYINPUT90), .A3(new_n440), .A4(new_n436), .ZN(new_n441));
  INV_X1    g255(.A(new_n427), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n419), .B1(new_n417), .B2(new_n426), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n322), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n439), .A2(new_n441), .B1(G475), .B2(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(G116), .B(G122), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(G107), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(new_n249), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT91), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(KEYINPUT13), .B1(new_n222), .B2(G143), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n453), .A2(new_n324), .ZN(new_n454));
  XNOR2_X1  g268(.A(G128), .B(G143), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n448), .A2(KEYINPUT91), .A3(new_n449), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n452), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n259), .A2(KEYINPUT14), .A3(G122), .ZN(new_n459));
  OAI211_X1 g273(.A(G107), .B(new_n459), .C1(new_n447), .C2(KEYINPUT14), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n455), .A2(G134), .ZN(new_n461));
  OR2_X1    g275(.A1(new_n455), .A2(G134), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n460), .A2(new_n449), .A3(new_n461), .A4(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(G217), .ZN(new_n465));
  NOR3_X1   g279(.A1(new_n318), .A2(new_n465), .A3(G953), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n458), .A2(new_n463), .A3(new_n466), .ZN(new_n469));
  AOI21_X1  g283(.A(G902), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G478), .ZN(new_n471));
  OR2_X1    g285(.A1(new_n471), .A2(KEYINPUT15), .ZN(new_n472));
  XOR2_X1   g286(.A(new_n470), .B(new_n472), .Z(new_n473));
  NAND2_X1  g287(.A1(new_n445), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n381), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT32), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT67), .B1(new_n327), .B2(G134), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n327), .A2(G134), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n325), .A2(KEYINPUT67), .ZN(new_n480));
  OAI21_X1  g294(.A(G131), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AND2_X1   g295(.A1(new_n481), .A2(new_n333), .ZN(new_n482));
  AOI211_X1 g296(.A(KEYINPUT1), .B(new_n222), .C1(new_n236), .C2(new_n203), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n234), .A2(KEYINPUT1), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n231), .B1(G128), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n482), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n334), .B(new_n205), .C1(new_n215), .C2(new_n212), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n486), .A2(new_n487), .A3(KEYINPUT30), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT70), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT70), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n486), .A2(new_n487), .A3(new_n490), .A4(KEYINPUT30), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT68), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n486), .A2(new_n487), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT30), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AOI211_X1 g310(.A(KEYINPUT68), .B(KEYINPUT30), .C1(new_n486), .C2(new_n487), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n492), .B(new_n285), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT31), .ZN(new_n499));
  INV_X1    g313(.A(new_n285), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n486), .A2(new_n487), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n503));
  INV_X1    g317(.A(G210), .ZN(new_n504));
  NOR3_X1   g318(.A1(new_n504), .A2(G237), .A3(G953), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n503), .B(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(KEYINPUT26), .B(G101), .ZN(new_n507));
  XOR2_X1   g321(.A(new_n506), .B(new_n507), .Z(new_n508));
  NOR2_X1   g322(.A1(new_n502), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n498), .A2(new_n499), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n502), .A2(KEYINPUT28), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT28), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n501), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n494), .A2(new_n285), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n511), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n508), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n510), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n509), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n238), .A2(new_n334), .B1(new_n335), .B2(new_n482), .ZN(new_n519));
  OAI21_X1  g333(.A(KEYINPUT68), .B1(new_n519), .B2(KEYINPUT30), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n494), .A2(new_n493), .A3(new_n495), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n520), .A2(new_n521), .B1(new_n489), .B2(new_n491), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n518), .B1(new_n522), .B2(new_n285), .ZN(new_n523));
  OAI21_X1  g337(.A(KEYINPUT72), .B1(new_n523), .B2(new_n499), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n498), .A2(new_n509), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT72), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n525), .A2(new_n526), .A3(KEYINPUT31), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n517), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(G472), .A2(G902), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n476), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT74), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n530), .A2(new_n476), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n532), .B1(new_n528), .B2(new_n534), .ZN(new_n535));
  AOI22_X1  g349(.A1(new_n523), .A2(new_n499), .B1(new_n508), .B2(new_n515), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n526), .B1(new_n525), .B2(KEYINPUT31), .ZN(new_n537));
  AOI211_X1 g351(.A(KEYINPUT72), .B(new_n499), .C1(new_n498), .C2(new_n509), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n539), .A2(KEYINPUT74), .A3(new_n533), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n501), .A2(KEYINPUT73), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT73), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n486), .A2(new_n487), .A3(new_n542), .A4(new_n500), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n541), .A2(new_n514), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT28), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n545), .A2(new_n513), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT29), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n508), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(G902), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n498), .A2(new_n508), .A3(new_n501), .ZN(new_n550));
  INV_X1    g364(.A(new_n508), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n515), .A2(new_n551), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n549), .B1(new_n553), .B2(KEYINPUT29), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(G472), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n531), .A2(new_n535), .A3(new_n540), .A4(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT77), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n465), .B1(G234), .B2(new_n322), .ZN(new_n558));
  XOR2_X1   g372(.A(KEYINPUT24), .B(G110), .Z(new_n559));
  XNOR2_X1  g373(.A(G119), .B(G128), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT23), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n562), .B1(new_n257), .B2(G128), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n222), .A2(KEYINPUT23), .A3(G119), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n563), .B(new_n564), .C1(G119), .C2(new_n222), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(G110), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n561), .B(new_n566), .C1(new_n410), .C2(new_n411), .ZN(new_n567));
  OAI22_X1  g381(.A1(new_n565), .A2(G110), .B1(new_n560), .B2(new_n559), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n414), .A2(new_n423), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n384), .A2(G221), .A3(G234), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(KEYINPUT76), .ZN(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT22), .B(G137), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n572), .B(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n567), .A2(new_n569), .A3(new_n574), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n578), .A2(KEYINPUT25), .A3(new_n322), .ZN(new_n579));
  AOI21_X1  g393(.A(KEYINPUT25), .B1(new_n578), .B2(new_n322), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n558), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n558), .A2(G902), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  AND3_X1   g398(.A1(new_n556), .A2(new_n557), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n557), .B1(new_n556), .B2(new_n584), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n475), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(G101), .ZN(G3));
  OAI21_X1  g402(.A(G472), .B1(new_n528), .B2(G902), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n539), .A2(new_n529), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n370), .ZN(new_n592));
  INV_X1    g406(.A(new_n584), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n470), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n595), .A2(KEYINPUT93), .A3(new_n471), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT93), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n597), .B1(new_n470), .B2(G478), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n468), .A2(new_n469), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(KEYINPUT33), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT33), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n468), .A2(new_n601), .A3(new_n469), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n471), .A2(G902), .ZN(new_n604));
  AOI22_X1  g418(.A1(new_n596), .A2(new_n598), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n445), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n312), .A2(new_n314), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n380), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n594), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT34), .B(G104), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G6));
  INV_X1    g427(.A(new_n473), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n444), .A2(G475), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT94), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n437), .B1(new_n616), .B2(KEYINPUT20), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(KEYINPUT95), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n616), .A2(KEYINPUT20), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT95), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n437), .B(new_n620), .C1(new_n616), .C2(KEYINPUT20), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n618), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n619), .B1(new_n618), .B2(new_n621), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n614), .B(new_n615), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n624), .A2(new_n609), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n594), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT35), .B(G107), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G9));
  NOR2_X1   g442(.A1(new_n574), .A2(KEYINPUT36), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n570), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n582), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n581), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n381), .A2(new_n474), .A3(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n591), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT37), .B(G110), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G12));
  NAND2_X1  g452(.A1(new_n608), .A2(new_n378), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n592), .A2(new_n633), .A3(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(G900), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n375), .A2(new_n641), .ZN(new_n642));
  AND2_X1   g456(.A1(new_n642), .A2(KEYINPUT96), .ZN(new_n643));
  INV_X1    g457(.A(new_n372), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n644), .B1(new_n642), .B2(KEYINPUT96), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n624), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n556), .A2(new_n640), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G128), .ZN(G30));
  XOR2_X1   g463(.A(new_n317), .B(KEYINPUT38), .Z(new_n650));
  XOR2_X1   g464(.A(new_n646), .B(KEYINPUT39), .Z(new_n651));
  NAND2_X1  g465(.A1(new_n370), .A2(new_n651), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n652), .A2(KEYINPUT40), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n633), .A2(new_n378), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n650), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n445), .A2(new_n473), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n535), .A2(new_n540), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n508), .B1(new_n498), .B2(new_n501), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n322), .B1(new_n544), .B2(new_n551), .ZN(new_n659));
  OAI21_X1  g473(.A(G472), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n531), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  OR2_X1    g476(.A1(new_n652), .A2(KEYINPUT40), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n655), .A2(new_n656), .A3(new_n662), .A4(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G143), .ZN(G45));
  NOR2_X1   g479(.A1(new_n607), .A2(new_n646), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n556), .A2(new_n640), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(KEYINPUT97), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT97), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n556), .A2(new_n640), .A3(new_n669), .A4(new_n666), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G146), .ZN(G48));
  NAND2_X1  g486(.A1(new_n368), .A2(new_n322), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(G469), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n674), .A2(new_n319), .A3(new_n369), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n675), .A2(new_n593), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n556), .A2(new_n610), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(KEYINPUT41), .B(G113), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G15));
  NAND3_X1  g493(.A1(new_n556), .A2(new_n625), .A3(new_n676), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G116), .ZN(G18));
  INV_X1    g495(.A(new_n377), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n632), .A2(new_n682), .ZN(new_n683));
  NOR4_X1   g497(.A1(new_n675), .A2(new_n639), .A3(new_n474), .A4(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n556), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G119), .ZN(G21));
  AND3_X1   g500(.A1(new_n498), .A2(new_n499), .A3(new_n509), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n499), .B1(new_n498), .B2(new_n509), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n551), .B1(new_n545), .B2(new_n513), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g504(.A(KEYINPUT98), .B1(new_n690), .B2(new_n530), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT98), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n525), .A2(KEYINPUT31), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n510), .ZN(new_n694));
  OAI211_X1 g508(.A(new_n692), .B(new_n529), .C1(new_n694), .C2(new_n689), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n674), .A2(new_n319), .A3(new_n369), .A4(new_n682), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n439), .A2(new_n441), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n615), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n608), .A2(new_n700), .A3(new_n614), .A4(new_n378), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n697), .A2(new_n702), .A3(new_n584), .A4(new_n589), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G122), .ZN(G24));
  INV_X1    g518(.A(G472), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n705), .B1(new_n539), .B2(new_n322), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n696), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n675), .A2(new_n639), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n707), .A2(new_n632), .A3(new_n666), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G125), .ZN(G27));
  AOI21_X1  g524(.A(new_n379), .B1(new_n315), .B2(new_n316), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT42), .ZN(new_n712));
  NOR4_X1   g526(.A1(new_n445), .A2(new_n712), .A3(new_n605), .A4(new_n646), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n711), .A2(new_n713), .A3(new_n370), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n539), .A2(new_n533), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n531), .A2(new_n555), .A3(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n714), .A2(new_n716), .A3(new_n584), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(KEYINPUT99), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT99), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n714), .A2(new_n716), .A3(new_n719), .A4(new_n584), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n711), .A2(new_n370), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n556), .A2(new_n584), .A3(new_n666), .A4(new_n721), .ZN(new_n722));
  AOI22_X1  g536(.A1(new_n718), .A2(new_n720), .B1(new_n722), .B2(new_n712), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n332), .ZN(G33));
  NAND4_X1  g538(.A1(new_n556), .A2(new_n647), .A3(new_n584), .A4(new_n721), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G134), .ZN(G36));
  XOR2_X1   g540(.A(new_n711), .B(KEYINPUT101), .Z(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n605), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n445), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(KEYINPUT43), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n635), .A2(new_n633), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n728), .B1(KEYINPUT44), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n361), .A2(KEYINPUT45), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT100), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n361), .A2(KEYINPUT45), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(new_n321), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n323), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n369), .B1(new_n739), .B2(KEYINPUT46), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT46), .ZN(new_n741));
  AOI211_X1 g555(.A(new_n741), .B(new_n323), .C1(new_n736), .C2(new_n738), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n319), .B(new_n651), .C1(new_n740), .C2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n733), .B(new_n744), .C1(KEYINPUT44), .C2(new_n732), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G137), .ZN(G39));
  OAI21_X1  g560(.A(new_n319), .B1(new_n740), .B2(new_n742), .ZN(new_n747));
  XOR2_X1   g561(.A(KEYINPUT102), .B(KEYINPUT47), .Z(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT47), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n750), .A2(KEYINPUT102), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n749), .B1(new_n747), .B2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n666), .ZN(new_n753));
  INV_X1    g567(.A(new_n711), .ZN(new_n754));
  NOR4_X1   g568(.A1(new_n556), .A2(new_n753), .A3(new_n584), .A4(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(KEYINPUT103), .ZN(new_n756));
  OR2_X1    g570(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G140), .ZN(G42));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n709), .A2(new_n648), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n760), .B1(new_n670), .B2(new_n668), .ZN(new_n761));
  INV_X1    g575(.A(new_n646), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n370), .A2(new_n633), .A3(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT107), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n763), .B(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n639), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n765), .A2(new_n662), .A3(new_n766), .A4(new_n656), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n759), .B1(new_n761), .B2(new_n767), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n709), .A2(new_n648), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n671), .A2(new_n769), .A3(new_n767), .A4(new_n759), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n591), .A2(new_n593), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n474), .B1(new_n445), .B2(new_n729), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n381), .A2(new_n774), .ZN(new_n775));
  AOI22_X1  g589(.A1(new_n634), .A2(new_n635), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n633), .A2(new_n614), .A3(new_n646), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n777), .B(new_n615), .C1(new_n622), .C2(new_n623), .ZN(new_n778));
  AOI22_X1  g592(.A1(new_n590), .A2(new_n476), .B1(G472), .B2(new_n554), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n778), .B1(new_n657), .B2(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n589), .A2(new_n632), .A3(new_n691), .A4(new_n695), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n781), .A2(new_n753), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n721), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n587), .A2(new_n725), .A3(new_n776), .A4(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT108), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n725), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n622), .A2(new_n623), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n556), .A2(new_n615), .A3(new_n788), .A4(new_n777), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n707), .A2(new_n632), .A3(new_n666), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n787), .B1(new_n791), .B2(new_n721), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n792), .A2(KEYINPUT108), .A3(new_n587), .A4(new_n776), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n786), .A2(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n680), .A2(new_n677), .A3(new_n685), .A4(new_n703), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT109), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n760), .A2(KEYINPUT52), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n718), .A2(new_n720), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n722), .A2(new_n712), .ZN(new_n799));
  OAI211_X1 g613(.A(KEYINPUT53), .B(new_n797), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n772), .A2(new_n794), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n671), .A2(new_n769), .A3(new_n767), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(KEYINPUT52), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT106), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n795), .A2(new_n805), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n696), .A2(new_n706), .A3(new_n593), .ZN(new_n807));
  AOI22_X1  g621(.A1(new_n807), .A2(new_n702), .B1(new_n556), .B2(new_n684), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n808), .A2(KEYINPUT106), .A3(new_n677), .A4(new_n680), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n723), .B1(new_n806), .B2(new_n809), .ZN(new_n810));
  AND4_X1   g624(.A1(new_n587), .A2(new_n725), .A3(new_n776), .A4(new_n783), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n804), .A2(new_n810), .A3(new_n811), .A4(new_n770), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n802), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n810), .A2(new_n811), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n797), .A2(new_n813), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n772), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n815), .B1(new_n819), .B2(new_n814), .ZN(new_n820));
  OAI21_X1  g634(.A(KEYINPUT110), .B1(new_n816), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT53), .B1(new_n772), .B2(new_n817), .ZN(new_n822));
  INV_X1    g636(.A(new_n818), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n812), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(KEYINPUT54), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT110), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n802), .A2(new_n814), .A3(new_n815), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(KEYINPUT111), .B(KEYINPUT51), .ZN(new_n829));
  INV_X1    g643(.A(new_n675), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n650), .A2(new_n379), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n731), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n807), .A2(new_n372), .A3(new_n832), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT114), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT50), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n835), .B(KEYINPUT50), .C1(new_n831), .C2(new_n833), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT50), .B1(new_n834), .B2(new_n835), .ZN(new_n842));
  INV_X1    g656(.A(new_n840), .ZN(new_n843));
  OAI21_X1  g657(.A(KEYINPUT115), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n728), .A2(new_n833), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n674), .A2(new_n369), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n319), .B1(new_n848), .B2(KEYINPUT112), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n849), .B1(KEYINPUT112), .B2(new_n848), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(KEYINPUT113), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n847), .B1(new_n752), .B2(new_n851), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n754), .A2(KEYINPUT116), .A3(new_n675), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT116), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n854), .B1(new_n830), .B2(new_n711), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n853), .A2(new_n855), .A3(new_n644), .ZN(new_n856));
  INV_X1    g670(.A(new_n662), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n856), .A2(new_n584), .A3(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT117), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n700), .A2(new_n729), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n856), .A2(new_n832), .ZN(new_n862));
  OR2_X1    g676(.A1(new_n862), .A2(new_n781), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n859), .B1(new_n858), .B2(new_n860), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n852), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n829), .B1(new_n845), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n858), .A2(new_n606), .ZN(new_n868));
  INV_X1    g682(.A(new_n833), .ZN(new_n869));
  AOI211_X1 g683(.A(new_n371), .B(G953), .C1(new_n869), .C2(new_n708), .ZN(new_n870));
  NOR2_X1   g684(.A1(KEYINPUT118), .A2(KEYINPUT48), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n593), .B1(new_n779), .B2(new_n715), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n871), .B1(new_n862), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n868), .A2(new_n870), .A3(new_n874), .ZN(new_n875));
  AND2_X1   g689(.A1(KEYINPUT118), .A2(KEYINPUT48), .ZN(new_n876));
  NOR4_X1   g690(.A1(new_n862), .A2(new_n873), .A3(new_n871), .A4(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n752), .A2(new_n850), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n846), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n880), .A2(KEYINPUT51), .A3(new_n840), .A4(new_n838), .ZN(new_n881));
  OR2_X1    g695(.A1(new_n864), .A2(new_n865), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n878), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n867), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n821), .A2(new_n828), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n371), .A2(new_n384), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n848), .A2(KEYINPUT49), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT104), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n584), .A2(new_n319), .A3(new_n378), .ZN(new_n890));
  AOI211_X1 g704(.A(new_n730), .B(new_n890), .C1(new_n848), .C2(KEYINPUT49), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n857), .A2(new_n650), .A3(new_n889), .A4(new_n891), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT105), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n887), .A2(new_n893), .ZN(G75));
  INV_X1    g708(.A(KEYINPUT56), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n300), .B(new_n308), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT55), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n802), .A2(new_n814), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(G902), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n895), .B(new_n898), .C1(new_n900), .C2(new_n504), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n384), .A2(G952), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(KEYINPUT120), .Z(new_n903));
  NAND2_X1  g717(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n322), .B1(new_n802), .B2(new_n814), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT56), .B1(new_n905), .B2(G210), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n907), .A2(KEYINPUT119), .A3(new_n897), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT119), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n909), .B1(new_n906), .B2(new_n898), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n904), .B1(new_n908), .B2(new_n910), .ZN(G51));
  XNOR2_X1  g725(.A(new_n368), .B(KEYINPUT121), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n815), .B1(new_n802), .B2(new_n814), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n816), .A2(new_n913), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n323), .B(KEYINPUT57), .Z(new_n915));
  OAI21_X1  g729(.A(new_n912), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n905), .A2(new_n736), .A3(new_n738), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n902), .B1(new_n916), .B2(new_n917), .ZN(G54));
  AND3_X1   g732(.A1(new_n905), .A2(KEYINPUT58), .A3(G475), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n919), .A2(new_n435), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n919), .A2(new_n435), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n920), .A2(new_n921), .A3(new_n902), .ZN(G60));
  NAND2_X1  g736(.A1(G478), .A2(G902), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT59), .Z(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n603), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n903), .B1(new_n914), .B2(new_n926), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n816), .A2(new_n820), .A3(KEYINPUT110), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n826), .B1(new_n825), .B2(new_n827), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n925), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n603), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n927), .B1(new_n930), .B2(new_n931), .ZN(G63));
  NAND2_X1  g746(.A1(G217), .A2(G902), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT60), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n934), .B1(new_n802), .B2(new_n814), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n630), .B(KEYINPUT123), .Z(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(KEYINPUT61), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n903), .B1(new_n935), .B2(new_n578), .ZN(new_n939));
  OR2_X1    g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT124), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n935), .A2(new_n941), .A3(new_n936), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n941), .B1(new_n935), .B2(new_n936), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n942), .A2(new_n939), .A3(new_n943), .ZN(new_n944));
  XOR2_X1   g758(.A(KEYINPUT122), .B(KEYINPUT61), .Z(new_n945));
  OAI21_X1  g759(.A(new_n940), .B1(new_n944), .B2(new_n945), .ZN(G66));
  OAI21_X1  g760(.A(G953), .B1(new_n376), .B2(new_n187), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n806), .A2(new_n809), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n587), .A2(new_n776), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n947), .B1(new_n951), .B2(G953), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n308), .B1(G898), .B2(new_n384), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(G69));
  INV_X1    g768(.A(KEYINPUT125), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n671), .A2(new_n769), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n955), .B1(new_n671), .B2(new_n769), .ZN(new_n957));
  OR2_X1    g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n743), .A2(new_n701), .A3(new_n873), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n959), .A2(new_n723), .A3(new_n787), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n958), .A2(new_n757), .A3(new_n960), .A4(new_n745), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n384), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n522), .B(new_n430), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n963), .B1(new_n354), .B2(G953), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n641), .B1(new_n963), .B2(new_n354), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n754), .A2(new_n652), .A3(new_n774), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(new_n585), .B2(new_n586), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n745), .B(new_n968), .C1(new_n756), .C2(new_n752), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n664), .B1(new_n956), .B2(new_n957), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n969), .B1(KEYINPUT62), .B2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT62), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n972), .B(new_n664), .C1(new_n956), .C2(new_n957), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n973), .A2(KEYINPUT126), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n973), .A2(KEYINPUT126), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n971), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(KEYINPUT127), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT127), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n971), .B(new_n978), .C1(new_n974), .C2(new_n975), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n963), .A2(new_n384), .ZN(new_n981));
  OAI221_X1 g795(.A(new_n965), .B1(new_n384), .B2(new_n966), .C1(new_n980), .C2(new_n981), .ZN(G72));
  NAND2_X1  g796(.A1(G472), .A2(G902), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT63), .Z(new_n984));
  OAI21_X1  g798(.A(new_n984), .B1(new_n961), .B2(new_n950), .ZN(new_n985));
  INV_X1    g799(.A(new_n550), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n902), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(new_n984), .ZN(new_n988));
  NOR3_X1   g802(.A1(new_n986), .A2(new_n658), .A3(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n989), .B1(new_n822), .B2(new_n824), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n977), .A2(new_n951), .A3(new_n979), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n984), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n991), .B1(new_n993), .B2(new_n658), .ZN(G57));
endmodule


