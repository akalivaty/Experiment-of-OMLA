

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U551 ( .A1(n778), .A2(n777), .ZN(n779) );
  NOR2_X2 U552 ( .A1(n530), .A2(n529), .ZN(G164) );
  OR2_X1 U553 ( .A1(n720), .A2(n719), .ZN(n723) );
  NAND2_X1 U554 ( .A1(n699), .A2(n794), .ZN(n724) );
  NOR2_X2 U555 ( .A1(G2104), .A2(n526), .ZN(n880) );
  NOR2_X1 U556 ( .A1(n525), .A2(G2105), .ZN(n549) );
  INV_X1 U557 ( .A(G2104), .ZN(n525) );
  XNOR2_X1 U558 ( .A(n520), .B(n519), .ZN(n573) );
  XNOR2_X1 U559 ( .A(n518), .B(KEYINPUT66), .ZN(n520) );
  INV_X1 U560 ( .A(KEYINPUT17), .ZN(n518) );
  AND2_X1 U561 ( .A1(n701), .A2(n760), .ZN(n702) );
  INV_X1 U562 ( .A(KEYINPUT103), .ZN(n773) );
  NOR2_X1 U563 ( .A1(n772), .A2(KEYINPUT33), .ZN(n774) );
  XNOR2_X1 U564 ( .A(n551), .B(n550), .ZN(n553) );
  INV_X1 U565 ( .A(KEYINPUT23), .ZN(n550) );
  INV_X1 U566 ( .A(KEYINPUT91), .ZN(n521) );
  BUF_X1 U567 ( .A(n697), .Z(G160) );
  OR2_X1 U568 ( .A1(n789), .A2(n788), .ZN(n516) );
  XOR2_X1 U569 ( .A(n544), .B(n543), .Z(n517) );
  INV_X1 U570 ( .A(KEYINPUT26), .ZN(n712) );
  BUF_X1 U571 ( .A(n724), .Z(n746) );
  INV_X1 U572 ( .A(KEYINPUT31), .ZN(n710) );
  NOR2_X1 U573 ( .A1(n724), .A2(G2084), .ZN(n700) );
  AND2_X1 U574 ( .A1(n753), .A2(n752), .ZN(n755) );
  NAND2_X1 U575 ( .A1(n665), .A2(G51), .ZN(n540) );
  XNOR2_X1 U576 ( .A(n698), .B(KEYINPUT92), .ZN(n793) );
  AND2_X1 U577 ( .A1(n790), .A2(n516), .ZN(n791) );
  INV_X1 U578 ( .A(G2105), .ZN(n526) );
  INV_X1 U579 ( .A(KEYINPUT65), .ZN(n538) );
  BUF_X1 U580 ( .A(n549), .Z(n875) );
  XOR2_X1 U581 ( .A(KEYINPUT1), .B(n537), .Z(n658) );
  XNOR2_X1 U582 ( .A(n522), .B(n521), .ZN(n523) );
  NOR2_X1 U583 ( .A1(n555), .A2(n554), .ZN(n697) );
  AND2_X1 U584 ( .A1(G2105), .A2(G2104), .ZN(n879) );
  NAND2_X1 U585 ( .A1(n879), .A2(G114), .ZN(n524) );
  NOR2_X1 U586 ( .A1(G2105), .A2(G2104), .ZN(n519) );
  NAND2_X1 U587 ( .A1(n573), .A2(G138), .ZN(n522) );
  NAND2_X1 U588 ( .A1(n524), .A2(n523), .ZN(n530) );
  NAND2_X1 U589 ( .A1(G102), .A2(n875), .ZN(n528) );
  NAND2_X1 U590 ( .A1(G126), .A2(n880), .ZN(n527) );
  NAND2_X1 U591 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U592 ( .A(KEYINPUT0), .B(G543), .Z(n641) );
  INV_X1 U593 ( .A(G651), .ZN(n536) );
  NOR2_X1 U594 ( .A1(n641), .A2(n536), .ZN(n657) );
  NAND2_X1 U595 ( .A1(n657), .A2(G76), .ZN(n531) );
  XNOR2_X1 U596 ( .A(KEYINPUT78), .B(n531), .ZN(n534) );
  NOR2_X1 U597 ( .A1(G651), .A2(G543), .ZN(n661) );
  NAND2_X1 U598 ( .A1(n661), .A2(G89), .ZN(n532) );
  XNOR2_X1 U599 ( .A(KEYINPUT4), .B(n532), .ZN(n533) );
  NAND2_X1 U600 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U601 ( .A(KEYINPUT5), .B(n535), .ZN(n545) );
  XNOR2_X1 U602 ( .A(KEYINPUT80), .B(KEYINPUT6), .ZN(n544) );
  NOR2_X1 U603 ( .A1(G543), .A2(n536), .ZN(n537) );
  NAND2_X1 U604 ( .A1(n658), .A2(G63), .ZN(n542) );
  NOR2_X1 U605 ( .A1(G651), .A2(n641), .ZN(n539) );
  XNOR2_X2 U606 ( .A(n539), .B(n538), .ZN(n665) );
  XOR2_X1 U607 ( .A(KEYINPUT79), .B(n540), .Z(n541) );
  NAND2_X1 U608 ( .A1(n542), .A2(n541), .ZN(n543) );
  NAND2_X1 U609 ( .A1(n545), .A2(n517), .ZN(n546) );
  XNOR2_X1 U610 ( .A(KEYINPUT7), .B(n546), .ZN(G168) );
  NAND2_X1 U611 ( .A1(n573), .A2(G137), .ZN(n548) );
  NAND2_X1 U612 ( .A1(n880), .A2(G125), .ZN(n547) );
  NAND2_X1 U613 ( .A1(n548), .A2(n547), .ZN(n555) );
  NAND2_X1 U614 ( .A1(G101), .A2(n549), .ZN(n551) );
  NAND2_X1 U615 ( .A1(n879), .A2(G113), .ZN(n552) );
  NAND2_X1 U616 ( .A1(n553), .A2(n552), .ZN(n554) );
  NAND2_X1 U617 ( .A1(G64), .A2(n658), .ZN(n557) );
  NAND2_X1 U618 ( .A1(G52), .A2(n665), .ZN(n556) );
  NAND2_X1 U619 ( .A1(n557), .A2(n556), .ZN(n563) );
  NAND2_X1 U620 ( .A1(n661), .A2(G90), .ZN(n558) );
  XOR2_X1 U621 ( .A(KEYINPUT67), .B(n558), .Z(n560) );
  NAND2_X1 U622 ( .A1(n657), .A2(G77), .ZN(n559) );
  NAND2_X1 U623 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U624 ( .A(KEYINPUT9), .B(n561), .Z(n562) );
  NOR2_X1 U625 ( .A1(n563), .A2(n562), .ZN(G171) );
  XOR2_X1 U626 ( .A(G2443), .B(G2446), .Z(n565) );
  XNOR2_X1 U627 ( .A(G2427), .B(G2451), .ZN(n564) );
  XNOR2_X1 U628 ( .A(n565), .B(n564), .ZN(n571) );
  XOR2_X1 U629 ( .A(G2430), .B(G2454), .Z(n567) );
  XNOR2_X1 U630 ( .A(G1341), .B(G1348), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n567), .B(n566), .ZN(n569) );
  XOR2_X1 U632 ( .A(G2435), .B(G2438), .Z(n568) );
  XNOR2_X1 U633 ( .A(n569), .B(n568), .ZN(n570) );
  XOR2_X1 U634 ( .A(n571), .B(n570), .Z(n572) );
  AND2_X1 U635 ( .A1(G14), .A2(n572), .ZN(G401) );
  AND2_X1 U636 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U637 ( .A1(G111), .A2(n879), .ZN(n576) );
  BUF_X1 U638 ( .A(n573), .Z(n574) );
  NAND2_X1 U639 ( .A1(G135), .A2(n574), .ZN(n575) );
  NAND2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n579) );
  NAND2_X1 U641 ( .A1(n880), .A2(G123), .ZN(n577) );
  XOR2_X1 U642 ( .A(KEYINPUT18), .B(n577), .Z(n578) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n581) );
  NAND2_X1 U644 ( .A1(n875), .A2(G99), .ZN(n580) );
  NAND2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n998) );
  XNOR2_X1 U646 ( .A(G2096), .B(n998), .ZN(n582) );
  OR2_X1 U647 ( .A1(G2100), .A2(n582), .ZN(G156) );
  INV_X1 U648 ( .A(G57), .ZN(G237) );
  XOR2_X1 U649 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U650 ( .A1(G7), .A2(G661), .ZN(n583) );
  XNOR2_X1 U651 ( .A(n583), .B(KEYINPUT70), .ZN(n584) );
  XNOR2_X1 U652 ( .A(KEYINPUT10), .B(n584), .ZN(G223) );
  INV_X1 U653 ( .A(G223), .ZN(n840) );
  NAND2_X1 U654 ( .A1(n840), .A2(G567), .ZN(n585) );
  XOR2_X1 U655 ( .A(KEYINPUT11), .B(n585), .Z(G234) );
  XOR2_X1 U656 ( .A(KEYINPUT12), .B(KEYINPUT72), .Z(n587) );
  NAND2_X1 U657 ( .A1(G81), .A2(n661), .ZN(n586) );
  XNOR2_X1 U658 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U659 ( .A(KEYINPUT71), .B(n588), .ZN(n590) );
  NAND2_X1 U660 ( .A1(n657), .A2(G68), .ZN(n589) );
  NAND2_X1 U661 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U662 ( .A(KEYINPUT13), .B(n591), .ZN(n597) );
  NAND2_X1 U663 ( .A1(G56), .A2(n658), .ZN(n592) );
  XOR2_X1 U664 ( .A(KEYINPUT14), .B(n592), .Z(n595) );
  NAND2_X1 U665 ( .A1(G43), .A2(n665), .ZN(n593) );
  XNOR2_X1 U666 ( .A(KEYINPUT73), .B(n593), .ZN(n594) );
  NOR2_X1 U667 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U668 ( .A1(n597), .A2(n596), .ZN(n934) );
  INV_X1 U669 ( .A(G860), .ZN(n622) );
  OR2_X1 U670 ( .A1(n934), .A2(n622), .ZN(G153) );
  XOR2_X1 U671 ( .A(G171), .B(KEYINPUT74), .Z(G301) );
  NAND2_X1 U672 ( .A1(G868), .A2(G301), .ZN(n598) );
  XNOR2_X1 U673 ( .A(n598), .B(KEYINPUT75), .ZN(n608) );
  NAND2_X1 U674 ( .A1(G79), .A2(n657), .ZN(n600) );
  NAND2_X1 U675 ( .A1(G54), .A2(n665), .ZN(n599) );
  NAND2_X1 U676 ( .A1(n600), .A2(n599), .ZN(n605) );
  NAND2_X1 U677 ( .A1(G92), .A2(n661), .ZN(n602) );
  NAND2_X1 U678 ( .A1(G66), .A2(n658), .ZN(n601) );
  NAND2_X1 U679 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U680 ( .A(KEYINPUT76), .B(n603), .ZN(n604) );
  NOR2_X1 U681 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X2 U682 ( .A(n606), .B(KEYINPUT15), .ZN(n922) );
  INV_X1 U683 ( .A(n922), .ZN(n629) );
  NOR2_X1 U684 ( .A1(n629), .A2(G868), .ZN(n607) );
  NOR2_X1 U685 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U686 ( .A(KEYINPUT77), .B(n609), .ZN(G284) );
  NAND2_X1 U687 ( .A1(G91), .A2(n661), .ZN(n610) );
  XNOR2_X1 U688 ( .A(n610), .B(KEYINPUT68), .ZN(n617) );
  NAND2_X1 U689 ( .A1(G78), .A2(n657), .ZN(n612) );
  NAND2_X1 U690 ( .A1(G65), .A2(n658), .ZN(n611) );
  NAND2_X1 U691 ( .A1(n612), .A2(n611), .ZN(n615) );
  NAND2_X1 U692 ( .A1(G53), .A2(n665), .ZN(n613) );
  XNOR2_X1 U693 ( .A(KEYINPUT69), .B(n613), .ZN(n614) );
  NOR2_X1 U694 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U695 ( .A1(n617), .A2(n616), .ZN(G299) );
  XNOR2_X1 U696 ( .A(KEYINPUT81), .B(G868), .ZN(n618) );
  NOR2_X1 U697 ( .A1(G286), .A2(n618), .ZN(n620) );
  NOR2_X1 U698 ( .A1(G868), .A2(G299), .ZN(n619) );
  NOR2_X1 U699 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U700 ( .A(KEYINPUT82), .B(n621), .ZN(G297) );
  NAND2_X1 U701 ( .A1(n622), .A2(G559), .ZN(n623) );
  NAND2_X1 U702 ( .A1(n623), .A2(n629), .ZN(n624) );
  XNOR2_X1 U703 ( .A(n624), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U704 ( .A1(G559), .A2(n922), .ZN(n625) );
  NAND2_X1 U705 ( .A1(G868), .A2(n625), .ZN(n626) );
  XNOR2_X1 U706 ( .A(n626), .B(KEYINPUT83), .ZN(n628) );
  NOR2_X1 U707 ( .A1(n934), .A2(G868), .ZN(n627) );
  NOR2_X1 U708 ( .A1(n628), .A2(n627), .ZN(G282) );
  NAND2_X1 U709 ( .A1(n629), .A2(G559), .ZN(n676) );
  XNOR2_X1 U710 ( .A(n934), .B(n676), .ZN(n630) );
  NOR2_X1 U711 ( .A1(n630), .A2(G860), .ZN(n637) );
  NAND2_X1 U712 ( .A1(G67), .A2(n658), .ZN(n632) );
  NAND2_X1 U713 ( .A1(G55), .A2(n665), .ZN(n631) );
  NAND2_X1 U714 ( .A1(n632), .A2(n631), .ZN(n636) );
  NAND2_X1 U715 ( .A1(G93), .A2(n661), .ZN(n634) );
  NAND2_X1 U716 ( .A1(G80), .A2(n657), .ZN(n633) );
  NAND2_X1 U717 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U718 ( .A1(n636), .A2(n635), .ZN(n670) );
  XNOR2_X1 U719 ( .A(n637), .B(n670), .ZN(G145) );
  NAND2_X1 U720 ( .A1(G49), .A2(n665), .ZN(n639) );
  NAND2_X1 U721 ( .A1(G74), .A2(G651), .ZN(n638) );
  NAND2_X1 U722 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U723 ( .A1(n658), .A2(n640), .ZN(n643) );
  NAND2_X1 U724 ( .A1(n641), .A2(G87), .ZN(n642) );
  NAND2_X1 U725 ( .A1(n643), .A2(n642), .ZN(G288) );
  NAND2_X1 U726 ( .A1(G86), .A2(n661), .ZN(n645) );
  NAND2_X1 U727 ( .A1(G61), .A2(n658), .ZN(n644) );
  NAND2_X1 U728 ( .A1(n645), .A2(n644), .ZN(n648) );
  NAND2_X1 U729 ( .A1(n657), .A2(G73), .ZN(n646) );
  XOR2_X1 U730 ( .A(KEYINPUT2), .B(n646), .Z(n647) );
  NOR2_X1 U731 ( .A1(n648), .A2(n647), .ZN(n650) );
  NAND2_X1 U732 ( .A1(n665), .A2(G48), .ZN(n649) );
  NAND2_X1 U733 ( .A1(n650), .A2(n649), .ZN(G305) );
  AND2_X1 U734 ( .A1(n658), .A2(G60), .ZN(n654) );
  NAND2_X1 U735 ( .A1(G85), .A2(n661), .ZN(n652) );
  NAND2_X1 U736 ( .A1(G72), .A2(n657), .ZN(n651) );
  NAND2_X1 U737 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U738 ( .A1(n654), .A2(n653), .ZN(n656) );
  NAND2_X1 U739 ( .A1(n665), .A2(G47), .ZN(n655) );
  NAND2_X1 U740 ( .A1(n656), .A2(n655), .ZN(G290) );
  NAND2_X1 U741 ( .A1(G75), .A2(n657), .ZN(n660) );
  NAND2_X1 U742 ( .A1(G62), .A2(n658), .ZN(n659) );
  NAND2_X1 U743 ( .A1(n660), .A2(n659), .ZN(n664) );
  NAND2_X1 U744 ( .A1(n661), .A2(G88), .ZN(n662) );
  XOR2_X1 U745 ( .A(KEYINPUT84), .B(n662), .Z(n663) );
  NOR2_X1 U746 ( .A1(n664), .A2(n663), .ZN(n667) );
  NAND2_X1 U747 ( .A1(n665), .A2(G50), .ZN(n666) );
  NAND2_X1 U748 ( .A1(n667), .A2(n666), .ZN(G303) );
  INV_X1 U749 ( .A(G303), .ZN(G166) );
  NOR2_X1 U750 ( .A1(n670), .A2(G868), .ZN(n668) );
  XOR2_X1 U751 ( .A(KEYINPUT86), .B(n668), .Z(n680) );
  XNOR2_X1 U752 ( .A(KEYINPUT19), .B(G299), .ZN(n669) );
  XNOR2_X1 U753 ( .A(n669), .B(G288), .ZN(n673) );
  XNOR2_X1 U754 ( .A(n670), .B(n934), .ZN(n671) );
  XNOR2_X1 U755 ( .A(n671), .B(G305), .ZN(n672) );
  XNOR2_X1 U756 ( .A(n673), .B(n672), .ZN(n675) );
  XNOR2_X1 U757 ( .A(G290), .B(G166), .ZN(n674) );
  XNOR2_X1 U758 ( .A(n675), .B(n674), .ZN(n844) );
  XOR2_X1 U759 ( .A(n844), .B(n676), .Z(n677) );
  NAND2_X1 U760 ( .A1(G868), .A2(n677), .ZN(n678) );
  XOR2_X1 U761 ( .A(KEYINPUT85), .B(n678), .Z(n679) );
  NAND2_X1 U762 ( .A1(n680), .A2(n679), .ZN(G295) );
  NAND2_X1 U763 ( .A1(G2078), .A2(G2084), .ZN(n681) );
  XOR2_X1 U764 ( .A(KEYINPUT20), .B(n681), .Z(n682) );
  NAND2_X1 U765 ( .A1(G2090), .A2(n682), .ZN(n683) );
  XNOR2_X1 U766 ( .A(KEYINPUT21), .B(n683), .ZN(n684) );
  NAND2_X1 U767 ( .A1(n684), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U768 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U769 ( .A1(G69), .A2(G120), .ZN(n685) );
  NOR2_X1 U770 ( .A1(G237), .A2(n685), .ZN(n686) );
  NAND2_X1 U771 ( .A1(G108), .A2(n686), .ZN(n890) );
  NAND2_X1 U772 ( .A1(G567), .A2(n890), .ZN(n687) );
  XNOR2_X1 U773 ( .A(KEYINPUT89), .B(n687), .ZN(n694) );
  XOR2_X1 U774 ( .A(KEYINPUT22), .B(KEYINPUT87), .Z(n689) );
  NAND2_X1 U775 ( .A1(G132), .A2(G82), .ZN(n688) );
  XNOR2_X1 U776 ( .A(n689), .B(n688), .ZN(n690) );
  NOR2_X1 U777 ( .A1(n690), .A2(G218), .ZN(n691) );
  NAND2_X1 U778 ( .A1(G96), .A2(n691), .ZN(n889) );
  NAND2_X1 U779 ( .A1(G2106), .A2(n889), .ZN(n692) );
  XOR2_X1 U780 ( .A(KEYINPUT88), .B(n692), .Z(n693) );
  NOR2_X1 U781 ( .A1(n694), .A2(n693), .ZN(G319) );
  INV_X1 U782 ( .A(G319), .ZN(n911) );
  NAND2_X1 U783 ( .A1(G661), .A2(G483), .ZN(n695) );
  NOR2_X1 U784 ( .A1(n911), .A2(n695), .ZN(n843) );
  NAND2_X1 U785 ( .A1(G36), .A2(n843), .ZN(n696) );
  XNOR2_X1 U786 ( .A(n696), .B(KEYINPUT90), .ZN(G176) );
  NAND2_X1 U787 ( .A1(n697), .A2(G40), .ZN(n698) );
  XNOR2_X1 U788 ( .A(n793), .B(KEYINPUT95), .ZN(n699) );
  NOR2_X1 U789 ( .A1(G164), .A2(G1384), .ZN(n794) );
  NAND2_X1 U790 ( .A1(G8), .A2(n724), .ZN(n769) );
  NOR2_X1 U791 ( .A1(G1966), .A2(n769), .ZN(n757) );
  NOR2_X1 U792 ( .A1(n757), .A2(n751), .ZN(n701) );
  XNOR2_X1 U793 ( .A(n700), .B(KEYINPUT97), .ZN(n760) );
  XNOR2_X1 U794 ( .A(n702), .B(KEYINPUT30), .ZN(n703) );
  INV_X1 U795 ( .A(n703), .ZN(n704) );
  NOR2_X1 U796 ( .A1(n704), .A2(G168), .ZN(n709) );
  INV_X1 U797 ( .A(n724), .ZN(n727) );
  NOR2_X1 U798 ( .A1(n727), .A2(G1961), .ZN(n705) );
  XOR2_X1 U799 ( .A(KEYINPUT98), .B(n705), .Z(n707) );
  XNOR2_X1 U800 ( .A(G2078), .B(KEYINPUT25), .ZN(n974) );
  NAND2_X1 U801 ( .A1(n727), .A2(n974), .ZN(n706) );
  NAND2_X1 U802 ( .A1(n707), .A2(n706), .ZN(n740) );
  NOR2_X1 U803 ( .A1(G171), .A2(n740), .ZN(n708) );
  NOR2_X1 U804 ( .A1(n709), .A2(n708), .ZN(n711) );
  XNOR2_X1 U805 ( .A(n711), .B(n710), .ZN(n744) );
  INV_X1 U806 ( .A(G1996), .ZN(n977) );
  NOR2_X1 U807 ( .A1(n724), .A2(n977), .ZN(n713) );
  XNOR2_X1 U808 ( .A(n713), .B(n712), .ZN(n715) );
  NAND2_X1 U809 ( .A1(n746), .A2(G1341), .ZN(n714) );
  NAND2_X1 U810 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U811 ( .A1(n934), .A2(n716), .ZN(n720) );
  NAND2_X1 U812 ( .A1(G1348), .A2(n746), .ZN(n718) );
  NAND2_X1 U813 ( .A1(G2067), .A2(n727), .ZN(n717) );
  NAND2_X1 U814 ( .A1(n718), .A2(n717), .ZN(n721) );
  NOR2_X1 U815 ( .A1(n922), .A2(n721), .ZN(n719) );
  NAND2_X1 U816 ( .A1(n922), .A2(n721), .ZN(n722) );
  NAND2_X1 U817 ( .A1(n723), .A2(n722), .ZN(n731) );
  INV_X1 U818 ( .A(G299), .ZN(n733) );
  INV_X1 U819 ( .A(n724), .ZN(n725) );
  NAND2_X1 U820 ( .A1(n725), .A2(G2072), .ZN(n726) );
  XNOR2_X1 U821 ( .A(n726), .B(KEYINPUT27), .ZN(n729) );
  INV_X1 U822 ( .A(G1956), .ZN(n909) );
  NOR2_X1 U823 ( .A1(n909), .A2(n727), .ZN(n728) );
  NOR2_X1 U824 ( .A1(n729), .A2(n728), .ZN(n732) );
  NAND2_X1 U825 ( .A1(n733), .A2(n732), .ZN(n730) );
  NAND2_X1 U826 ( .A1(n731), .A2(n730), .ZN(n737) );
  NOR2_X1 U827 ( .A1(n733), .A2(n732), .ZN(n735) );
  XNOR2_X1 U828 ( .A(KEYINPUT28), .B(KEYINPUT99), .ZN(n734) );
  XNOR2_X1 U829 ( .A(n735), .B(n734), .ZN(n736) );
  NAND2_X1 U830 ( .A1(n737), .A2(n736), .ZN(n739) );
  INV_X1 U831 ( .A(KEYINPUT29), .ZN(n738) );
  XNOR2_X1 U832 ( .A(n739), .B(n738), .ZN(n742) );
  NAND2_X1 U833 ( .A1(n740), .A2(G171), .ZN(n741) );
  NAND2_X1 U834 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U835 ( .A1(n744), .A2(n743), .ZN(n756) );
  AND2_X1 U836 ( .A1(G286), .A2(G8), .ZN(n745) );
  NAND2_X1 U837 ( .A1(n756), .A2(n745), .ZN(n753) );
  INV_X1 U838 ( .A(G8), .ZN(n751) );
  NOR2_X1 U839 ( .A1(G1971), .A2(n769), .ZN(n748) );
  NOR2_X1 U840 ( .A1(G2090), .A2(n746), .ZN(n747) );
  NOR2_X1 U841 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U842 ( .A1(n749), .A2(G303), .ZN(n750) );
  OR2_X1 U843 ( .A1(n751), .A2(n750), .ZN(n752) );
  XOR2_X1 U844 ( .A(KEYINPUT101), .B(KEYINPUT32), .Z(n754) );
  XNOR2_X1 U845 ( .A(n755), .B(n754), .ZN(n765) );
  XNOR2_X1 U846 ( .A(n756), .B(KEYINPUT100), .ZN(n759) );
  INV_X1 U847 ( .A(n757), .ZN(n758) );
  AND2_X1 U848 ( .A1(n759), .A2(n758), .ZN(n763) );
  INV_X1 U849 ( .A(n760), .ZN(n761) );
  NAND2_X1 U850 ( .A1(G8), .A2(n761), .ZN(n762) );
  NAND2_X1 U851 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U852 ( .A1(n765), .A2(n764), .ZN(n782) );
  NOR2_X1 U853 ( .A1(G1976), .A2(G288), .ZN(n775) );
  NOR2_X1 U854 ( .A1(G1971), .A2(G303), .ZN(n766) );
  NOR2_X1 U855 ( .A1(n775), .A2(n766), .ZN(n931) );
  NAND2_X1 U856 ( .A1(n782), .A2(n931), .ZN(n767) );
  NAND2_X1 U857 ( .A1(G1976), .A2(G288), .ZN(n937) );
  NAND2_X1 U858 ( .A1(n767), .A2(n937), .ZN(n768) );
  XNOR2_X1 U859 ( .A(n768), .B(KEYINPUT102), .ZN(n770) );
  BUF_X1 U860 ( .A(n769), .Z(n788) );
  NOR2_X1 U861 ( .A1(n770), .A2(n788), .ZN(n771) );
  XNOR2_X1 U862 ( .A(n771), .B(KEYINPUT64), .ZN(n772) );
  XNOR2_X1 U863 ( .A(n774), .B(n773), .ZN(n778) );
  NAND2_X1 U864 ( .A1(n775), .A2(KEYINPUT33), .ZN(n776) );
  NOR2_X1 U865 ( .A1(n788), .A2(n776), .ZN(n777) );
  XNOR2_X1 U866 ( .A(n779), .B(KEYINPUT104), .ZN(n781) );
  XNOR2_X1 U867 ( .A(G1981), .B(G305), .ZN(n924) );
  INV_X1 U868 ( .A(n924), .ZN(n780) );
  NAND2_X1 U869 ( .A1(n781), .A2(n780), .ZN(n792) );
  NOR2_X1 U870 ( .A1(G2090), .A2(G303), .ZN(n783) );
  NAND2_X1 U871 ( .A1(G8), .A2(n783), .ZN(n784) );
  NAND2_X1 U872 ( .A1(n782), .A2(n784), .ZN(n785) );
  NAND2_X1 U873 ( .A1(n785), .A2(n788), .ZN(n790) );
  NOR2_X1 U874 ( .A1(G1981), .A2(G305), .ZN(n786) );
  XOR2_X1 U875 ( .A(n786), .B(KEYINPUT24), .Z(n787) );
  XNOR2_X1 U876 ( .A(KEYINPUT96), .B(n787), .ZN(n789) );
  NAND2_X1 U877 ( .A1(n792), .A2(n791), .ZN(n824) );
  XNOR2_X1 U878 ( .A(G1986), .B(G290), .ZN(n929) );
  NOR2_X1 U879 ( .A1(n793), .A2(n794), .ZN(n834) );
  NAND2_X1 U880 ( .A1(n929), .A2(n834), .ZN(n822) );
  NAND2_X1 U881 ( .A1(G95), .A2(n875), .ZN(n796) );
  NAND2_X1 U882 ( .A1(G131), .A2(n574), .ZN(n795) );
  NAND2_X1 U883 ( .A1(n796), .A2(n795), .ZN(n800) );
  NAND2_X1 U884 ( .A1(G107), .A2(n879), .ZN(n798) );
  NAND2_X1 U885 ( .A1(G119), .A2(n880), .ZN(n797) );
  NAND2_X1 U886 ( .A1(n798), .A2(n797), .ZN(n799) );
  OR2_X1 U887 ( .A1(n800), .A2(n799), .ZN(n855) );
  AND2_X1 U888 ( .A1(n855), .A2(G1991), .ZN(n809) );
  NAND2_X1 U889 ( .A1(G117), .A2(n879), .ZN(n802) );
  NAND2_X1 U890 ( .A1(G141), .A2(n574), .ZN(n801) );
  NAND2_X1 U891 ( .A1(n802), .A2(n801), .ZN(n805) );
  NAND2_X1 U892 ( .A1(n875), .A2(G105), .ZN(n803) );
  XOR2_X1 U893 ( .A(KEYINPUT38), .B(n803), .Z(n804) );
  NOR2_X1 U894 ( .A1(n805), .A2(n804), .ZN(n807) );
  NAND2_X1 U895 ( .A1(n880), .A2(G129), .ZN(n806) );
  NAND2_X1 U896 ( .A1(n807), .A2(n806), .ZN(n871) );
  AND2_X1 U897 ( .A1(G1996), .A2(n871), .ZN(n808) );
  NOR2_X1 U898 ( .A1(n809), .A2(n808), .ZN(n1004) );
  XNOR2_X1 U899 ( .A(KEYINPUT93), .B(n834), .ZN(n810) );
  NOR2_X1 U900 ( .A1(n1004), .A2(n810), .ZN(n827) );
  XOR2_X1 U901 ( .A(KEYINPUT94), .B(n827), .Z(n820) );
  NAND2_X1 U902 ( .A1(G104), .A2(n875), .ZN(n812) );
  NAND2_X1 U903 ( .A1(G140), .A2(n574), .ZN(n811) );
  NAND2_X1 U904 ( .A1(n812), .A2(n811), .ZN(n813) );
  XNOR2_X1 U905 ( .A(KEYINPUT34), .B(n813), .ZN(n818) );
  NAND2_X1 U906 ( .A1(G116), .A2(n879), .ZN(n815) );
  NAND2_X1 U907 ( .A1(G128), .A2(n880), .ZN(n814) );
  NAND2_X1 U908 ( .A1(n815), .A2(n814), .ZN(n816) );
  XOR2_X1 U909 ( .A(KEYINPUT35), .B(n816), .Z(n817) );
  NOR2_X1 U910 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U911 ( .A(KEYINPUT36), .B(n819), .ZN(n859) );
  XNOR2_X1 U912 ( .A(KEYINPUT37), .B(G2067), .ZN(n832) );
  NOR2_X1 U913 ( .A1(n859), .A2(n832), .ZN(n1016) );
  NAND2_X1 U914 ( .A1(n834), .A2(n1016), .ZN(n830) );
  AND2_X1 U915 ( .A1(n820), .A2(n830), .ZN(n821) );
  AND2_X1 U916 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U917 ( .A1(n824), .A2(n823), .ZN(n837) );
  NOR2_X1 U918 ( .A1(G1996), .A2(n871), .ZN(n1011) );
  NOR2_X1 U919 ( .A1(G1991), .A2(n855), .ZN(n1000) );
  NOR2_X1 U920 ( .A1(G1986), .A2(G290), .ZN(n825) );
  NOR2_X1 U921 ( .A1(n1000), .A2(n825), .ZN(n826) );
  NOR2_X1 U922 ( .A1(n827), .A2(n826), .ZN(n828) );
  NOR2_X1 U923 ( .A1(n1011), .A2(n828), .ZN(n829) );
  XNOR2_X1 U924 ( .A(n829), .B(KEYINPUT39), .ZN(n831) );
  NAND2_X1 U925 ( .A1(n831), .A2(n830), .ZN(n833) );
  NAND2_X1 U926 ( .A1(n859), .A2(n832), .ZN(n1013) );
  NAND2_X1 U927 ( .A1(n833), .A2(n1013), .ZN(n835) );
  NAND2_X1 U928 ( .A1(n835), .A2(n834), .ZN(n836) );
  NAND2_X1 U929 ( .A1(n837), .A2(n836), .ZN(n839) );
  XOR2_X1 U930 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n838) );
  XNOR2_X1 U931 ( .A(n839), .B(n838), .ZN(G329) );
  NAND2_X1 U932 ( .A1(G2106), .A2(n840), .ZN(G217) );
  AND2_X1 U933 ( .A1(G15), .A2(G2), .ZN(n841) );
  NAND2_X1 U934 ( .A1(G661), .A2(n841), .ZN(G259) );
  NAND2_X1 U935 ( .A1(G3), .A2(G1), .ZN(n842) );
  NAND2_X1 U936 ( .A1(n843), .A2(n842), .ZN(G188) );
  XNOR2_X1 U937 ( .A(G286), .B(n844), .ZN(n845) );
  XNOR2_X1 U938 ( .A(n845), .B(n922), .ZN(n846) );
  XOR2_X1 U939 ( .A(G171), .B(n846), .Z(n914) );
  NOR2_X1 U940 ( .A1(G37), .A2(n914), .ZN(G397) );
  NAND2_X1 U941 ( .A1(G124), .A2(n880), .ZN(n847) );
  XNOR2_X1 U942 ( .A(n847), .B(KEYINPUT44), .ZN(n850) );
  NAND2_X1 U943 ( .A1(G112), .A2(n879), .ZN(n848) );
  XNOR2_X1 U944 ( .A(n848), .B(KEYINPUT108), .ZN(n849) );
  NAND2_X1 U945 ( .A1(n850), .A2(n849), .ZN(n854) );
  NAND2_X1 U946 ( .A1(G100), .A2(n875), .ZN(n852) );
  NAND2_X1 U947 ( .A1(G136), .A2(n574), .ZN(n851) );
  NAND2_X1 U948 ( .A1(n852), .A2(n851), .ZN(n853) );
  NOR2_X1 U949 ( .A1(n854), .A2(n853), .ZN(G162) );
  XOR2_X1 U950 ( .A(KEYINPUT48), .B(KEYINPUT111), .Z(n857) );
  XOR2_X1 U951 ( .A(G164), .B(n855), .Z(n856) );
  XNOR2_X1 U952 ( .A(n857), .B(n856), .ZN(n858) );
  XNOR2_X1 U953 ( .A(KEYINPUT46), .B(n858), .ZN(n861) );
  XNOR2_X1 U954 ( .A(n859), .B(KEYINPUT112), .ZN(n860) );
  XNOR2_X1 U955 ( .A(n861), .B(n860), .ZN(n870) );
  NAND2_X1 U956 ( .A1(G103), .A2(n875), .ZN(n863) );
  NAND2_X1 U957 ( .A1(G139), .A2(n574), .ZN(n862) );
  NAND2_X1 U958 ( .A1(n863), .A2(n862), .ZN(n869) );
  NAND2_X1 U959 ( .A1(n880), .A2(G127), .ZN(n864) );
  XNOR2_X1 U960 ( .A(n864), .B(KEYINPUT110), .ZN(n866) );
  NAND2_X1 U961 ( .A1(G115), .A2(n879), .ZN(n865) );
  NAND2_X1 U962 ( .A1(n866), .A2(n865), .ZN(n867) );
  XOR2_X1 U963 ( .A(KEYINPUT47), .B(n867), .Z(n868) );
  NOR2_X1 U964 ( .A1(n869), .A2(n868), .ZN(n1005) );
  XOR2_X1 U965 ( .A(n870), .B(n1005), .Z(n873) );
  XOR2_X1 U966 ( .A(G160), .B(n871), .Z(n872) );
  XNOR2_X1 U967 ( .A(n873), .B(n872), .ZN(n874) );
  XNOR2_X1 U968 ( .A(G162), .B(n874), .ZN(n888) );
  NAND2_X1 U969 ( .A1(G106), .A2(n875), .ZN(n877) );
  NAND2_X1 U970 ( .A1(G142), .A2(n574), .ZN(n876) );
  NAND2_X1 U971 ( .A1(n877), .A2(n876), .ZN(n878) );
  XNOR2_X1 U972 ( .A(n878), .B(KEYINPUT45), .ZN(n885) );
  NAND2_X1 U973 ( .A1(G118), .A2(n879), .ZN(n882) );
  NAND2_X1 U974 ( .A1(G130), .A2(n880), .ZN(n881) );
  NAND2_X1 U975 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U976 ( .A(KEYINPUT109), .B(n883), .ZN(n884) );
  NAND2_X1 U977 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U978 ( .A(n886), .B(n998), .ZN(n887) );
  XOR2_X1 U979 ( .A(n888), .B(n887), .Z(n913) );
  NOR2_X1 U980 ( .A1(G37), .A2(n913), .ZN(G395) );
  INV_X1 U982 ( .A(G132), .ZN(G219) );
  INV_X1 U983 ( .A(G120), .ZN(G236) );
  INV_X1 U984 ( .A(G96), .ZN(G221) );
  INV_X1 U985 ( .A(G82), .ZN(G220) );
  INV_X1 U986 ( .A(G69), .ZN(G235) );
  NOR2_X1 U987 ( .A1(n890), .A2(n889), .ZN(G325) );
  INV_X1 U988 ( .A(G325), .ZN(G261) );
  XOR2_X1 U989 ( .A(G2096), .B(KEYINPUT43), .Z(n892) );
  XNOR2_X1 U990 ( .A(G2067), .B(G2678), .ZN(n891) );
  XNOR2_X1 U991 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U992 ( .A(n893), .B(KEYINPUT42), .Z(n895) );
  XNOR2_X1 U993 ( .A(G2072), .B(G2090), .ZN(n894) );
  XNOR2_X1 U994 ( .A(n895), .B(n894), .ZN(n899) );
  XOR2_X1 U995 ( .A(KEYINPUT106), .B(G2100), .Z(n897) );
  XNOR2_X1 U996 ( .A(G2078), .B(G2084), .ZN(n896) );
  XNOR2_X1 U997 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U998 ( .A(n899), .B(n898), .ZN(G227) );
  XOR2_X1 U999 ( .A(G1981), .B(G1961), .Z(n901) );
  XNOR2_X1 U1000 ( .A(G1986), .B(G1966), .ZN(n900) );
  XNOR2_X1 U1001 ( .A(n901), .B(n900), .ZN(n905) );
  XOR2_X1 U1002 ( .A(G1976), .B(G1971), .Z(n903) );
  XNOR2_X1 U1003 ( .A(G1996), .B(G1991), .ZN(n902) );
  XNOR2_X1 U1004 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1005 ( .A(n905), .B(n904), .Z(n907) );
  XNOR2_X1 U1006 ( .A(KEYINPUT107), .B(G2474), .ZN(n906) );
  XNOR2_X1 U1007 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1008 ( .A(KEYINPUT41), .B(n908), .ZN(n910) );
  XNOR2_X1 U1009 ( .A(n910), .B(n909), .ZN(G229) );
  NOR2_X1 U1010 ( .A1(n911), .A2(G401), .ZN(n912) );
  XNOR2_X1 U1011 ( .A(n912), .B(KEYINPUT113), .ZN(n918) );
  AND2_X1 U1012 ( .A1(n914), .A2(n913), .ZN(n915) );
  NOR2_X1 U1013 ( .A1(G37), .A2(n915), .ZN(n916) );
  XNOR2_X1 U1014 ( .A(n916), .B(KEYINPUT114), .ZN(n917) );
  NOR2_X1 U1015 ( .A1(n918), .A2(n917), .ZN(n921) );
  NOR2_X1 U1016 ( .A1(G227), .A2(G229), .ZN(n919) );
  XOR2_X1 U1017 ( .A(KEYINPUT49), .B(n919), .Z(n920) );
  NAND2_X1 U1018 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1021 ( .A(G16), .B(KEYINPUT56), .ZN(n944) );
  XNOR2_X1 U1022 ( .A(n922), .B(G1348), .ZN(n927) );
  XOR2_X1 U1023 ( .A(G1966), .B(G168), .Z(n923) );
  NOR2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1025 ( .A(KEYINPUT57), .B(n925), .ZN(n926) );
  NOR2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n942) );
  XNOR2_X1 U1027 ( .A(G1956), .B(G299), .ZN(n928) );
  NOR2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n940) );
  XNOR2_X1 U1030 ( .A(G171), .B(G1961), .ZN(n933) );
  NAND2_X1 U1031 ( .A1(G1971), .A2(G303), .ZN(n932) );
  NAND2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n936) );
  XNOR2_X1 U1033 ( .A(G1341), .B(n934), .ZN(n935) );
  NOR2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n938) );
  NAND2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1037 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1038 ( .A1(n944), .A2(n943), .ZN(n1030) );
  XOR2_X1 U1039 ( .A(G1966), .B(G21), .Z(n956) );
  XNOR2_X1 U1040 ( .A(KEYINPUT123), .B(G1341), .ZN(n945) );
  XNOR2_X1 U1041 ( .A(n945), .B(G19), .ZN(n951) );
  XOR2_X1 U1042 ( .A(KEYINPUT124), .B(G4), .Z(n947) );
  XNOR2_X1 U1043 ( .A(G1348), .B(KEYINPUT59), .ZN(n946) );
  XNOR2_X1 U1044 ( .A(n947), .B(n946), .ZN(n949) );
  XNOR2_X1 U1045 ( .A(G1981), .B(G6), .ZN(n948) );
  NOR2_X1 U1046 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n953) );
  XNOR2_X1 U1048 ( .A(G20), .B(G1956), .ZN(n952) );
  NOR2_X1 U1049 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1050 ( .A(KEYINPUT60), .B(n954), .ZN(n955) );
  NAND2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n969) );
  XNOR2_X1 U1052 ( .A(KEYINPUT125), .B(G1971), .ZN(n957) );
  XNOR2_X1 U1053 ( .A(n957), .B(G22), .ZN(n962) );
  XNOR2_X1 U1054 ( .A(G1976), .B(KEYINPUT126), .ZN(n958) );
  XNOR2_X1 U1055 ( .A(n958), .B(G23), .ZN(n960) );
  XNOR2_X1 U1056 ( .A(G24), .B(G1986), .ZN(n959) );
  NOR2_X1 U1057 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1059 ( .A(n963), .B(KEYINPUT58), .ZN(n964) );
  XNOR2_X1 U1060 ( .A(n964), .B(KEYINPUT127), .ZN(n967) );
  XOR2_X1 U1061 ( .A(G1961), .B(KEYINPUT122), .Z(n965) );
  XNOR2_X1 U1062 ( .A(G5), .B(n965), .ZN(n966) );
  NAND2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1065 ( .A(KEYINPUT61), .B(n970), .ZN(n972) );
  INV_X1 U1066 ( .A(G16), .ZN(n971) );
  NAND2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1068 ( .A1(n973), .A2(G11), .ZN(n1028) );
  XOR2_X1 U1069 ( .A(n974), .B(G27), .Z(n976) );
  XNOR2_X1 U1070 ( .A(G1991), .B(G25), .ZN(n975) );
  NOR2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n985) );
  XNOR2_X1 U1072 ( .A(G32), .B(n977), .ZN(n978) );
  NAND2_X1 U1073 ( .A1(n978), .A2(G28), .ZN(n983) );
  XNOR2_X1 U1074 ( .A(G2067), .B(G26), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(G2072), .B(G33), .ZN(n979) );
  NOR2_X1 U1076 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1077 ( .A(n981), .B(KEYINPUT117), .ZN(n982) );
  NOR2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1079 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1080 ( .A(n986), .B(KEYINPUT53), .ZN(n987) );
  XNOR2_X1 U1081 ( .A(KEYINPUT118), .B(n987), .ZN(n994) );
  XNOR2_X1 U1082 ( .A(G2090), .B(G35), .ZN(n992) );
  XOR2_X1 U1083 ( .A(G34), .B(KEYINPUT120), .Z(n989) );
  XNOR2_X1 U1084 ( .A(G2084), .B(KEYINPUT54), .ZN(n988) );
  XNOR2_X1 U1085 ( .A(n989), .B(n988), .ZN(n990) );
  XNOR2_X1 U1086 ( .A(n990), .B(KEYINPUT119), .ZN(n991) );
  NOR2_X1 U1087 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1088 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1089 ( .A(KEYINPUT55), .B(n995), .ZN(n996) );
  NOR2_X1 U1090 ( .A1(G29), .A2(n996), .ZN(n997) );
  XNOR2_X1 U1091 ( .A(n997), .B(KEYINPUT121), .ZN(n1026) );
  XNOR2_X1 U1092 ( .A(G160), .B(G2084), .ZN(n999) );
  NAND2_X1 U1093 ( .A1(n999), .A2(n998), .ZN(n1001) );
  NOR2_X1 U1094 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1095 ( .A(KEYINPUT115), .B(n1002), .Z(n1003) );
  NAND2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1020) );
  XOR2_X1 U1097 ( .A(G2072), .B(n1005), .Z(n1007) );
  XOR2_X1 U1098 ( .A(G164), .B(G2078), .Z(n1006) );
  NOR2_X1 U1099 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1100 ( .A(KEYINPUT50), .B(n1008), .ZN(n1009) );
  XNOR2_X1 U1101 ( .A(n1009), .B(KEYINPUT116), .ZN(n1018) );
  XOR2_X1 U1102 ( .A(G2090), .B(G162), .Z(n1010) );
  NOR2_X1 U1103 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1104 ( .A(KEYINPUT51), .B(n1012), .Z(n1014) );
  NAND2_X1 U1105 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1106 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1109 ( .A(n1021), .B(KEYINPUT52), .ZN(n1023) );
  INV_X1 U1110 ( .A(KEYINPUT55), .ZN(n1022) );
  NAND2_X1 U1111 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1112 ( .A1(G29), .A2(n1024), .ZN(n1025) );
  NAND2_X1 U1113 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1116 ( .A(KEYINPUT62), .B(n1031), .Z(G311) );
  INV_X1 U1117 ( .A(G311), .ZN(G150) );
endmodule

