

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587;

  NOR2_X1 U323 ( .A1(n523), .A2(n472), .ZN(n569) );
  XNOR2_X1 U324 ( .A(n438), .B(n437), .ZN(n447) );
  AND2_X1 U325 ( .A1(n399), .A2(n523), .ZN(n378) );
  INV_X1 U326 ( .A(n349), .ZN(n346) );
  XOR2_X1 U327 ( .A(KEYINPUT94), .B(n403), .Z(n523) );
  XOR2_X1 U328 ( .A(G176GAT), .B(G120GAT), .Z(n291) );
  XOR2_X1 U329 ( .A(KEYINPUT103), .B(n452), .Z(n292) );
  XNOR2_X1 U330 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n455) );
  XNOR2_X1 U331 ( .A(n436), .B(n291), .ZN(n437) );
  XNOR2_X1 U332 ( .A(n445), .B(n444), .ZN(n446) );
  AND2_X1 U333 ( .A1(n569), .A2(n473), .ZN(n475) );
  XNOR2_X1 U334 ( .A(KEYINPUT48), .B(KEYINPUT114), .ZN(n467) );
  NOR2_X1 U335 ( .A1(n585), .A2(n406), .ZN(n408) );
  XNOR2_X1 U336 ( .A(n345), .B(G197GAT), .ZN(n349) );
  XNOR2_X1 U337 ( .A(n447), .B(n446), .ZN(n451) );
  XNOR2_X1 U338 ( .A(n378), .B(KEYINPUT95), .ZN(n532) );
  NAND2_X1 U339 ( .A1(n405), .A2(n404), .ZN(n486) );
  XOR2_X1 U340 ( .A(n451), .B(n450), .Z(n463) );
  XNOR2_X1 U341 ( .A(n479), .B(n478), .ZN(n566) );
  XOR2_X1 U342 ( .A(n391), .B(n390), .Z(n534) );
  XOR2_X1 U343 ( .A(n361), .B(n360), .Z(n525) );
  XNOR2_X1 U344 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U345 ( .A(G36GAT), .B(KEYINPUT104), .ZN(n453) );
  XNOR2_X1 U346 ( .A(n483), .B(n482), .ZN(G1351GAT) );
  XNOR2_X1 U347 ( .A(n454), .B(n453), .ZN(G1329GAT) );
  XOR2_X1 U348 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n294) );
  XNOR2_X1 U349 ( .A(G85GAT), .B(KEYINPUT64), .ZN(n293) );
  XNOR2_X1 U350 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U351 ( .A(n295), .B(G92GAT), .Z(n297) );
  XOR2_X1 U352 ( .A(G106GAT), .B(KEYINPUT72), .Z(n442) );
  XNOR2_X1 U353 ( .A(G218GAT), .B(n442), .ZN(n296) );
  XNOR2_X1 U354 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U355 ( .A(G50GAT), .B(KEYINPUT76), .Z(n335) );
  XOR2_X1 U356 ( .A(n298), .B(n335), .Z(n301) );
  XNOR2_X1 U357 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n299) );
  XNOR2_X1 U358 ( .A(n299), .B(KEYINPUT7), .ZN(n415) );
  XOR2_X1 U359 ( .A(G43GAT), .B(G134GAT), .Z(n383) );
  XNOR2_X1 U360 ( .A(n415), .B(n383), .ZN(n300) );
  XNOR2_X1 U361 ( .A(n301), .B(n300), .ZN(n310) );
  XOR2_X1 U362 ( .A(KEYINPUT78), .B(KEYINPUT10), .Z(n303) );
  XNOR2_X1 U363 ( .A(G162GAT), .B(KEYINPUT77), .ZN(n302) );
  XNOR2_X1 U364 ( .A(n303), .B(n302), .ZN(n308) );
  XNOR2_X1 U365 ( .A(G36GAT), .B(G190GAT), .ZN(n304) );
  XNOR2_X1 U366 ( .A(n304), .B(KEYINPUT79), .ZN(n353) );
  XOR2_X1 U367 ( .A(n353), .B(G99GAT), .Z(n306) );
  NAND2_X1 U368 ( .A1(G232GAT), .A2(G233GAT), .ZN(n305) );
  XNOR2_X1 U369 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U370 ( .A(n308), .B(n307), .Z(n309) );
  XOR2_X1 U371 ( .A(n310), .B(n309), .Z(n544) );
  XOR2_X1 U372 ( .A(KEYINPUT36), .B(n544), .Z(n585) );
  XOR2_X1 U373 ( .A(G8GAT), .B(KEYINPUT80), .Z(n350) );
  XOR2_X1 U374 ( .A(G22GAT), .B(G78GAT), .Z(n334) );
  XOR2_X1 U375 ( .A(n350), .B(n334), .Z(n312) );
  XNOR2_X1 U376 ( .A(G155GAT), .B(G211GAT), .ZN(n311) );
  XNOR2_X1 U377 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U378 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n314) );
  NAND2_X1 U379 ( .A1(G231GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U380 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U381 ( .A(n316), .B(n315), .Z(n318) );
  XOR2_X1 U382 ( .A(G15GAT), .B(G1GAT), .Z(n412) );
  XNOR2_X1 U383 ( .A(n412), .B(KEYINPUT14), .ZN(n317) );
  XNOR2_X1 U384 ( .A(n318), .B(n317), .ZN(n326) );
  XOR2_X1 U385 ( .A(G57GAT), .B(G127GAT), .Z(n320) );
  XNOR2_X1 U386 ( .A(G183GAT), .B(G71GAT), .ZN(n319) );
  XNOR2_X1 U387 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U388 ( .A(KEYINPUT81), .B(KEYINPUT82), .Z(n322) );
  XNOR2_X1 U389 ( .A(KEYINPUT13), .B(G64GAT), .ZN(n321) );
  XNOR2_X1 U390 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U391 ( .A(n324), .B(n323), .Z(n325) );
  XOR2_X1 U392 ( .A(n326), .B(n325), .Z(n565) );
  INV_X1 U393 ( .A(n565), .ZN(n579) );
  XNOR2_X1 U394 ( .A(KEYINPUT28), .B(KEYINPUT65), .ZN(n348) );
  XOR2_X1 U395 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n328) );
  XNOR2_X1 U396 ( .A(G162GAT), .B(KEYINPUT89), .ZN(n327) );
  XNOR2_X1 U397 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U398 ( .A(n329), .B(G155GAT), .Z(n331) );
  XNOR2_X1 U399 ( .A(G141GAT), .B(G148GAT), .ZN(n330) );
  XNOR2_X1 U400 ( .A(n331), .B(n330), .ZN(n375) );
  XOR2_X1 U401 ( .A(KEYINPUT24), .B(KEYINPUT90), .Z(n333) );
  XNOR2_X1 U402 ( .A(G204GAT), .B(KEYINPUT22), .ZN(n332) );
  XNOR2_X1 U403 ( .A(n333), .B(n332), .ZN(n339) );
  XOR2_X1 U404 ( .A(KEYINPUT23), .B(G106GAT), .Z(n337) );
  XNOR2_X1 U405 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U406 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U407 ( .A(n339), .B(n338), .Z(n341) );
  NAND2_X1 U408 ( .A1(G228GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U409 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U410 ( .A(n375), .B(n342), .ZN(n347) );
  XOR2_X1 U411 ( .A(KEYINPUT21), .B(G218GAT), .Z(n344) );
  XNOR2_X1 U412 ( .A(KEYINPUT88), .B(G211GAT), .ZN(n343) );
  XNOR2_X1 U413 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U414 ( .A(n347), .B(n346), .Z(n473) );
  XNOR2_X1 U415 ( .A(n348), .B(n473), .ZN(n537) );
  XNOR2_X1 U416 ( .A(n350), .B(n349), .ZN(n352) );
  NAND2_X1 U417 ( .A1(G226GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U418 ( .A(n352), .B(n351), .ZN(n354) );
  XOR2_X1 U419 ( .A(n354), .B(n353), .Z(n361) );
  XNOR2_X1 U420 ( .A(G204GAT), .B(G92GAT), .ZN(n355) );
  XNOR2_X1 U421 ( .A(n355), .B(G64GAT), .ZN(n436) );
  XNOR2_X1 U422 ( .A(G183GAT), .B(KEYINPUT19), .ZN(n356) );
  XNOR2_X1 U423 ( .A(n356), .B(KEYINPUT18), .ZN(n357) );
  XOR2_X1 U424 ( .A(n357), .B(KEYINPUT17), .Z(n359) );
  XNOR2_X1 U425 ( .A(G169GAT), .B(G176GAT), .ZN(n358) );
  XNOR2_X1 U426 ( .A(n359), .B(n358), .ZN(n382) );
  XNOR2_X1 U427 ( .A(n436), .B(n382), .ZN(n360) );
  XNOR2_X1 U428 ( .A(n525), .B(KEYINPUT27), .ZN(n399) );
  XOR2_X1 U429 ( .A(G85GAT), .B(G57GAT), .Z(n431) );
  XOR2_X1 U430 ( .A(KEYINPUT91), .B(G134GAT), .Z(n363) );
  XNOR2_X1 U431 ( .A(G29GAT), .B(G1GAT), .ZN(n362) );
  XNOR2_X1 U432 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U433 ( .A(n431), .B(n364), .Z(n366) );
  NAND2_X1 U434 ( .A1(G225GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U435 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U436 ( .A(n367), .B(KEYINPUT1), .Z(n371) );
  XOR2_X1 U437 ( .A(G120GAT), .B(G127GAT), .Z(n369) );
  XNOR2_X1 U438 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n368) );
  XNOR2_X1 U439 ( .A(n369), .B(n368), .ZN(n384) );
  XNOR2_X1 U440 ( .A(n384), .B(KEYINPUT4), .ZN(n370) );
  XNOR2_X1 U441 ( .A(n371), .B(n370), .ZN(n377) );
  XOR2_X1 U442 ( .A(KEYINPUT6), .B(KEYINPUT93), .Z(n373) );
  XNOR2_X1 U443 ( .A(KEYINPUT5), .B(KEYINPUT92), .ZN(n372) );
  XNOR2_X1 U444 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U445 ( .A(n375), .B(n374), .Z(n376) );
  XOR2_X1 U446 ( .A(n377), .B(n376), .Z(n403) );
  NOR2_X1 U447 ( .A1(n537), .A2(n532), .ZN(n393) );
  XOR2_X1 U448 ( .A(KEYINPUT84), .B(KEYINPUT86), .Z(n380) );
  XNOR2_X1 U449 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n379) );
  XNOR2_X1 U450 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U451 ( .A(n382), .B(n381), .ZN(n391) );
  XOR2_X1 U452 ( .A(n384), .B(n383), .Z(n386) );
  NAND2_X1 U453 ( .A1(G227GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U454 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U455 ( .A(G99GAT), .B(G71GAT), .Z(n443) );
  XOR2_X1 U456 ( .A(n387), .B(n443), .Z(n389) );
  XNOR2_X1 U457 ( .A(G190GAT), .B(KEYINPUT85), .ZN(n388) );
  XNOR2_X1 U458 ( .A(n389), .B(n388), .ZN(n390) );
  INV_X1 U459 ( .A(n534), .ZN(n477) );
  XOR2_X1 U460 ( .A(n477), .B(KEYINPUT87), .Z(n392) );
  NAND2_X1 U461 ( .A1(n393), .A2(n392), .ZN(n405) );
  NAND2_X1 U462 ( .A1(n534), .A2(n525), .ZN(n394) );
  NAND2_X1 U463 ( .A1(n394), .A2(n473), .ZN(n395) );
  XNOR2_X1 U464 ( .A(n395), .B(KEYINPUT97), .ZN(n396) );
  XNOR2_X1 U465 ( .A(n396), .B(KEYINPUT25), .ZN(n401) );
  NOR2_X1 U466 ( .A1(n534), .A2(n473), .ZN(n398) );
  XNOR2_X1 U467 ( .A(KEYINPUT96), .B(KEYINPUT26), .ZN(n397) );
  XNOR2_X1 U468 ( .A(n398), .B(n397), .ZN(n568) );
  NAND2_X1 U469 ( .A1(n568), .A2(n399), .ZN(n400) );
  NAND2_X1 U470 ( .A1(n401), .A2(n400), .ZN(n402) );
  NAND2_X1 U471 ( .A1(n403), .A2(n402), .ZN(n404) );
  NAND2_X1 U472 ( .A1(n579), .A2(n486), .ZN(n406) );
  XNOR2_X1 U473 ( .A(KEYINPUT102), .B(KEYINPUT37), .ZN(n407) );
  XNOR2_X1 U474 ( .A(n408), .B(n407), .ZN(n520) );
  XOR2_X1 U475 ( .A(G197GAT), .B(G22GAT), .Z(n410) );
  XNOR2_X1 U476 ( .A(G43GAT), .B(G141GAT), .ZN(n409) );
  XNOR2_X1 U477 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U478 ( .A(n411), .B(G36GAT), .Z(n414) );
  XNOR2_X1 U479 ( .A(n412), .B(G50GAT), .ZN(n413) );
  XNOR2_X1 U480 ( .A(n414), .B(n413), .ZN(n419) );
  XOR2_X1 U481 ( .A(n415), .B(KEYINPUT67), .Z(n417) );
  NAND2_X1 U482 ( .A1(G229GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U483 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U484 ( .A(n419), .B(n418), .Z(n427) );
  XOR2_X1 U485 ( .A(KEYINPUT69), .B(KEYINPUT66), .Z(n421) );
  XNOR2_X1 U486 ( .A(G169GAT), .B(G113GAT), .ZN(n420) );
  XNOR2_X1 U487 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U488 ( .A(G8GAT), .B(KEYINPUT30), .Z(n423) );
  XNOR2_X1 U489 ( .A(KEYINPUT68), .B(KEYINPUT29), .ZN(n422) );
  XNOR2_X1 U490 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U491 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U492 ( .A(n427), .B(n426), .Z(n570) );
  INV_X1 U493 ( .A(n570), .ZN(n558) );
  XOR2_X1 U494 ( .A(KEYINPUT32), .B(KEYINPUT73), .Z(n429) );
  XNOR2_X1 U495 ( .A(G148GAT), .B(G78GAT), .ZN(n428) );
  XNOR2_X1 U496 ( .A(n429), .B(n428), .ZN(n433) );
  INV_X1 U497 ( .A(n433), .ZN(n430) );
  NAND2_X1 U498 ( .A1(n430), .A2(n431), .ZN(n435) );
  INV_X1 U499 ( .A(n431), .ZN(n432) );
  NAND2_X1 U500 ( .A1(n433), .A2(n432), .ZN(n434) );
  NAND2_X1 U501 ( .A1(n435), .A2(n434), .ZN(n438) );
  XOR2_X1 U502 ( .A(KEYINPUT74), .B(KEYINPUT33), .Z(n440) );
  NAND2_X1 U503 ( .A1(G230GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U504 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U505 ( .A(KEYINPUT71), .B(n441), .ZN(n445) );
  XNOR2_X1 U506 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U507 ( .A(KEYINPUT31), .B(KEYINPUT70), .Z(n449) );
  XNOR2_X1 U508 ( .A(KEYINPUT75), .B(KEYINPUT13), .ZN(n448) );
  XNOR2_X1 U509 ( .A(n449), .B(n448), .ZN(n450) );
  INV_X1 U510 ( .A(n463), .ZN(n576) );
  NAND2_X1 U511 ( .A1(n558), .A2(n576), .ZN(n488) );
  NOR2_X1 U512 ( .A1(n520), .A2(n488), .ZN(n452) );
  XNOR2_X1 U513 ( .A(KEYINPUT38), .B(n292), .ZN(n507) );
  NAND2_X1 U514 ( .A1(n507), .A2(n525), .ZN(n454) );
  INV_X1 U515 ( .A(KEYINPUT119), .ZN(n479) );
  XOR2_X1 U516 ( .A(KEYINPUT41), .B(n463), .Z(n509) );
  NAND2_X1 U517 ( .A1(n509), .A2(n558), .ZN(n456) );
  XNOR2_X1 U518 ( .A(n456), .B(n455), .ZN(n457) );
  NAND2_X1 U519 ( .A1(n457), .A2(n579), .ZN(n458) );
  XNOR2_X1 U520 ( .A(n458), .B(KEYINPUT113), .ZN(n459) );
  INV_X1 U521 ( .A(n544), .ZN(n556) );
  NAND2_X1 U522 ( .A1(n459), .A2(n556), .ZN(n460) );
  XNOR2_X1 U523 ( .A(n460), .B(KEYINPUT47), .ZN(n466) );
  NOR2_X1 U524 ( .A1(n585), .A2(n579), .ZN(n461) );
  XNOR2_X1 U525 ( .A(KEYINPUT45), .B(n461), .ZN(n462) );
  NAND2_X1 U526 ( .A1(n462), .A2(n570), .ZN(n464) );
  NOR2_X1 U527 ( .A1(n464), .A2(n463), .ZN(n465) );
  NOR2_X1 U528 ( .A1(n466), .A2(n465), .ZN(n468) );
  XNOR2_X1 U529 ( .A(n468), .B(n467), .ZN(n533) );
  XNOR2_X1 U530 ( .A(KEYINPUT117), .B(n525), .ZN(n469) );
  NOR2_X1 U531 ( .A1(n533), .A2(n469), .ZN(n471) );
  INV_X1 U532 ( .A(KEYINPUT54), .ZN(n470) );
  XNOR2_X1 U533 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U534 ( .A(KEYINPUT55), .B(KEYINPUT118), .ZN(n474) );
  XNOR2_X1 U535 ( .A(n475), .B(n474), .ZN(n476) );
  NOR2_X1 U536 ( .A1(n477), .A2(n476), .ZN(n478) );
  NAND2_X1 U537 ( .A1(n566), .A2(n544), .ZN(n483) );
  XOR2_X1 U538 ( .A(KEYINPUT122), .B(KEYINPUT58), .Z(n481) );
  INV_X1 U539 ( .A(G190GAT), .ZN(n480) );
  NAND2_X1 U540 ( .A1(n556), .A2(n565), .ZN(n484) );
  XNOR2_X1 U541 ( .A(n484), .B(KEYINPUT16), .ZN(n485) );
  XNOR2_X1 U542 ( .A(n485), .B(KEYINPUT83), .ZN(n487) );
  NAND2_X1 U543 ( .A1(n487), .A2(n486), .ZN(n511) );
  NOR2_X1 U544 ( .A1(n488), .A2(n511), .ZN(n497) );
  NAND2_X1 U545 ( .A1(n497), .A2(n523), .ZN(n489) );
  XNOR2_X1 U546 ( .A(n489), .B(KEYINPUT34), .ZN(n490) );
  XNOR2_X1 U547 ( .A(G1GAT), .B(n490), .ZN(G1324GAT) );
  XOR2_X1 U548 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n492) );
  NAND2_X1 U549 ( .A1(n497), .A2(n525), .ZN(n491) );
  XNOR2_X1 U550 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U551 ( .A(G8GAT), .B(n493), .ZN(G1325GAT) );
  XOR2_X1 U552 ( .A(KEYINPUT35), .B(KEYINPUT100), .Z(n495) );
  NAND2_X1 U553 ( .A1(n497), .A2(n534), .ZN(n494) );
  XNOR2_X1 U554 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U555 ( .A(G15GAT), .B(n496), .ZN(G1326GAT) );
  NAND2_X1 U556 ( .A1(n537), .A2(n497), .ZN(n498) );
  XNOR2_X1 U557 ( .A(n498), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U558 ( .A1(n507), .A2(n523), .ZN(n501) );
  XNOR2_X1 U559 ( .A(G29GAT), .B(KEYINPUT101), .ZN(n499) );
  XNOR2_X1 U560 ( .A(n499), .B(KEYINPUT39), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n501), .B(n500), .ZN(G1328GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n503) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(KEYINPUT106), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n503), .B(n502), .ZN(n504) );
  XOR2_X1 U565 ( .A(KEYINPUT105), .B(n504), .Z(n506) );
  NAND2_X1 U566 ( .A1(n507), .A2(n534), .ZN(n505) );
  XNOR2_X1 U567 ( .A(n506), .B(n505), .ZN(G1330GAT) );
  NAND2_X1 U568 ( .A1(n507), .A2(n537), .ZN(n508) );
  XNOR2_X1 U569 ( .A(n508), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U570 ( .A(KEYINPUT42), .B(KEYINPUT109), .Z(n513) );
  NAND2_X1 U571 ( .A1(n570), .A2(n509), .ZN(n510) );
  XNOR2_X1 U572 ( .A(n510), .B(KEYINPUT108), .ZN(n521) );
  NOR2_X1 U573 ( .A1(n521), .A2(n511), .ZN(n517) );
  NAND2_X1 U574 ( .A1(n517), .A2(n523), .ZN(n512) );
  XNOR2_X1 U575 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U576 ( .A(G57GAT), .B(n514), .ZN(G1332GAT) );
  NAND2_X1 U577 ( .A1(n525), .A2(n517), .ZN(n515) );
  XNOR2_X1 U578 ( .A(n515), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U579 ( .A1(n534), .A2(n517), .ZN(n516) );
  XNOR2_X1 U580 ( .A(n516), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U581 ( .A(G78GAT), .B(KEYINPUT43), .Z(n519) );
  NAND2_X1 U582 ( .A1(n517), .A2(n537), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n519), .B(n518), .ZN(G1335GAT) );
  NOR2_X1 U584 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U585 ( .A(n522), .B(KEYINPUT110), .ZN(n528) );
  NAND2_X1 U586 ( .A1(n528), .A2(n523), .ZN(n524) );
  XNOR2_X1 U587 ( .A(n524), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U588 ( .A1(n528), .A2(n525), .ZN(n526) );
  XNOR2_X1 U589 ( .A(n526), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U590 ( .A1(n528), .A2(n534), .ZN(n527) );
  XNOR2_X1 U591 ( .A(n527), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT111), .B(KEYINPUT44), .Z(n530) );
  NAND2_X1 U593 ( .A1(n528), .A2(n537), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  NOR2_X1 U596 ( .A1(n533), .A2(n532), .ZN(n548) );
  NAND2_X1 U597 ( .A1(n548), .A2(n534), .ZN(n535) );
  XOR2_X1 U598 ( .A(KEYINPUT115), .B(n535), .Z(n536) );
  NOR2_X1 U599 ( .A1(n537), .A2(n536), .ZN(n545) );
  NAND2_X1 U600 ( .A1(n545), .A2(n558), .ZN(n538) );
  XNOR2_X1 U601 ( .A(n538), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n540) );
  NAND2_X1 U603 ( .A1(n545), .A2(n509), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U605 ( .A(G120GAT), .B(n541), .ZN(G1341GAT) );
  NAND2_X1 U606 ( .A1(n545), .A2(n565), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n542), .B(KEYINPUT50), .ZN(n543) );
  XNOR2_X1 U608 ( .A(G127GAT), .B(n543), .ZN(G1342GAT) );
  XOR2_X1 U609 ( .A(G134GAT), .B(KEYINPUT51), .Z(n547) );
  NAND2_X1 U610 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  NAND2_X1 U612 ( .A1(n548), .A2(n568), .ZN(n555) );
  NOR2_X1 U613 ( .A1(n570), .A2(n555), .ZN(n549) );
  XOR2_X1 U614 ( .A(G141GAT), .B(n549), .Z(G1344GAT) );
  INV_X1 U615 ( .A(n509), .ZN(n550) );
  NOR2_X1 U616 ( .A1(n550), .A2(n555), .ZN(n552) );
  XNOR2_X1 U617 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(n553), .ZN(G1345GAT) );
  NOR2_X1 U620 ( .A1(n579), .A2(n555), .ZN(n554) );
  XOR2_X1 U621 ( .A(G155GAT), .B(n554), .Z(G1346GAT) );
  NOR2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U623 ( .A(G162GAT), .B(n557), .Z(G1347GAT) );
  XNOR2_X1 U624 ( .A(G169GAT), .B(KEYINPUT120), .ZN(n560) );
  NAND2_X1 U625 ( .A1(n558), .A2(n566), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(G1348GAT) );
  NAND2_X1 U627 ( .A1(n566), .A2(n509), .ZN(n562) );
  XOR2_X1 U628 ( .A(KEYINPUT57), .B(KEYINPUT56), .Z(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n564) );
  XOR2_X1 U630 ( .A(G176GAT), .B(KEYINPUT121), .Z(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(G1349GAT) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n584) );
  NOR2_X1 U635 ( .A1(n570), .A2(n584), .ZN(n575) );
  XOR2_X1 U636 ( .A(KEYINPUT60), .B(KEYINPUT124), .Z(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(KEYINPUT123), .B(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1352GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n584), .ZN(n578) );
  XNOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  NOR2_X1 U644 ( .A1(n579), .A2(n584), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G211GAT), .B(KEYINPUT125), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1354GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n583) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(n587) );
  NOR2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U651 ( .A(n587), .B(n586), .Z(G1355GAT) );
endmodule

