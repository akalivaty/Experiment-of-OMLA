

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578;

  INV_X1 U321 ( .A(n572), .ZN(n486) );
  XNOR2_X1 U322 ( .A(n304), .B(n303), .ZN(n305) );
  NAND2_X1 U323 ( .A1(n404), .A2(n563), .ZN(n406) );
  XNOR2_X2 U324 ( .A(n306), .B(n305), .ZN(n568) );
  NOR2_X2 U325 ( .A1(n461), .A2(n561), .ZN(n450) );
  XNOR2_X1 U326 ( .A(n568), .B(n307), .ZN(n404) );
  NOR2_X1 U327 ( .A1(n541), .A2(n458), .ZN(n524) );
  NOR2_X1 U328 ( .A1(n576), .A2(n487), .ZN(n489) );
  XOR2_X1 U329 ( .A(n425), .B(n424), .Z(n516) );
  XNOR2_X1 U330 ( .A(KEYINPUT45), .B(KEYINPUT117), .ZN(n383) );
  XNOR2_X1 U331 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U332 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U333 ( .A(KEYINPUT123), .B(KEYINPUT54), .ZN(n427) );
  XNOR2_X1 U334 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U335 ( .A(n428), .B(n427), .ZN(n449) );
  XNOR2_X1 U336 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U337 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U338 ( .A(n492), .B(n491), .ZN(n501) );
  INV_X1 U339 ( .A(KEYINPUT40), .ZN(n498) );
  XNOR2_X1 U340 ( .A(n453), .B(G176GAT), .ZN(n454) );
  XNOR2_X1 U341 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U342 ( .A(n455), .B(n454), .ZN(G1349GAT) );
  XOR2_X1 U343 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n290) );
  XNOR2_X1 U344 ( .A(KEYINPUT75), .B(KEYINPUT73), .ZN(n289) );
  XOR2_X1 U345 ( .A(n290), .B(n289), .Z(n306) );
  XNOR2_X1 U346 ( .A(G71GAT), .B(G57GAT), .ZN(n291) );
  XNOR2_X1 U347 ( .A(n291), .B(KEYINPUT13), .ZN(n349) );
  XOR2_X1 U348 ( .A(KEYINPUT76), .B(n349), .Z(n293) );
  NAND2_X1 U349 ( .A1(G230GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U350 ( .A(n293), .B(n292), .ZN(n296) );
  XOR2_X1 U351 ( .A(G64GAT), .B(G92GAT), .Z(n295) );
  XNOR2_X1 U352 ( .A(G176GAT), .B(G204GAT), .ZN(n294) );
  XNOR2_X1 U353 ( .A(n295), .B(n294), .ZN(n415) );
  XOR2_X1 U354 ( .A(n296), .B(n415), .Z(n299) );
  XNOR2_X1 U355 ( .A(G106GAT), .B(G78GAT), .ZN(n297) );
  XNOR2_X1 U356 ( .A(n297), .B(G148GAT), .ZN(n337) );
  XNOR2_X1 U357 ( .A(G120GAT), .B(n337), .ZN(n298) );
  XNOR2_X1 U358 ( .A(n299), .B(n298), .ZN(n301) );
  INV_X1 U359 ( .A(KEYINPUT72), .ZN(n300) );
  XNOR2_X1 U360 ( .A(n301), .B(n300), .ZN(n304) );
  XNOR2_X1 U361 ( .A(G99GAT), .B(G85GAT), .ZN(n302) );
  XNOR2_X1 U362 ( .A(n302), .B(KEYINPUT74), .ZN(n378) );
  XNOR2_X1 U363 ( .A(n378), .B(KEYINPUT32), .ZN(n303) );
  XOR2_X1 U364 ( .A(KEYINPUT64), .B(KEYINPUT41), .Z(n307) );
  XOR2_X1 U365 ( .A(KEYINPUT111), .B(n404), .Z(n529) );
  XOR2_X1 U366 ( .A(KEYINPUT88), .B(KEYINPUT17), .Z(n309) );
  XNOR2_X1 U367 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n308) );
  XNOR2_X1 U368 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U369 ( .A(G169GAT), .B(n310), .Z(n419) );
  XOR2_X1 U370 ( .A(G183GAT), .B(KEYINPUT85), .Z(n312) );
  XNOR2_X1 U371 ( .A(KEYINPUT90), .B(KEYINPUT89), .ZN(n311) );
  XNOR2_X1 U372 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U373 ( .A(G176GAT), .B(KEYINPUT20), .Z(n314) );
  XNOR2_X1 U374 ( .A(KEYINPUT87), .B(KEYINPUT86), .ZN(n313) );
  XNOR2_X1 U375 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U376 ( .A(n316), .B(n315), .Z(n329) );
  XOR2_X1 U377 ( .A(KEYINPUT84), .B(KEYINPUT0), .Z(n318) );
  XNOR2_X1 U378 ( .A(G134GAT), .B(KEYINPUT83), .ZN(n317) );
  XNOR2_X1 U379 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U380 ( .A(n319), .B(KEYINPUT82), .Z(n321) );
  XNOR2_X1 U381 ( .A(G113GAT), .B(G120GAT), .ZN(n320) );
  XNOR2_X1 U382 ( .A(n321), .B(n320), .ZN(n440) );
  XOR2_X1 U383 ( .A(G15GAT), .B(G127GAT), .Z(n355) );
  XOR2_X1 U384 ( .A(G71GAT), .B(G99GAT), .Z(n323) );
  XNOR2_X1 U385 ( .A(G43GAT), .B(G190GAT), .ZN(n322) );
  XNOR2_X1 U386 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U387 ( .A(n355), .B(n324), .Z(n326) );
  NAND2_X1 U388 ( .A1(G227GAT), .A2(G233GAT), .ZN(n325) );
  XNOR2_X1 U389 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U390 ( .A(n440), .B(n327), .ZN(n328) );
  XNOR2_X1 U391 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U392 ( .A(n419), .B(n330), .ZN(n526) );
  XOR2_X1 U393 ( .A(G204GAT), .B(KEYINPUT23), .Z(n332) );
  XNOR2_X1 U394 ( .A(KEYINPUT93), .B(KEYINPUT24), .ZN(n331) );
  XNOR2_X1 U395 ( .A(n332), .B(n331), .ZN(n346) );
  XOR2_X1 U396 ( .A(KEYINPUT91), .B(KEYINPUT22), .Z(n334) );
  NAND2_X1 U397 ( .A1(G228GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U398 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U399 ( .A(n335), .B(G211GAT), .Z(n339) );
  XNOR2_X1 U400 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n336) );
  XNOR2_X1 U401 ( .A(n336), .B(KEYINPUT2), .ZN(n429) );
  XNOR2_X1 U402 ( .A(n337), .B(n429), .ZN(n338) );
  XNOR2_X1 U403 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U404 ( .A(G22GAT), .B(G155GAT), .Z(n354) );
  XOR2_X1 U405 ( .A(n340), .B(n354), .Z(n344) );
  XOR2_X1 U406 ( .A(G50GAT), .B(G162GAT), .Z(n377) );
  XOR2_X1 U407 ( .A(KEYINPUT92), .B(KEYINPUT21), .Z(n342) );
  XNOR2_X1 U408 ( .A(G197GAT), .B(G218GAT), .ZN(n341) );
  XNOR2_X1 U409 ( .A(n342), .B(n341), .ZN(n417) );
  XNOR2_X1 U410 ( .A(n377), .B(n417), .ZN(n343) );
  XNOR2_X1 U411 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U412 ( .A(n346), .B(n345), .Z(n461) );
  XOR2_X1 U413 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n348) );
  XNOR2_X1 U414 ( .A(KEYINPUT12), .B(KEYINPUT14), .ZN(n347) );
  XNOR2_X1 U415 ( .A(n348), .B(n347), .ZN(n362) );
  XNOR2_X1 U416 ( .A(G8GAT), .B(G183GAT), .ZN(n350) );
  XNOR2_X1 U417 ( .A(n350), .B(G211GAT), .ZN(n414) );
  XOR2_X1 U418 ( .A(n414), .B(KEYINPUT15), .Z(n352) );
  NAND2_X1 U419 ( .A1(G231GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U420 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U421 ( .A(n349), .B(n353), .Z(n357) );
  XNOR2_X1 U422 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U423 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U424 ( .A(n358), .B(G64GAT), .ZN(n360) );
  XOR2_X1 U425 ( .A(KEYINPUT71), .B(G1GAT), .Z(n391) );
  XOR2_X1 U426 ( .A(n391), .B(G78GAT), .Z(n359) );
  XNOR2_X1 U427 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U428 ( .A(n362), .B(n361), .ZN(n572) );
  XOR2_X1 U429 ( .A(KEYINPUT70), .B(KEYINPUT8), .Z(n364) );
  XNOR2_X1 U430 ( .A(G43GAT), .B(G29GAT), .ZN(n363) );
  XNOR2_X1 U431 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U432 ( .A(KEYINPUT7), .B(n365), .Z(n398) );
  XOR2_X1 U433 ( .A(G92GAT), .B(G218GAT), .Z(n367) );
  XNOR2_X1 U434 ( .A(G134GAT), .B(G106GAT), .ZN(n366) );
  XNOR2_X1 U435 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U436 ( .A(KEYINPUT78), .B(KEYINPUT77), .Z(n369) );
  XNOR2_X1 U437 ( .A(KEYINPUT65), .B(KEYINPUT66), .ZN(n368) );
  XNOR2_X1 U438 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U439 ( .A(n371), .B(n370), .Z(n376) );
  XOR2_X1 U440 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n373) );
  NAND2_X1 U441 ( .A1(G232GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U442 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U443 ( .A(KEYINPUT9), .B(n374), .ZN(n375) );
  XNOR2_X1 U444 ( .A(n376), .B(n375), .ZN(n381) );
  XOR2_X1 U445 ( .A(G36GAT), .B(G190GAT), .Z(n421) );
  XOR2_X1 U446 ( .A(n377), .B(n421), .Z(n379) );
  XOR2_X1 U447 ( .A(n398), .B(n382), .Z(n558) );
  XOR2_X1 U448 ( .A(KEYINPUT36), .B(n558), .Z(n576) );
  NOR2_X1 U449 ( .A1(n486), .A2(n576), .ZN(n384) );
  NOR2_X1 U450 ( .A1(n385), .A2(n568), .ZN(n403) );
  XOR2_X1 U451 ( .A(KEYINPUT68), .B(G8GAT), .Z(n387) );
  XNOR2_X1 U452 ( .A(G197GAT), .B(G22GAT), .ZN(n386) );
  XNOR2_X1 U453 ( .A(n387), .B(n386), .ZN(n402) );
  XOR2_X1 U454 ( .A(G141GAT), .B(G113GAT), .Z(n389) );
  XNOR2_X1 U455 ( .A(G50GAT), .B(G36GAT), .ZN(n388) );
  XNOR2_X1 U456 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U457 ( .A(n390), .B(G15GAT), .Z(n393) );
  XNOR2_X1 U458 ( .A(G169GAT), .B(n391), .ZN(n392) );
  XNOR2_X1 U459 ( .A(n393), .B(n392), .ZN(n397) );
  XOR2_X1 U460 ( .A(KEYINPUT69), .B(KEYINPUT30), .Z(n395) );
  NAND2_X1 U461 ( .A1(G229GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U462 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U463 ( .A(n397), .B(n396), .Z(n400) );
  XNOR2_X1 U464 ( .A(n398), .B(KEYINPUT29), .ZN(n399) );
  XNOR2_X1 U465 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U466 ( .A(n402), .B(n401), .ZN(n544) );
  NAND2_X1 U467 ( .A1(n403), .A2(n544), .ZN(n412) );
  INV_X1 U468 ( .A(n544), .ZN(n563) );
  XOR2_X1 U469 ( .A(KEYINPUT46), .B(KEYINPUT115), .Z(n405) );
  XNOR2_X1 U470 ( .A(n406), .B(n405), .ZN(n408) );
  XOR2_X1 U471 ( .A(KEYINPUT114), .B(n486), .Z(n554) );
  NOR2_X1 U472 ( .A1(n554), .A2(n558), .ZN(n407) );
  NAND2_X1 U473 ( .A1(n408), .A2(n407), .ZN(n410) );
  XOR2_X1 U474 ( .A(KEYINPUT116), .B(KEYINPUT47), .Z(n409) );
  XNOR2_X1 U475 ( .A(n410), .B(n409), .ZN(n411) );
  NAND2_X1 U476 ( .A1(n412), .A2(n411), .ZN(n413) );
  XNOR2_X1 U477 ( .A(n413), .B(KEYINPUT48), .ZN(n543) );
  XNOR2_X1 U478 ( .A(n415), .B(n414), .ZN(n425) );
  XOR2_X1 U479 ( .A(KEYINPUT99), .B(KEYINPUT98), .Z(n416) );
  XOR2_X1 U480 ( .A(n421), .B(n420), .Z(n423) );
  NAND2_X1 U481 ( .A1(G226GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U482 ( .A(n423), .B(n422), .ZN(n424) );
  INV_X1 U483 ( .A(n516), .ZN(n426) );
  NAND2_X1 U484 ( .A1(n543), .A2(n426), .ZN(n428) );
  XNOR2_X1 U485 ( .A(n429), .B(KEYINPUT97), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n430), .B(KEYINPUT94), .ZN(n434) );
  XOR2_X1 U487 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n432) );
  XNOR2_X1 U488 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n431) );
  XNOR2_X1 U489 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U490 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U491 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n436) );
  XNOR2_X1 U492 ( .A(G1GAT), .B(G57GAT), .ZN(n435) );
  XNOR2_X1 U493 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U494 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U495 ( .A(n440), .B(n439), .ZN(n448) );
  NAND2_X1 U496 ( .A1(G225GAT), .A2(G233GAT), .ZN(n446) );
  XOR2_X1 U497 ( .A(G85GAT), .B(G155GAT), .Z(n442) );
  XNOR2_X1 U498 ( .A(G127GAT), .B(G148GAT), .ZN(n441) );
  XNOR2_X1 U499 ( .A(n442), .B(n441), .ZN(n444) );
  XOR2_X1 U500 ( .A(G29GAT), .B(G162GAT), .Z(n443) );
  XNOR2_X1 U501 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U502 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U503 ( .A(n448), .B(n447), .ZN(n513) );
  NAND2_X1 U504 ( .A1(n449), .A2(n513), .ZN(n561) );
  XNOR2_X1 U505 ( .A(n450), .B(KEYINPUT55), .ZN(n451) );
  NOR2_X1 U506 ( .A1(n526), .A2(n451), .ZN(n452) );
  XNOR2_X1 U507 ( .A(KEYINPUT124), .B(n452), .ZN(n557) );
  NAND2_X1 U508 ( .A1(n529), .A2(n557), .ZN(n455) );
  XOR2_X1 U509 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n453) );
  NOR2_X1 U510 ( .A1(n568), .A2(n544), .ZN(n490) );
  XNOR2_X1 U511 ( .A(n516), .B(KEYINPUT27), .ZN(n464) );
  NOR2_X1 U512 ( .A1(n464), .A2(n513), .ZN(n456) );
  XOR2_X1 U513 ( .A(KEYINPUT100), .B(n456), .Z(n541) );
  XOR2_X1 U514 ( .A(n461), .B(KEYINPUT67), .Z(n457) );
  XOR2_X1 U515 ( .A(KEYINPUT28), .B(n457), .Z(n520) );
  INV_X1 U516 ( .A(n520), .ZN(n458) );
  NAND2_X1 U517 ( .A1(n524), .A2(n526), .ZN(n470) );
  NOR2_X1 U518 ( .A1(n526), .A2(n516), .ZN(n459) );
  NOR2_X1 U519 ( .A1(n461), .A2(n459), .ZN(n460) );
  XOR2_X1 U520 ( .A(KEYINPUT25), .B(n460), .Z(n466) );
  XOR2_X1 U521 ( .A(KEYINPUT101), .B(KEYINPUT26), .Z(n463) );
  NAND2_X1 U522 ( .A1(n461), .A2(n526), .ZN(n462) );
  XNOR2_X1 U523 ( .A(n463), .B(n462), .ZN(n562) );
  NOR2_X1 U524 ( .A1(n562), .A2(n464), .ZN(n465) );
  NOR2_X1 U525 ( .A1(n466), .A2(n465), .ZN(n467) );
  XOR2_X1 U526 ( .A(KEYINPUT102), .B(n467), .Z(n468) );
  NAND2_X1 U527 ( .A1(n468), .A2(n513), .ZN(n469) );
  NAND2_X1 U528 ( .A1(n470), .A2(n469), .ZN(n485) );
  NOR2_X1 U529 ( .A1(n486), .A2(n558), .ZN(n471) );
  XNOR2_X1 U530 ( .A(n471), .B(KEYINPUT16), .ZN(n472) );
  XOR2_X1 U531 ( .A(KEYINPUT81), .B(n472), .Z(n473) );
  AND2_X1 U532 ( .A1(n485), .A2(n473), .ZN(n503) );
  NAND2_X1 U533 ( .A1(n490), .A2(n503), .ZN(n482) );
  NOR2_X1 U534 ( .A1(n513), .A2(n482), .ZN(n475) );
  XNOR2_X1 U535 ( .A(KEYINPUT103), .B(KEYINPUT34), .ZN(n474) );
  XNOR2_X1 U536 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U537 ( .A(G1GAT), .B(n476), .ZN(G1324GAT) );
  NOR2_X1 U538 ( .A1(n516), .A2(n482), .ZN(n477) );
  XOR2_X1 U539 ( .A(G8GAT), .B(n477), .Z(G1325GAT) );
  NOR2_X1 U540 ( .A1(n482), .A2(n526), .ZN(n481) );
  XOR2_X1 U541 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n479) );
  XNOR2_X1 U542 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n478) );
  XNOR2_X1 U543 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U544 ( .A(n481), .B(n480), .ZN(G1326GAT) );
  NOR2_X1 U545 ( .A1(n520), .A2(n482), .ZN(n483) );
  XOR2_X1 U546 ( .A(KEYINPUT106), .B(n483), .Z(n484) );
  XNOR2_X1 U547 ( .A(G22GAT), .B(n484), .ZN(G1327GAT) );
  NAND2_X1 U548 ( .A1(n486), .A2(n485), .ZN(n487) );
  XNOR2_X1 U549 ( .A(KEYINPUT107), .B(KEYINPUT37), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n489), .B(n488), .ZN(n512) );
  NAND2_X1 U551 ( .A1(n512), .A2(n490), .ZN(n492) );
  XNOR2_X1 U552 ( .A(KEYINPUT108), .B(KEYINPUT38), .ZN(n491) );
  NOR2_X1 U553 ( .A1(n513), .A2(n501), .ZN(n494) );
  XNOR2_X1 U554 ( .A(KEYINPUT39), .B(KEYINPUT109), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U556 ( .A(G29GAT), .B(n495), .Z(G1328GAT) );
  NOR2_X1 U557 ( .A1(n516), .A2(n501), .ZN(n496) );
  XOR2_X1 U558 ( .A(KEYINPUT110), .B(n496), .Z(n497) );
  XNOR2_X1 U559 ( .A(G36GAT), .B(n497), .ZN(G1329GAT) );
  NOR2_X1 U560 ( .A1(n526), .A2(n501), .ZN(n499) );
  XNOR2_X1 U561 ( .A(G43GAT), .B(n500), .ZN(G1330GAT) );
  NOR2_X1 U562 ( .A1(n520), .A2(n501), .ZN(n502) );
  XOR2_X1 U563 ( .A(G50GAT), .B(n502), .Z(G1331GAT) );
  AND2_X1 U564 ( .A1(n544), .A2(n529), .ZN(n511) );
  NAND2_X1 U565 ( .A1(n511), .A2(n503), .ZN(n508) );
  NOR2_X1 U566 ( .A1(n513), .A2(n508), .ZN(n504) );
  XOR2_X1 U567 ( .A(G57GAT), .B(n504), .Z(n505) );
  XNOR2_X1 U568 ( .A(KEYINPUT42), .B(n505), .ZN(G1332GAT) );
  NOR2_X1 U569 ( .A1(n516), .A2(n508), .ZN(n506) );
  XOR2_X1 U570 ( .A(G64GAT), .B(n506), .Z(G1333GAT) );
  NOR2_X1 U571 ( .A1(n526), .A2(n508), .ZN(n507) );
  XOR2_X1 U572 ( .A(G71GAT), .B(n507), .Z(G1334GAT) );
  NOR2_X1 U573 ( .A1(n520), .A2(n508), .ZN(n510) );
  XNOR2_X1 U574 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n510), .B(n509), .ZN(G1335GAT) );
  NAND2_X1 U576 ( .A1(n512), .A2(n511), .ZN(n519) );
  NOR2_X1 U577 ( .A1(n513), .A2(n519), .ZN(n514) );
  XOR2_X1 U578 ( .A(KEYINPUT112), .B(n514), .Z(n515) );
  XNOR2_X1 U579 ( .A(G85GAT), .B(n515), .ZN(G1336GAT) );
  NOR2_X1 U580 ( .A1(n516), .A2(n519), .ZN(n517) );
  XOR2_X1 U581 ( .A(G92GAT), .B(n517), .Z(G1337GAT) );
  NOR2_X1 U582 ( .A1(n526), .A2(n519), .ZN(n518) );
  XOR2_X1 U583 ( .A(G99GAT), .B(n518), .Z(G1338GAT) );
  NOR2_X1 U584 ( .A1(n520), .A2(n519), .ZN(n522) );
  XNOR2_X1 U585 ( .A(KEYINPUT44), .B(KEYINPUT113), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U587 ( .A(G106GAT), .B(n523), .ZN(G1339GAT) );
  NAND2_X1 U588 ( .A1(n543), .A2(n524), .ZN(n525) );
  NOR2_X1 U589 ( .A1(n526), .A2(n525), .ZN(n538) );
  NAND2_X1 U590 ( .A1(n538), .A2(n563), .ZN(n527) );
  XNOR2_X1 U591 ( .A(n527), .B(KEYINPUT118), .ZN(n528) );
  XNOR2_X1 U592 ( .A(G113GAT), .B(n528), .ZN(G1340GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT49), .B(KEYINPUT120), .Z(n531) );
  NAND2_X1 U594 ( .A1(n538), .A2(n529), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n531), .B(n530), .ZN(n533) );
  XOR2_X1 U596 ( .A(G120GAT), .B(KEYINPUT119), .Z(n532) );
  XNOR2_X1 U597 ( .A(n533), .B(n532), .ZN(G1341GAT) );
  XNOR2_X1 U598 ( .A(G127GAT), .B(KEYINPUT122), .ZN(n537) );
  XOR2_X1 U599 ( .A(KEYINPUT50), .B(KEYINPUT121), .Z(n535) );
  NAND2_X1 U600 ( .A1(n538), .A2(n554), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(G1342GAT) );
  XOR2_X1 U603 ( .A(G134GAT), .B(KEYINPUT51), .Z(n540) );
  NAND2_X1 U604 ( .A1(n538), .A2(n558), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(G1343GAT) );
  NOR2_X1 U606 ( .A1(n562), .A2(n541), .ZN(n542) );
  NAND2_X1 U607 ( .A1(n543), .A2(n542), .ZN(n546) );
  NOR2_X1 U608 ( .A1(n544), .A2(n546), .ZN(n545) );
  XOR2_X1 U609 ( .A(G141GAT), .B(n545), .Z(G1344GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n548) );
  INV_X1 U611 ( .A(n546), .ZN(n551) );
  NAND2_X1 U612 ( .A1(n551), .A2(n404), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(n549), .ZN(G1345GAT) );
  NAND2_X1 U615 ( .A1(n572), .A2(n551), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n550), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U617 ( .A1(n551), .A2(n558), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n552), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U619 ( .A1(n557), .A2(n563), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U621 ( .A(G183GAT), .B(KEYINPUT125), .Z(n556) );
  NAND2_X1 U622 ( .A1(n554), .A2(n557), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(G1350GAT) );
  XNOR2_X1 U624 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n560) );
  NAND2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(G1351GAT) );
  XNOR2_X1 U627 ( .A(KEYINPUT59), .B(KEYINPUT126), .ZN(n567) );
  XOR2_X1 U628 ( .A(G197GAT), .B(KEYINPUT60), .Z(n565) );
  NOR2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n574) );
  NAND2_X1 U630 ( .A1(n574), .A2(n563), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(G1352GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n570) );
  NAND2_X1 U634 ( .A1(n574), .A2(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XOR2_X1 U636 ( .A(G204GAT), .B(n571), .Z(G1353GAT) );
  NAND2_X1 U637 ( .A1(n572), .A2(n574), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n573), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U639 ( .A(n574), .ZN(n575) );
  NOR2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U641 ( .A(KEYINPUT62), .B(n577), .Z(n578) );
  XNOR2_X1 U642 ( .A(G218GAT), .B(n578), .ZN(G1355GAT) );
endmodule

