

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795;

  INV_X1 U374 ( .A(n565), .ZN(n622) );
  NOR2_X1 U375 ( .A1(G953), .A2(G237), .ZN(n550) );
  XNOR2_X1 U376 ( .A(n388), .B(n380), .ZN(n700) );
  NOR2_X2 U377 ( .A1(n769), .A2(n768), .ZN(n770) );
  NOR2_X2 U378 ( .A1(n667), .A2(n768), .ZN(n669) );
  XNOR2_X2 U379 ( .A(n512), .B(n511), .ZN(n751) );
  XNOR2_X1 U380 ( .A(n522), .B(n521), .ZN(n593) );
  XNOR2_X1 U381 ( .A(n461), .B(n467), .ZN(n771) );
  XNOR2_X1 U382 ( .A(n479), .B(n478), .ZN(n513) );
  AND2_X1 U383 ( .A1(n365), .A2(n364), .ZN(n363) );
  NAND2_X1 U384 ( .A1(n370), .A2(n358), .ZN(n369) );
  NAND2_X1 U385 ( .A1(n394), .A2(n393), .ZN(n392) );
  NAND2_X1 U386 ( .A1(n564), .A2(n722), .ZN(n676) );
  AND2_X1 U387 ( .A1(n376), .A2(n375), .ZN(n374) );
  XNOR2_X1 U388 ( .A(n420), .B(KEYINPUT35), .ZN(n792) );
  NAND2_X1 U389 ( .A1(n373), .A2(n407), .ZN(n372) );
  XNOR2_X1 U390 ( .A(n442), .B(KEYINPUT31), .ZN(n718) );
  XNOR2_X1 U391 ( .A(n451), .B(n450), .ZN(n793) );
  XNOR2_X1 U392 ( .A(n403), .B(KEYINPUT39), .ZN(n653) );
  NOR2_X1 U393 ( .A1(n707), .A2(KEYINPUT103), .ZN(n407) );
  OR2_X1 U394 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U395 ( .A(n510), .B(n509), .ZN(n389) );
  NOR2_X1 U396 ( .A1(n728), .A2(n620), .ZN(n603) );
  XNOR2_X1 U397 ( .A(n452), .B(KEYINPUT38), .ZN(n736) );
  NAND2_X1 U398 ( .A1(n417), .A2(n413), .ZN(n577) );
  XOR2_X1 U399 ( .A(n765), .B(n764), .Z(n766) );
  AND2_X1 U400 ( .A1(n419), .A2(n418), .ZN(n417) );
  OR2_X1 U401 ( .A1(n678), .A2(G902), .ZN(n449) );
  XNOR2_X1 U402 ( .A(n443), .B(G134), .ZN(n541) );
  XNOR2_X1 U403 ( .A(n547), .B(n513), .ZN(n461) );
  XNOR2_X1 U404 ( .A(n514), .B(G113), .ZN(n547) );
  XNOR2_X1 U405 ( .A(n538), .B(KEYINPUT16), .ZN(n467) );
  XNOR2_X1 U406 ( .A(G122), .B(G104), .ZN(n514) );
  XNOR2_X1 U407 ( .A(KEYINPUT77), .B(G110), .ZN(n378) );
  XNOR2_X1 U408 ( .A(G119), .B(G101), .ZN(n479) );
  NOR2_X1 U409 ( .A1(n645), .A2(n473), .ZN(n408) );
  NAND2_X1 U410 ( .A1(n416), .A2(n415), .ZN(n414) );
  NOR2_X1 U411 ( .A1(n795), .A2(n793), .ZN(n615) );
  NAND2_X1 U412 ( .A1(n470), .A2(n457), .ZN(n368) );
  AND2_X1 U413 ( .A1(n658), .A2(n657), .ZN(n457) );
  XNOR2_X1 U414 ( .A(n371), .B(n406), .ZN(n588) );
  NAND2_X1 U415 ( .A1(n387), .A2(n574), .ZN(n386) );
  NAND2_X1 U416 ( .A1(n352), .A2(n676), .ZN(n387) );
  NAND2_X1 U417 ( .A1(n676), .A2(n351), .ZN(n385) );
  INV_X1 U418 ( .A(n728), .ZN(n390) );
  XNOR2_X1 U419 ( .A(n557), .B(n556), .ZN(n558) );
  BUF_X1 U420 ( .A(n577), .Z(n610) );
  XNOR2_X1 U421 ( .A(n402), .B(n480), .ZN(n401) );
  XNOR2_X1 U422 ( .A(n423), .B(n475), .ZN(n402) );
  NAND2_X1 U423 ( .A1(n456), .A2(n469), .ZN(n370) );
  NOR2_X1 U424 ( .A1(n656), .A2(n424), .ZN(n456) );
  XNOR2_X1 U425 ( .A(G902), .B(KEYINPUT15), .ZN(n519) );
  INV_X1 U426 ( .A(n792), .ZN(n468) );
  XNOR2_X1 U427 ( .A(n410), .B(n409), .ZN(n781) );
  XNOR2_X1 U428 ( .A(KEYINPUT73), .B(KEYINPUT10), .ZN(n409) );
  XNOR2_X1 U429 ( .A(n411), .B(G140), .ZN(n410) );
  INV_X1 U430 ( .A(G125), .ZN(n411) );
  XNOR2_X1 U431 ( .A(n624), .B(n623), .ZN(n647) );
  NOR2_X1 U432 ( .A1(n620), .A2(n621), .ZN(n412) );
  INV_X1 U433 ( .A(KEYINPUT102), .ZN(n454) );
  NAND2_X1 U434 ( .A1(n389), .A2(n390), .ZN(n455) );
  NAND2_X1 U435 ( .A1(n725), .A2(KEYINPUT110), .ZN(n471) );
  XNOR2_X1 U436 ( .A(n728), .B(n448), .ZN(n565) );
  XNOR2_X1 U437 ( .A(KEYINPUT109), .B(KEYINPUT6), .ZN(n448) );
  NAND2_X1 U438 ( .A1(n392), .A2(n391), .ZN(n398) );
  AND2_X1 U439 ( .A1(n396), .A2(n655), .ZN(n395) );
  XNOR2_X1 U440 ( .A(KEYINPUT24), .B(G119), .ZN(n482) );
  INV_X1 U441 ( .A(KEYINPUT23), .ZN(n484) );
  XNOR2_X1 U442 ( .A(G128), .B(KEYINPUT76), .ZN(n485) );
  XNOR2_X1 U443 ( .A(n781), .B(G146), .ZN(n377) );
  XOR2_X1 U444 ( .A(KEYINPUT106), .B(G122), .Z(n539) );
  INV_X1 U445 ( .A(KEYINPUT64), .ZN(n489) );
  AND2_X1 U446 ( .A1(n368), .A2(KEYINPUT66), .ZN(n361) );
  XNOR2_X1 U447 ( .A(G140), .B(G107), .ZN(n503) );
  XNOR2_X1 U448 ( .A(G104), .B(G101), .ZN(n504) );
  XNOR2_X1 U449 ( .A(n384), .B(n546), .ZN(n383) );
  XNOR2_X1 U450 ( .A(n515), .B(G137), .ZN(n384) );
  NAND2_X1 U451 ( .A1(n386), .A2(n385), .ZN(n592) );
  NAND2_X1 U452 ( .A1(n751), .A2(KEYINPUT34), .ZN(n422) );
  AND2_X1 U453 ( .A1(n445), .A2(n560), .ZN(n444) );
  NOR2_X1 U454 ( .A1(n612), .A2(n611), .ZN(n632) );
  NAND2_X1 U455 ( .A1(n390), .A2(n605), .ZN(n607) );
  AND2_X1 U456 ( .A1(KEYINPUT110), .A2(KEYINPUT67), .ZN(n431) );
  INV_X1 U457 ( .A(KEYINPUT67), .ZN(n426) );
  NOR2_X1 U458 ( .A1(n460), .A2(n641), .ZN(n375) );
  NOR2_X1 U459 ( .A1(n580), .A2(n439), .ZN(n460) );
  INV_X1 U460 ( .A(KEYINPUT103), .ZN(n439) );
  INV_X1 U461 ( .A(KEYINPUT108), .ZN(n406) );
  INV_X1 U462 ( .A(G237), .ZN(n520) );
  XNOR2_X1 U463 ( .A(n476), .B(n477), .ZN(n423) );
  XOR2_X1 U464 ( .A(KEYINPUT5), .B(KEYINPUT81), .Z(n476) );
  NAND2_X1 U465 ( .A1(n397), .A2(KEYINPUT48), .ZN(n396) );
  INV_X1 U466 ( .A(n408), .ZN(n397) );
  XNOR2_X1 U467 ( .A(n782), .B(KEYINPUT82), .ZN(n656) );
  NAND2_X1 U468 ( .A1(n359), .A2(n658), .ZN(n424) );
  AND2_X1 U469 ( .A1(n783), .A2(G224), .ZN(n465) );
  INV_X1 U470 ( .A(KEYINPUT90), .ZN(n459) );
  NAND2_X1 U471 ( .A1(G237), .A2(G234), .ZN(n526) );
  XNOR2_X1 U472 ( .A(n577), .B(n508), .ZN(n563) );
  INV_X1 U473 ( .A(KEYINPUT3), .ZN(n478) );
  XNOR2_X1 U474 ( .A(n555), .B(n554), .ZN(n691) );
  NAND2_X1 U475 ( .A1(n404), .A2(n633), .ZN(n403) );
  AND2_X1 U476 ( .A1(n608), .A2(n632), .ZN(n404) );
  NAND2_X1 U477 ( .A1(n576), .A2(n575), .ZN(n442) );
  INV_X1 U478 ( .A(G953), .ZN(n437) );
  XNOR2_X1 U479 ( .A(n377), .B(n488), .ZN(n492) );
  XNOR2_X1 U480 ( .A(n543), .B(n542), .ZN(n663) );
  NAND2_X1 U481 ( .A1(n362), .A2(n361), .ZN(n360) );
  XNOR2_X1 U482 ( .A(n505), .B(n381), .ZN(n380) );
  INV_X1 U483 ( .A(n452), .ZN(n650) );
  XNOR2_X1 U484 ( .A(KEYINPUT112), .B(KEYINPUT42), .ZN(n450) );
  NAND2_X1 U485 ( .A1(n354), .A2(n421), .ZN(n420) );
  NAND2_X1 U486 ( .A1(n636), .A2(n452), .ZN(n675) );
  AND2_X1 U487 ( .A1(n432), .A2(n430), .ZN(n429) );
  INV_X1 U488 ( .A(n580), .ZN(n707) );
  AND2_X1 U489 ( .A1(n584), .A2(n566), .ZN(n379) );
  AND2_X1 U490 ( .A1(n573), .A2(KEYINPUT44), .ZN(n351) );
  AND2_X1 U491 ( .A1(n468), .A2(n573), .ZN(n352) );
  XOR2_X1 U492 ( .A(G107), .B(G116), .Z(n538) );
  BUF_X1 U493 ( .A(n563), .Z(n725) );
  NAND2_X2 U494 ( .A1(n363), .A2(n360), .ZN(n687) );
  AND2_X1 U495 ( .A1(n427), .A2(n426), .ZN(n353) );
  AND2_X1 U496 ( .A1(n422), .A2(n444), .ZN(n354) );
  NAND2_X1 U497 ( .A1(n398), .A2(n395), .ZN(n782) );
  AND2_X1 U498 ( .A1(n566), .A2(n472), .ZN(n355) );
  AND2_X1 U499 ( .A1(n726), .A2(n610), .ZN(n356) );
  INV_X1 U500 ( .A(G902), .ZN(n415) );
  AND2_X1 U501 ( .A1(n471), .A2(n728), .ZN(n357) );
  INV_X1 U502 ( .A(KEYINPUT48), .ZN(n393) );
  OR2_X1 U503 ( .A1(n661), .A2(KEYINPUT89), .ZN(n358) );
  AND2_X1 U504 ( .A1(n661), .A2(KEYINPUT89), .ZN(n359) );
  INV_X1 U505 ( .A(n367), .ZN(n755) );
  NAND2_X1 U506 ( .A1(n458), .A2(n469), .ZN(n367) );
  NOR2_X1 U507 ( .A1(n369), .A2(n755), .ZN(n362) );
  NAND2_X1 U508 ( .A1(n369), .A2(n662), .ZN(n364) );
  NAND2_X1 U509 ( .A1(n366), .A2(n662), .ZN(n365) );
  NAND2_X1 U510 ( .A1(n367), .A2(n368), .ZN(n366) );
  NAND2_X1 U511 ( .A1(n374), .A2(n372), .ZN(n371) );
  INV_X1 U512 ( .A(n718), .ZN(n373) );
  NAND2_X1 U513 ( .A1(n718), .A2(KEYINPUT103), .ZN(n376) );
  XNOR2_X1 U514 ( .A(n377), .B(n553), .ZN(n554) );
  XNOR2_X1 U515 ( .A(n378), .B(n515), .ZN(n466) );
  XNOR2_X1 U516 ( .A(n382), .B(n378), .ZN(n381) );
  AND2_X1 U517 ( .A1(n569), .A2(n379), .ZN(n704) );
  XNOR2_X2 U518 ( .A(n441), .B(KEYINPUT22), .ZN(n569) );
  NAND2_X1 U519 ( .A1(n783), .A2(G227), .ZN(n382) );
  XNOR2_X2 U520 ( .A(n541), .B(n383), .ZN(n388) );
  XNOR2_X2 U521 ( .A(n453), .B(G143), .ZN(n443) );
  XNOR2_X1 U522 ( .A(n401), .B(n388), .ZN(n678) );
  XNOR2_X1 U523 ( .A(n388), .B(n405), .ZN(n786) );
  NAND2_X1 U524 ( .A1(n389), .A2(n622), .ZN(n512) );
  NAND2_X1 U525 ( .A1(n356), .A2(n728), .ZN(n578) );
  INV_X1 U526 ( .A(n400), .ZN(n394) );
  XNOR2_X1 U527 ( .A(n615), .B(KEYINPUT46), .ZN(n400) );
  NAND2_X1 U528 ( .A1(n400), .A2(n399), .ZN(n391) );
  NAND2_X1 U529 ( .A1(n408), .A2(n393), .ZN(n399) );
  NAND2_X1 U530 ( .A1(n653), .A2(n717), .ZN(n614) );
  INV_X1 U531 ( .A(n781), .ZN(n405) );
  XNOR2_X2 U532 ( .A(n455), .B(n454), .ZN(n576) );
  NAND2_X1 U533 ( .A1(n434), .A2(n357), .ZN(n433) );
  INV_X1 U534 ( .A(n621), .ZN(n717) );
  NAND2_X1 U535 ( .A1(n412), .A2(n622), .ZN(n624) );
  NAND2_X1 U536 ( .A1(n582), .A2(n583), .ZN(n621) );
  NAND2_X1 U537 ( .A1(n700), .A2(n507), .ZN(n419) );
  OR2_X1 U538 ( .A1(n700), .A2(n414), .ZN(n413) );
  INV_X1 U539 ( .A(n507), .ZN(n416) );
  NAND2_X1 U540 ( .A1(n507), .A2(G902), .ZN(n418) );
  OR2_X1 U541 ( .A1(n751), .A2(n446), .ZN(n421) );
  NAND2_X1 U542 ( .A1(n429), .A2(n425), .ZN(n564) );
  NAND2_X1 U543 ( .A1(n428), .A2(n353), .ZN(n425) );
  NAND2_X1 U544 ( .A1(n435), .A2(KEYINPUT110), .ZN(n427) );
  INV_X1 U545 ( .A(n433), .ZN(n428) );
  NAND2_X1 U546 ( .A1(n435), .A2(n431), .ZN(n430) );
  NAND2_X1 U547 ( .A1(n433), .A2(KEYINPUT67), .ZN(n432) );
  NAND2_X1 U548 ( .A1(n569), .A2(n355), .ZN(n434) );
  INV_X1 U549 ( .A(n569), .ZN(n435) );
  NAND2_X1 U550 ( .A1(n469), .A2(n436), .ZN(n470) );
  INV_X1 U551 ( .A(n656), .ZN(n436) );
  AND2_X1 U552 ( .A1(n469), .A2(n659), .ZN(n754) );
  AND2_X1 U553 ( .A1(n469), .A2(n437), .ZN(n778) );
  XNOR2_X2 U554 ( .A(n438), .B(KEYINPUT45), .ZN(n469) );
  NAND2_X1 U555 ( .A1(n592), .A2(n591), .ZN(n438) );
  NAND2_X1 U556 ( .A1(n579), .A2(KEYINPUT34), .ZN(n445) );
  XNOR2_X2 U557 ( .A(n534), .B(n533), .ZN(n579) );
  NAND2_X1 U558 ( .A1(n563), .A2(n726), .ZN(n510) );
  BUF_X1 U559 ( .A(n718), .Z(n440) );
  NOR2_X2 U560 ( .A1(n579), .A2(n562), .ZN(n441) );
  XNOR2_X2 U561 ( .A(n499), .B(n498), .ZN(n601) );
  XNOR2_X1 U562 ( .A(n607), .B(n606), .ZN(n633) );
  XNOR2_X1 U563 ( .A(n660), .B(n459), .ZN(n458) );
  XNOR2_X1 U564 ( .A(n443), .B(n518), .ZN(n463) );
  NAND2_X1 U565 ( .A1(n575), .A2(n447), .ZN(n446) );
  INV_X1 U566 ( .A(KEYINPUT34), .ZN(n447) );
  XNOR2_X2 U567 ( .A(n449), .B(n481), .ZN(n728) );
  NOR2_X1 U568 ( .A1(n750), .A2(n617), .ZN(n451) );
  BUF_X2 U569 ( .A(n593), .Z(n452) );
  XNOR2_X2 U570 ( .A(G128), .B(KEYINPUT65), .ZN(n453) );
  NAND2_X1 U571 ( .A1(n687), .A2(G478), .ZN(n664) );
  NAND2_X1 U572 ( .A1(n687), .A2(G210), .ZN(n767) );
  XNOR2_X1 U573 ( .A(n462), .B(n771), .ZN(n764) );
  XNOR2_X1 U574 ( .A(n464), .B(n463), .ZN(n462) );
  XNOR2_X1 U575 ( .A(n465), .B(n466), .ZN(n464) );
  INV_X1 U576 ( .A(KEYINPUT110), .ZN(n472) );
  OR2_X1 U577 ( .A1(n644), .A2(n643), .ZN(n473) );
  XNOR2_X1 U578 ( .A(n485), .B(n484), .ZN(n486) );
  INV_X1 U579 ( .A(KEYINPUT111), .ZN(n623) );
  INV_X1 U580 ( .A(KEYINPUT30), .ZN(n606) );
  XNOR2_X1 U581 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U582 ( .A(n559), .B(n558), .ZN(n583) );
  INV_X1 U583 ( .A(KEYINPUT40), .ZN(n613) );
  INV_X1 U584 ( .A(KEYINPUT125), .ZN(n668) );
  XNOR2_X1 U585 ( .A(n614), .B(n613), .ZN(n795) );
  XNOR2_X2 U586 ( .A(G146), .B(KEYINPUT4), .ZN(n515) );
  INV_X1 U587 ( .A(KEYINPUT74), .ZN(n474) );
  XNOR2_X1 U588 ( .A(n474), .B(G131), .ZN(n546) );
  XNOR2_X1 U589 ( .A(G116), .B(G113), .ZN(n475) );
  NAND2_X1 U590 ( .A1(n550), .A2(G210), .ZN(n477) );
  INV_X1 U591 ( .A(n513), .ZN(n480) );
  XNOR2_X1 U592 ( .A(G472), .B(KEYINPUT101), .ZN(n481) );
  XOR2_X1 U593 ( .A(G137), .B(G110), .Z(n483) );
  XNOR2_X1 U594 ( .A(n483), .B(n482), .ZN(n487) );
  XNOR2_X2 U595 ( .A(n489), .B(G953), .ZN(n783) );
  NAND2_X1 U596 ( .A1(n783), .A2(G234), .ZN(n490) );
  XOR2_X1 U597 ( .A(KEYINPUT8), .B(n490), .Z(n535) );
  NAND2_X1 U598 ( .A1(G221), .A2(n535), .ZN(n491) );
  XNOR2_X1 U599 ( .A(n492), .B(n491), .ZN(n684) );
  NOR2_X1 U600 ( .A1(n684), .A2(G902), .ZN(n499) );
  XOR2_X1 U601 ( .A(KEYINPUT25), .B(KEYINPUT99), .Z(n495) );
  NAND2_X1 U602 ( .A1(n519), .A2(G234), .ZN(n493) );
  XNOR2_X1 U603 ( .A(n493), .B(KEYINPUT20), .ZN(n500) );
  NAND2_X1 U604 ( .A1(n500), .A2(G217), .ZN(n494) );
  XNOR2_X1 U605 ( .A(n495), .B(n494), .ZN(n497) );
  INV_X1 U606 ( .A(KEYINPUT83), .ZN(n496) );
  XNOR2_X1 U607 ( .A(n497), .B(n496), .ZN(n498) );
  NAND2_X1 U608 ( .A1(G221), .A2(n500), .ZN(n501) );
  XNOR2_X1 U609 ( .A(n501), .B(KEYINPUT21), .ZN(n723) );
  INV_X1 U610 ( .A(KEYINPUT100), .ZN(n502) );
  XNOR2_X1 U611 ( .A(n723), .B(n502), .ZN(n561) );
  AND2_X2 U612 ( .A1(n601), .A2(n561), .ZN(n726) );
  XNOR2_X1 U613 ( .A(n504), .B(n503), .ZN(n505) );
  INV_X1 U614 ( .A(KEYINPUT75), .ZN(n506) );
  XNOR2_X1 U615 ( .A(n506), .B(G469), .ZN(n507) );
  XNOR2_X1 U616 ( .A(KEYINPUT68), .B(KEYINPUT1), .ZN(n508) );
  INV_X1 U617 ( .A(KEYINPUT80), .ZN(n509) );
  XOR2_X1 U618 ( .A(KEYINPUT33), .B(KEYINPUT78), .Z(n511) );
  XNOR2_X1 U619 ( .A(KEYINPUT18), .B(G125), .ZN(n517) );
  XNOR2_X1 U620 ( .A(KEYINPUT93), .B(KEYINPUT17), .ZN(n516) );
  XNOR2_X1 U621 ( .A(n517), .B(n516), .ZN(n518) );
  INV_X1 U622 ( .A(n519), .ZN(n661) );
  OR2_X2 U623 ( .A1(n764), .A2(n661), .ZN(n522) );
  NAND2_X1 U624 ( .A1(n415), .A2(n520), .ZN(n523) );
  AND2_X1 U625 ( .A1(n523), .A2(G210), .ZN(n521) );
  NAND2_X1 U626 ( .A1(n523), .A2(G214), .ZN(n525) );
  INV_X1 U627 ( .A(KEYINPUT95), .ZN(n524) );
  XNOR2_X1 U628 ( .A(n525), .B(n524), .ZN(n605) );
  AND2_X2 U629 ( .A1(n593), .A2(n605), .ZN(n626) );
  XNOR2_X1 U630 ( .A(n626), .B(KEYINPUT19), .ZN(n616) );
  XNOR2_X1 U631 ( .A(n526), .B(KEYINPUT96), .ZN(n527) );
  XNOR2_X1 U632 ( .A(KEYINPUT14), .B(n527), .ZN(n529) );
  NAND2_X1 U633 ( .A1(n529), .A2(G952), .ZN(n528) );
  XOR2_X1 U634 ( .A(KEYINPUT97), .B(n528), .Z(n749) );
  NOR2_X1 U635 ( .A1(n749), .A2(G953), .ZN(n599) );
  NAND2_X1 U636 ( .A1(G902), .A2(n529), .ZN(n597) );
  XOR2_X1 U637 ( .A(G898), .B(KEYINPUT98), .Z(n776) );
  NAND2_X1 U638 ( .A1(G953), .A2(n776), .ZN(n773) );
  NOR2_X1 U639 ( .A1(n597), .A2(n773), .ZN(n530) );
  NOR2_X1 U640 ( .A1(n599), .A2(n530), .ZN(n531) );
  OR2_X2 U641 ( .A1(n616), .A2(n531), .ZN(n534) );
  INV_X1 U642 ( .A(KEYINPUT71), .ZN(n532) );
  XNOR2_X1 U643 ( .A(n532), .B(KEYINPUT0), .ZN(n533) );
  XNOR2_X1 U644 ( .A(G478), .B(KEYINPUT107), .ZN(n545) );
  XOR2_X1 U645 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n537) );
  NAND2_X1 U646 ( .A1(G217), .A2(n535), .ZN(n536) );
  XNOR2_X1 U647 ( .A(n537), .B(n536), .ZN(n543) );
  XNOR2_X1 U648 ( .A(n538), .B(n539), .ZN(n540) );
  XNOR2_X1 U649 ( .A(n541), .B(n540), .ZN(n542) );
  NOR2_X1 U650 ( .A1(n663), .A2(G902), .ZN(n544) );
  XNOR2_X1 U651 ( .A(n545), .B(n544), .ZN(n581) );
  XOR2_X1 U652 ( .A(KEYINPUT104), .B(n546), .Z(n549) );
  XNOR2_X1 U653 ( .A(n547), .B(G143), .ZN(n548) );
  XNOR2_X1 U654 ( .A(n549), .B(n548), .ZN(n555) );
  XOR2_X1 U655 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n552) );
  NAND2_X1 U656 ( .A1(n550), .A2(G214), .ZN(n551) );
  XNOR2_X1 U657 ( .A(n552), .B(n551), .ZN(n553) );
  NOR2_X1 U658 ( .A1(G902), .A2(n691), .ZN(n559) );
  XNOR2_X1 U659 ( .A(KEYINPUT105), .B(KEYINPUT13), .ZN(n557) );
  INV_X1 U660 ( .A(G475), .ZN(n556) );
  NAND2_X1 U661 ( .A1(n581), .A2(n583), .ZN(n635) );
  XOR2_X1 U662 ( .A(KEYINPUT84), .B(n635), .Z(n560) );
  NOR2_X1 U663 ( .A1(n583), .A2(n581), .ZN(n737) );
  NAND2_X1 U664 ( .A1(n737), .A2(n561), .ZN(n562) );
  INV_X1 U665 ( .A(n725), .ZN(n566) );
  INV_X1 U666 ( .A(n601), .ZN(n722) );
  XOR2_X1 U667 ( .A(KEYINPUT85), .B(n565), .Z(n568) );
  NOR2_X1 U668 ( .A1(n566), .A2(n601), .ZN(n567) );
  AND2_X1 U669 ( .A1(n568), .A2(n567), .ZN(n570) );
  NAND2_X1 U670 ( .A1(n570), .A2(n569), .ZN(n572) );
  INV_X1 U671 ( .A(KEYINPUT32), .ZN(n571) );
  XNOR2_X1 U672 ( .A(n572), .B(n571), .ZN(n794) );
  INV_X1 U673 ( .A(n794), .ZN(n573) );
  INV_X1 U674 ( .A(KEYINPUT44), .ZN(n574) );
  INV_X1 U675 ( .A(n579), .ZN(n575) );
  INV_X1 U676 ( .A(n581), .ZN(n582) );
  OR2_X1 U677 ( .A1(n583), .A2(n582), .ZN(n652) );
  NAND2_X1 U678 ( .A1(n621), .A2(n652), .ZN(n740) );
  INV_X1 U679 ( .A(n740), .ZN(n641) );
  NAND2_X1 U680 ( .A1(n792), .A2(KEYINPUT44), .ZN(n586) );
  NOR2_X1 U681 ( .A1(n622), .A2(n722), .ZN(n584) );
  INV_X1 U682 ( .A(n704), .ZN(n585) );
  NAND2_X1 U683 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U684 ( .A1(n588), .A2(n587), .ZN(n590) );
  INV_X1 U685 ( .A(KEYINPUT91), .ZN(n589) );
  XNOR2_X1 U686 ( .A(n590), .B(n589), .ZN(n591) );
  INV_X1 U687 ( .A(KEYINPUT41), .ZN(n595) );
  INV_X1 U688 ( .A(n605), .ZN(n735) );
  NOR2_X1 U689 ( .A1(n736), .A2(n735), .ZN(n739) );
  NAND2_X1 U690 ( .A1(n739), .A2(n737), .ZN(n594) );
  XNOR2_X1 U691 ( .A(n595), .B(n594), .ZN(n750) );
  OR2_X1 U692 ( .A1(n783), .A2(G900), .ZN(n596) );
  NOR2_X1 U693 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U694 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U695 ( .A(KEYINPUT86), .B(n600), .Z(n609) );
  NOR2_X1 U696 ( .A1(n723), .A2(n601), .ZN(n602) );
  NAND2_X1 U697 ( .A1(n609), .A2(n602), .ZN(n620) );
  XNOR2_X1 U698 ( .A(KEYINPUT28), .B(n603), .ZN(n604) );
  NAND2_X1 U699 ( .A1(n604), .A2(n610), .ZN(n617) );
  INV_X1 U700 ( .A(n736), .ZN(n608) );
  NAND2_X1 U701 ( .A1(n726), .A2(n609), .ZN(n612) );
  INV_X1 U702 ( .A(n610), .ZN(n611) );
  NOR2_X1 U703 ( .A1(n617), .A2(n616), .ZN(n714) );
  NAND2_X1 U704 ( .A1(n641), .A2(KEYINPUT88), .ZN(n618) );
  NAND2_X1 U705 ( .A1(n714), .A2(n618), .ZN(n619) );
  NAND2_X1 U706 ( .A1(n619), .A2(KEYINPUT47), .ZN(n631) );
  INV_X1 U707 ( .A(n647), .ZN(n625) );
  NAND2_X1 U708 ( .A1(n626), .A2(n625), .ZN(n629) );
  XOR2_X1 U709 ( .A(KEYINPUT113), .B(KEYINPUT36), .Z(n627) );
  XOR2_X1 U710 ( .A(n627), .B(KEYINPUT92), .Z(n628) );
  XNOR2_X1 U711 ( .A(n629), .B(n628), .ZN(n630) );
  NAND2_X1 U712 ( .A1(n630), .A2(n725), .ZN(n674) );
  NAND2_X1 U713 ( .A1(n631), .A2(n674), .ZN(n645) );
  NAND2_X1 U714 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U715 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U716 ( .A(KEYINPUT47), .B(KEYINPUT72), .Z(n637) );
  NAND2_X1 U717 ( .A1(n637), .A2(n740), .ZN(n638) );
  XNOR2_X1 U718 ( .A(n638), .B(KEYINPUT79), .ZN(n639) );
  NAND2_X1 U719 ( .A1(n714), .A2(n639), .ZN(n640) );
  NAND2_X1 U720 ( .A1(n675), .A2(n640), .ZN(n644) );
  AND2_X1 U721 ( .A1(n641), .A2(KEYINPUT47), .ZN(n642) );
  NOR2_X1 U722 ( .A1(KEYINPUT88), .A2(n642), .ZN(n643) );
  OR2_X1 U723 ( .A1(n725), .A2(n735), .ZN(n646) );
  NOR2_X1 U724 ( .A1(n647), .A2(n646), .ZN(n649) );
  INV_X1 U725 ( .A(KEYINPUT43), .ZN(n648) );
  XNOR2_X1 U726 ( .A(n649), .B(n648), .ZN(n651) );
  NAND2_X1 U727 ( .A1(n651), .A2(n650), .ZN(n672) );
  INV_X1 U728 ( .A(n652), .ZN(n711) );
  AND2_X1 U729 ( .A1(n653), .A2(n711), .ZN(n721) );
  INV_X1 U730 ( .A(n721), .ZN(n654) );
  AND2_X1 U731 ( .A1(n672), .A2(n654), .ZN(n655) );
  INV_X1 U732 ( .A(KEYINPUT89), .ZN(n657) );
  INV_X1 U733 ( .A(KEYINPUT2), .ZN(n658) );
  INV_X1 U734 ( .A(n782), .ZN(n659) );
  NAND2_X1 U735 ( .A1(n659), .A2(KEYINPUT2), .ZN(n660) );
  INV_X1 U736 ( .A(KEYINPUT66), .ZN(n662) );
  XNOR2_X1 U737 ( .A(n664), .B(n663), .ZN(n667) );
  INV_X1 U738 ( .A(n783), .ZN(n666) );
  INV_X1 U739 ( .A(G952), .ZN(n665) );
  NAND2_X1 U740 ( .A1(n666), .A2(n665), .ZN(n694) );
  INV_X1 U741 ( .A(n694), .ZN(n768) );
  XNOR2_X1 U742 ( .A(n669), .B(n668), .ZN(G63) );
  NAND2_X1 U743 ( .A1(n440), .A2(n711), .ZN(n670) );
  XNOR2_X1 U744 ( .A(n670), .B(G116), .ZN(G18) );
  XOR2_X1 U745 ( .A(G140), .B(KEYINPUT119), .Z(n671) );
  XNOR2_X1 U746 ( .A(n672), .B(n671), .ZN(G42) );
  XOR2_X1 U747 ( .A(G125), .B(KEYINPUT37), .Z(n673) );
  XNOR2_X1 U748 ( .A(n674), .B(n673), .ZN(G27) );
  XNOR2_X1 U749 ( .A(n675), .B(G143), .ZN(G45) );
  XNOR2_X1 U750 ( .A(n676), .B(G110), .ZN(G12) );
  NAND2_X1 U751 ( .A1(n687), .A2(G472), .ZN(n680) );
  XOR2_X1 U752 ( .A(KEYINPUT114), .B(KEYINPUT62), .Z(n677) );
  XNOR2_X1 U753 ( .A(n678), .B(n677), .ZN(n679) );
  XNOR2_X1 U754 ( .A(n680), .B(n679), .ZN(n681) );
  NAND2_X1 U755 ( .A1(n681), .A2(n694), .ZN(n683) );
  XOR2_X1 U756 ( .A(KEYINPUT115), .B(KEYINPUT63), .Z(n682) );
  XNOR2_X1 U757 ( .A(n683), .B(n682), .ZN(G57) );
  NAND2_X1 U758 ( .A1(n687), .A2(G217), .ZN(n685) );
  XNOR2_X1 U759 ( .A(n684), .B(n685), .ZN(n686) );
  NOR2_X1 U760 ( .A1(n686), .A2(n768), .ZN(G66) );
  NAND2_X1 U761 ( .A1(n687), .A2(G475), .ZN(n693) );
  XOR2_X1 U762 ( .A(KEYINPUT94), .B(KEYINPUT124), .Z(n689) );
  XNOR2_X1 U763 ( .A(KEYINPUT59), .B(KEYINPUT69), .ZN(n688) );
  XNOR2_X1 U764 ( .A(n689), .B(n688), .ZN(n690) );
  XNOR2_X1 U765 ( .A(n691), .B(n690), .ZN(n692) );
  XNOR2_X1 U766 ( .A(n693), .B(n692), .ZN(n695) );
  NAND2_X1 U767 ( .A1(n695), .A2(n694), .ZN(n697) );
  XOR2_X1 U768 ( .A(KEYINPUT70), .B(KEYINPUT60), .Z(n696) );
  XNOR2_X1 U769 ( .A(n697), .B(n696), .ZN(G60) );
  NAND2_X1 U770 ( .A1(n687), .A2(G469), .ZN(n702) );
  XNOR2_X1 U771 ( .A(KEYINPUT58), .B(KEYINPUT123), .ZN(n698) );
  XNOR2_X1 U772 ( .A(n698), .B(KEYINPUT57), .ZN(n699) );
  XNOR2_X1 U773 ( .A(n700), .B(n699), .ZN(n701) );
  XNOR2_X1 U774 ( .A(n702), .B(n701), .ZN(n703) );
  NOR2_X1 U775 ( .A1(n703), .A2(n768), .ZN(G54) );
  XOR2_X1 U776 ( .A(G101), .B(n704), .Z(G3) );
  NAND2_X1 U777 ( .A1(n707), .A2(n717), .ZN(n705) );
  XNOR2_X1 U778 ( .A(n705), .B(KEYINPUT116), .ZN(n706) );
  XNOR2_X1 U779 ( .A(G104), .B(n706), .ZN(G6) );
  XOR2_X1 U780 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n709) );
  NAND2_X1 U781 ( .A1(n707), .A2(n711), .ZN(n708) );
  XNOR2_X1 U782 ( .A(n709), .B(n708), .ZN(n710) );
  XNOR2_X1 U783 ( .A(G107), .B(n710), .ZN(G9) );
  XOR2_X1 U784 ( .A(G128), .B(KEYINPUT29), .Z(n713) );
  NAND2_X1 U785 ( .A1(n714), .A2(n711), .ZN(n712) );
  XNOR2_X1 U786 ( .A(n713), .B(n712), .ZN(G30) );
  XOR2_X1 U787 ( .A(G146), .B(KEYINPUT117), .Z(n716) );
  NAND2_X1 U788 ( .A1(n714), .A2(n717), .ZN(n715) );
  XNOR2_X1 U789 ( .A(n716), .B(n715), .ZN(G48) );
  NAND2_X1 U790 ( .A1(n440), .A2(n717), .ZN(n719) );
  XNOR2_X1 U791 ( .A(n719), .B(KEYINPUT118), .ZN(n720) );
  XNOR2_X1 U792 ( .A(G113), .B(n720), .ZN(G15) );
  XOR2_X1 U793 ( .A(G134), .B(n721), .Z(G36) );
  XOR2_X1 U794 ( .A(KEYINPUT120), .B(KEYINPUT52), .Z(n747) );
  NAND2_X1 U795 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U796 ( .A(n724), .B(KEYINPUT49), .ZN(n731) );
  NOR2_X1 U797 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U798 ( .A(KEYINPUT50), .B(n727), .Z(n729) );
  NAND2_X1 U799 ( .A1(n729), .A2(n728), .ZN(n730) );
  NOR2_X1 U800 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U801 ( .A1(n732), .A2(n576), .ZN(n733) );
  XOR2_X1 U802 ( .A(KEYINPUT51), .B(n733), .Z(n734) );
  NOR2_X1 U803 ( .A1(n750), .A2(n734), .ZN(n745) );
  NAND2_X1 U804 ( .A1(n736), .A2(n735), .ZN(n738) );
  NAND2_X1 U805 ( .A1(n738), .A2(n737), .ZN(n742) );
  NAND2_X1 U806 ( .A1(n740), .A2(n739), .ZN(n741) );
  AND2_X1 U807 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U808 ( .A1(n751), .A2(n743), .ZN(n744) );
  NOR2_X1 U809 ( .A1(n745), .A2(n744), .ZN(n746) );
  XOR2_X1 U810 ( .A(n747), .B(n746), .Z(n748) );
  NOR2_X1 U811 ( .A1(n749), .A2(n748), .ZN(n753) );
  NOR2_X1 U812 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U813 ( .A1(n753), .A2(n752), .ZN(n758) );
  NOR2_X1 U814 ( .A1(n754), .A2(KEYINPUT2), .ZN(n756) );
  OR2_X1 U815 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U816 ( .A1(n758), .A2(n757), .ZN(n759) );
  XOR2_X1 U817 ( .A(KEYINPUT121), .B(n759), .Z(n760) );
  NOR2_X1 U818 ( .A1(G953), .A2(n760), .ZN(n761) );
  XNOR2_X1 U819 ( .A(KEYINPUT53), .B(n761), .ZN(G75) );
  XOR2_X1 U820 ( .A(KEYINPUT122), .B(KEYINPUT54), .Z(n763) );
  XNOR2_X1 U821 ( .A(KEYINPUT87), .B(KEYINPUT55), .ZN(n762) );
  XNOR2_X1 U822 ( .A(n763), .B(n762), .ZN(n765) );
  XNOR2_X1 U823 ( .A(n767), .B(n766), .ZN(n769) );
  XNOR2_X1 U824 ( .A(n770), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U825 ( .A(n771), .B(G110), .Z(n772) );
  NAND2_X1 U826 ( .A1(n773), .A2(n772), .ZN(n780) );
  NAND2_X1 U827 ( .A1(G953), .A2(G224), .ZN(n774) );
  XOR2_X1 U828 ( .A(KEYINPUT61), .B(n774), .Z(n775) );
  NOR2_X1 U829 ( .A1(n776), .A2(n775), .ZN(n777) );
  NOR2_X1 U830 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U831 ( .A(n780), .B(n779), .ZN(G69) );
  XNOR2_X1 U832 ( .A(n782), .B(n786), .ZN(n784) );
  NAND2_X1 U833 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U834 ( .A(n785), .B(KEYINPUT126), .ZN(n791) );
  XOR2_X1 U835 ( .A(G227), .B(n786), .Z(n787) );
  XNOR2_X1 U836 ( .A(n787), .B(KEYINPUT127), .ZN(n788) );
  NAND2_X1 U837 ( .A1(n788), .A2(G900), .ZN(n789) );
  NAND2_X1 U838 ( .A1(G953), .A2(n789), .ZN(n790) );
  NAND2_X1 U839 ( .A1(n791), .A2(n790), .ZN(G72) );
  XOR2_X1 U840 ( .A(G122), .B(n792), .Z(G24) );
  XOR2_X1 U841 ( .A(G137), .B(n793), .Z(G39) );
  XOR2_X1 U842 ( .A(G119), .B(n794), .Z(G21) );
  XOR2_X1 U843 ( .A(n795), .B(G131), .Z(G33) );
endmodule

