//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1233,
    new_n1234, new_n1235, new_n1236;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  NAND2_X1  g0009(.A1(G107), .A2(G264), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n210), .B1(new_n206), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G50), .A2(G226), .ZN(new_n213));
  INV_X1    g0013(.A(G232), .ZN(new_n214));
  INV_X1    g0014(.A(G116), .ZN(new_n215));
  INV_X1    g0015(.A(G270), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n213), .B1(new_n202), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI211_X1 g0017(.A(new_n212), .B(new_n217), .C1(G87), .C2(G250), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G68), .A2(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  XOR2_X1   g0020(.A(KEYINPUT65), .B(G244), .Z(new_n221));
  OAI211_X1 g0021(.A(new_n218), .B(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G20), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XOR2_X1   g0024(.A(KEYINPUT66), .B(KEYINPUT1), .Z(new_n225));
  XNOR2_X1  g0025(.A(new_n224), .B(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n223), .A2(G13), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT64), .Z(new_n228));
  OAI211_X1 g0028(.A(new_n228), .B(G250), .C1(G257), .C2(G264), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT0), .ZN(new_n230));
  NAND3_X1  g0030(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n231));
  OAI21_X1  g0031(.A(G50), .B1(G58), .B2(G68), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n226), .B(new_n230), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G226), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G264), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n216), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G107), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(new_n215), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G1), .A2(G13), .ZN(new_n252));
  AND2_X1   g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G13), .A3(G20), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(G33), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n253), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  XOR2_X1   g0058(.A(KEYINPUT15), .B(G87), .Z(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n255), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G20), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G97), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT19), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G87), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n267), .A2(new_n206), .A3(new_n207), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n263), .A2(G33), .A3(G97), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n266), .A2(new_n268), .B1(new_n265), .B2(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT3), .B(G33), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(new_n263), .A3(G68), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n260), .B(new_n262), .C1(new_n273), .C2(new_n253), .ZN(new_n274));
  INV_X1    g0074(.A(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT3), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT3), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G33), .ZN(new_n278));
  INV_X1    g0078(.A(G1698), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n276), .A2(new_n278), .A3(G238), .A4(new_n279), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n276), .A2(new_n278), .A3(G244), .A4(G1698), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G116), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G33), .A2(G41), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n284), .A2(G1), .A3(G13), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G179), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n254), .A2(G45), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n285), .A2(G250), .A3(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n289), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G274), .ZN(new_n292));
  AOI21_X1  g0092(.A(KEYINPUT82), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  AND3_X1   g0093(.A1(new_n290), .A2(new_n292), .A3(KEYINPUT82), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n287), .B(new_n288), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n290), .A2(new_n292), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT82), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n290), .A2(new_n292), .A3(KEYINPUT82), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n298), .A2(new_n299), .B1(new_n286), .B2(new_n283), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n274), .B(new_n295), .C1(new_n300), .C2(G169), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n253), .B1(new_n270), .B2(new_n272), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n257), .A2(new_n267), .ZN(new_n303));
  NOR3_X1   g0103(.A1(new_n302), .A2(new_n303), .A3(new_n261), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n287), .B(G190), .C1(new_n293), .C2(new_n294), .ZN(new_n305));
  INV_X1    g0105(.A(G200), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n304), .B(new_n305), .C1(new_n300), .C2(new_n306), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n301), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n255), .A2(G97), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n257), .A2(new_n206), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n276), .A2(new_n278), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT7), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n311), .A2(new_n312), .A3(new_n263), .ZN(new_n313));
  AOI21_X1  g0113(.A(G20), .B1(new_n276), .B2(new_n278), .ZN(new_n314));
  AND2_X1   g0114(.A1(KEYINPUT74), .A2(KEYINPUT7), .ZN(new_n315));
  NOR2_X1   g0115(.A1(KEYINPUT74), .A2(KEYINPUT7), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n313), .B(G107), .C1(new_n314), .C2(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(G20), .A2(G33), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G77), .ZN(new_n321));
  NAND2_X1  g0121(.A1(G97), .A2(G107), .ZN(new_n322));
  AOI21_X1  g0122(.A(KEYINPUT6), .B1(new_n208), .B2(new_n322), .ZN(new_n323));
  AND3_X1   g0123(.A1(new_n207), .A2(KEYINPUT6), .A3(G97), .ZN(new_n324));
  OAI21_X1  g0124(.A(G20), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n319), .A2(new_n321), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n251), .A2(new_n252), .ZN(new_n327));
  AOI211_X1 g0127(.A(new_n309), .B(new_n310), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n276), .A2(new_n278), .A3(G244), .A4(new_n279), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT4), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n271), .A2(KEYINPUT4), .A3(G244), .A4(new_n279), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n271), .A2(G250), .A3(G1698), .ZN(new_n333));
  NAND2_X1  g0133(.A1(G33), .A2(G283), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n331), .A2(new_n332), .A3(new_n333), .A4(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n286), .ZN(new_n336));
  XNOR2_X1  g0136(.A(KEYINPUT5), .B(G41), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n291), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n338), .A2(G257), .A3(new_n285), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT81), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n337), .A2(G274), .A3(new_n291), .ZN(new_n341));
  AND3_X1   g0141(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n340), .B1(new_n339), .B2(new_n341), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n336), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G200), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n336), .B(G190), .C1(new_n342), .C2(new_n343), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n328), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G169), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n326), .A2(new_n327), .ZN(new_n350));
  INV_X1    g0150(.A(new_n309), .ZN(new_n351));
  INV_X1    g0151(.A(new_n310), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n336), .B(new_n288), .C1(new_n342), .C2(new_n343), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n349), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  AND3_X1   g0155(.A1(new_n308), .A2(new_n347), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT8), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(G58), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n360), .A2(new_n263), .A3(G33), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n320), .A2(G150), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT69), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n204), .A2(new_n363), .A3(G20), .ZN(new_n364));
  NOR3_X1   g0164(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT69), .B1(new_n365), .B2(new_n263), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n361), .A2(new_n362), .A3(new_n364), .A4(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n255), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n367), .A2(new_n327), .B1(new_n201), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT70), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(new_n263), .B2(G1), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n253), .A2(new_n255), .A3(new_n371), .ZN(new_n372));
  NOR3_X1   g0172(.A1(new_n370), .A2(new_n263), .A3(G1), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(G50), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n369), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(KEYINPUT71), .A2(KEYINPUT9), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT71), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT9), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n376), .A2(new_n377), .A3(new_n380), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n369), .A2(new_n378), .A3(new_n379), .A4(new_n375), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n254), .B1(G41), .B2(G45), .ZN(new_n384));
  INV_X1    g0184(.A(G274), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n271), .A2(G223), .A3(G1698), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n271), .A2(G222), .A3(new_n279), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n387), .B(new_n388), .C1(new_n220), .C2(new_n271), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n386), .B1(new_n389), .B2(new_n286), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n285), .A2(new_n384), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  OR2_X1    g0192(.A1(KEYINPUT68), .A2(G226), .ZN(new_n393));
  NAND2_X1  g0193(.A1(KEYINPUT68), .A2(G226), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(G200), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n389), .A2(new_n286), .ZN(new_n398));
  INV_X1    g0198(.A(new_n386), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n398), .A2(G190), .A3(new_n399), .A4(new_n395), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT72), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n390), .A2(KEYINPUT72), .A3(G190), .A4(new_n395), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n383), .A2(new_n397), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT10), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n383), .A2(new_n404), .A3(KEYINPUT10), .A4(new_n397), .ZN(new_n408));
  AND2_X1   g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n271), .A2(G226), .A3(new_n279), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n271), .A2(G232), .A3(G1698), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(new_n411), .A3(new_n264), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n386), .B1(new_n412), .B2(new_n286), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT13), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n392), .A2(G238), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n414), .B1(new_n413), .B2(new_n415), .ZN(new_n417));
  OAI21_X1  g0217(.A(G200), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n263), .A2(G33), .A3(G77), .ZN(new_n419));
  INV_X1    g0219(.A(new_n320), .ZN(new_n420));
  OAI221_X1 g0220(.A(new_n419), .B1(new_n263), .B2(G68), .C1(new_n420), .C2(new_n201), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n327), .ZN(new_n422));
  XNOR2_X1  g0222(.A(new_n422), .B(KEYINPUT11), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n374), .A2(G68), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n368), .A2(new_n203), .ZN(new_n425));
  XNOR2_X1  g0225(.A(new_n425), .B(KEYINPUT12), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n423), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n412), .A2(new_n286), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n429), .A2(new_n415), .A3(new_n399), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT13), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n431), .A2(G190), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n418), .A2(new_n428), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT73), .ZN(new_n435));
  XNOR2_X1  g0235(.A(new_n434), .B(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n396), .A2(new_n348), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n437), .B(new_n376), .C1(G179), .C2(new_n396), .ZN(new_n438));
  INV_X1    g0238(.A(new_n259), .ZN(new_n439));
  NOR3_X1   g0239(.A1(new_n439), .A2(G20), .A3(new_n275), .ZN(new_n440));
  INV_X1    g0240(.A(new_n360), .ZN(new_n441));
  OAI22_X1  g0241(.A1(new_n441), .A2(new_n420), .B1(new_n263), .B2(new_n220), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n327), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n368), .A2(new_n220), .ZN(new_n444));
  INV_X1    g0244(.A(new_n373), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n253), .A2(new_n255), .A3(new_n445), .A4(new_n371), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n443), .B(new_n444), .C1(new_n220), .C2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n271), .A2(G238), .A3(G1698), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n448), .B1(new_n207), .B2(new_n271), .ZN(new_n449));
  NOR3_X1   g0249(.A1(new_n311), .A2(new_n214), .A3(G1698), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n286), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OR2_X1    g0251(.A1(new_n391), .A2(new_n221), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n451), .A2(new_n399), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n447), .B1(G200), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(G190), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n454), .B1(new_n455), .B2(new_n453), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n409), .A2(new_n436), .A3(new_n438), .A4(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n447), .B1(new_n453), .B2(G179), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n453), .A2(new_n348), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(G169), .B1(new_n416), .B2(new_n417), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT14), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT14), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n463), .B(G169), .C1(new_n416), .C2(new_n417), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n431), .A2(G179), .A3(new_n432), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n462), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n460), .B1(new_n466), .B2(new_n427), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT75), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n314), .A2(new_n468), .A3(new_n317), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT75), .B1(new_n314), .B2(KEYINPUT7), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n311), .A2(new_n317), .A3(new_n263), .ZN(new_n471));
  OAI211_X1 g0271(.A(G68), .B(new_n469), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT76), .ZN(new_n473));
  INV_X1    g0273(.A(G159), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n473), .B1(new_n420), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n320), .A2(KEYINPUT76), .A3(G159), .ZN(new_n476));
  XNOR2_X1  g0276(.A(G58), .B(G68), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n475), .A2(new_n476), .B1(new_n477), .B2(G20), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n472), .A2(KEYINPUT16), .A3(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n313), .B(G68), .C1(new_n314), .C2(new_n318), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n478), .ZN(new_n481));
  XNOR2_X1  g0281(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n479), .A2(new_n327), .A3(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n276), .A2(new_n278), .A3(G226), .A4(G1698), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n276), .A2(new_n278), .A3(G223), .A4(new_n279), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G33), .A2(G87), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n386), .B1(new_n488), .B2(new_n286), .ZN(new_n489));
  OAI21_X1  g0289(.A(KEYINPUT79), .B1(new_n391), .B2(new_n214), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT79), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n285), .A2(new_n384), .A3(new_n491), .A4(G232), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n306), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n489), .A2(new_n455), .A3(new_n493), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n360), .A2(new_n368), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(new_n374), .B2(new_n441), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT78), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n498), .B1(new_n446), .B2(new_n360), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT78), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n484), .A2(new_n497), .A3(new_n505), .ZN(new_n506));
  XNOR2_X1  g0306(.A(new_n506), .B(KEYINPUT17), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n484), .A2(new_n505), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n494), .A2(G169), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n489), .A2(G179), .A3(new_n493), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(KEYINPUT18), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT80), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n508), .A2(KEYINPUT18), .A3(new_n511), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI211_X1 g0315(.A(KEYINPUT80), .B(KEYINPUT18), .C1(new_n508), .C2(new_n511), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n467), .B(new_n507), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n457), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n276), .A2(new_n278), .A3(new_n263), .A4(G87), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT22), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT22), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n271), .A2(new_n521), .A3(new_n263), .A4(G87), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n282), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n263), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n263), .A2(G107), .ZN(new_n526));
  XNOR2_X1  g0326(.A(new_n526), .B(KEYINPUT23), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT24), .ZN(new_n528));
  OR2_X1    g0328(.A1(new_n528), .A2(KEYINPUT84), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n523), .A2(new_n525), .A3(new_n527), .A4(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n530), .A2(KEYINPUT84), .A3(new_n528), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n520), .A2(new_n522), .B1(new_n263), .B2(new_n524), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n528), .A2(KEYINPUT84), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n532), .A2(new_n527), .A3(new_n529), .A4(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n531), .A2(new_n327), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n258), .A2(G107), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n255), .A2(G107), .ZN(new_n537));
  XNOR2_X1  g0337(.A(new_n537), .B(KEYINPUT25), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n535), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n271), .A2(G257), .A3(G1698), .ZN(new_n540));
  NAND2_X1  g0340(.A1(G33), .A2(G294), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n276), .A2(new_n278), .A3(G250), .A4(new_n279), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n286), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n286), .B1(new_n291), .B2(new_n337), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G264), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n341), .A3(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT85), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n341), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n550), .B1(new_n543), .B2(new_n286), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n551), .A2(KEYINPUT85), .A3(new_n546), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n549), .A2(new_n455), .A3(new_n552), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n544), .A2(new_n341), .A3(new_n546), .ZN(new_n554));
  OAI21_X1  g0354(.A(KEYINPUT86), .B1(new_n554), .B2(G200), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT86), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n547), .A2(new_n556), .A3(new_n306), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n553), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n539), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n535), .A2(new_n536), .A3(new_n538), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n348), .B1(new_n549), .B2(new_n552), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n547), .A2(new_n288), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n251), .A2(new_n252), .B1(G20), .B2(new_n215), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n334), .B(new_n263), .C1(G33), .C2(new_n206), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(KEYINPUT20), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT83), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n565), .A2(new_n566), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT20), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT83), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n565), .A2(new_n572), .A3(new_n566), .A4(KEYINPUT20), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n568), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n258), .A2(G116), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n368), .A2(new_n215), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n271), .A2(G257), .A3(new_n279), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n271), .A2(G264), .A3(G1698), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n311), .A2(G303), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n286), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n545), .A2(G270), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n341), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n577), .A2(new_n584), .A3(G169), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(KEYINPUT21), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT21), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n577), .A2(new_n584), .A3(new_n587), .A4(G169), .ZN(new_n588));
  INV_X1    g0388(.A(new_n577), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n589), .A2(new_n584), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n586), .A2(new_n588), .B1(new_n590), .B2(G179), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n584), .A2(G200), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n592), .B(new_n589), .C1(new_n455), .C2(new_n584), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  AND4_X1   g0394(.A1(new_n356), .A2(new_n518), .A3(new_n564), .A4(new_n594), .ZN(G372));
  NAND2_X1  g0395(.A1(new_n508), .A2(new_n511), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT18), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n598), .A2(new_n514), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n418), .A2(new_n428), .A3(new_n433), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n507), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n600), .B1(new_n602), .B2(new_n467), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT87), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n600), .B(KEYINPUT87), .C1(new_n602), .C2(new_n467), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(new_n409), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n563), .A2(new_n591), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n608), .A2(new_n356), .A3(new_n559), .ZN(new_n609));
  INV_X1    g0409(.A(new_n301), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n353), .A2(new_n354), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n308), .A2(new_n611), .A3(KEYINPUT26), .A4(new_n349), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT26), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n301), .A2(new_n307), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n613), .B1(new_n355), .B2(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n610), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n609), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n518), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n607), .A2(new_n618), .A3(new_n438), .ZN(G369));
  INV_X1    g0419(.A(new_n591), .ZN(new_n620));
  INV_X1    g0420(.A(G13), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n621), .A2(G20), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n254), .ZN(new_n623));
  OR2_X1    g0423(.A1(new_n623), .A2(KEYINPUT27), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(KEYINPUT27), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n624), .A2(G213), .A3(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(G343), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n564), .A2(new_n620), .A3(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n564), .B1(new_n539), .B2(new_n629), .ZN(new_n631));
  OR2_X1    g0431(.A1(new_n563), .A2(new_n629), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n591), .A2(new_n628), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n630), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n589), .A2(new_n629), .ZN(new_n637));
  MUX2_X1   g0437(.A(new_n594), .B(new_n620), .S(new_n637), .Z(new_n638));
  AND2_X1   g0438(.A1(new_n638), .A2(G330), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n608), .A2(new_n559), .A3(new_n629), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(G399));
  INV_X1    g0444(.A(KEYINPUT89), .ZN(new_n645));
  INV_X1    g0445(.A(new_n228), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT88), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n646), .A2(new_n647), .A3(G41), .ZN(new_n648));
  INV_X1    g0448(.A(G41), .ZN(new_n649));
  AOI21_X1  g0449(.A(KEYINPUT88), .B1(new_n228), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n645), .B1(new_n652), .B2(new_n232), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n651), .A2(new_n254), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n268), .A2(G116), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(KEYINPUT89), .B2(new_n656), .ZN(new_n658));
  XNOR2_X1  g0458(.A(new_n658), .B(KEYINPUT28), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT30), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n339), .A2(new_n341), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(KEYINPUT81), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n662), .A2(new_n663), .B1(new_n286), .B2(new_n335), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n582), .A2(new_n583), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n554), .A2(G179), .A3(new_n300), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n660), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  AND4_X1   g0468(.A1(G179), .A2(new_n300), .A3(new_n546), .A4(new_n551), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n669), .A2(KEYINPUT30), .A3(new_n664), .A4(new_n665), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n344), .A2(new_n547), .A3(new_n584), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n672), .A2(G179), .A3(new_n300), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(new_n629), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n564), .A2(new_n356), .A3(new_n594), .A4(new_n629), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n675), .B1(new_n676), .B2(KEYINPUT31), .ZN(new_n677));
  OAI211_X1 g0477(.A(KEYINPUT31), .B(new_n628), .C1(new_n671), .C2(new_n673), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT90), .ZN(new_n679));
  OAI21_X1  g0479(.A(G330), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n617), .A2(new_n629), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT29), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n628), .B1(new_n609), .B2(new_n616), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(KEYINPUT29), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n680), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n659), .B1(new_n688), .B2(G1), .ZN(G364));
  NOR2_X1   g0489(.A1(new_n263), .A2(G179), .ZN(new_n690));
  NOR2_X1   g0490(.A1(G190), .A2(G200), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n693), .A2(G329), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n263), .A2(new_n288), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G200), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(new_n455), .ZN(new_n697));
  AOI211_X1 g0497(.A(new_n271), .B(new_n694), .C1(G326), .C2(new_n697), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n695), .A2(KEYINPUT93), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n455), .A2(G200), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n695), .A2(KEYINPUT93), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  AND3_X1   g0503(.A1(new_n699), .A2(new_n701), .A3(new_n691), .ZN(new_n704));
  AOI22_X1  g0504(.A1(G322), .A2(new_n703), .B1(new_n704), .B2(G311), .ZN(new_n705));
  INV_X1    g0505(.A(G283), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n690), .A2(new_n455), .A3(G200), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n690), .A2(G190), .A3(G200), .ZN(new_n708));
  INV_X1    g0508(.A(G303), .ZN(new_n709));
  OAI22_X1  g0509(.A1(new_n706), .A2(new_n707), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n696), .A2(G190), .ZN(new_n711));
  XNOR2_X1  g0511(.A(KEYINPUT33), .B(G317), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n700), .A2(new_n288), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G20), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(G294), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n698), .A2(new_n705), .A3(new_n713), .A4(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n708), .A2(new_n267), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n693), .A2(G159), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT32), .ZN(new_n720));
  AOI211_X1 g0520(.A(new_n718), .B(new_n720), .C1(G68), .C2(new_n711), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n707), .A2(new_n207), .ZN(new_n722));
  AOI211_X1 g0522(.A(new_n311), .B(new_n722), .C1(G50), .C2(new_n697), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  XOR2_X1   g0524(.A(new_n702), .B(KEYINPUT94), .Z(new_n725));
  INV_X1    g0525(.A(new_n704), .ZN(new_n726));
  OAI221_X1 g0526(.A(new_n724), .B1(new_n202), .B2(new_n725), .C1(new_n220), .C2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n715), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(new_n206), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n717), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n252), .B1(G20), .B2(new_n348), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n228), .A2(new_n311), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n732), .B(KEYINPUT91), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n734), .B1(new_n246), .B2(G45), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n735), .B1(G45), .B2(new_n232), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n228), .A2(new_n271), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G355), .ZN(new_n739));
  OAI211_X1 g0539(.A(new_n736), .B(new_n739), .C1(G116), .C2(new_n228), .ZN(new_n740));
  NOR2_X1   g0540(.A1(G13), .A2(G33), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(new_n263), .ZN(new_n742));
  XOR2_X1   g0542(.A(new_n742), .B(KEYINPUT92), .Z(new_n743));
  INV_X1    g0543(.A(new_n731), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AOI22_X1  g0545(.A1(new_n730), .A2(new_n731), .B1(new_n740), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n622), .A2(G45), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n654), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n746), .B(new_n749), .C1(new_n638), .C2(new_n743), .ZN(new_n750));
  XOR2_X1   g0550(.A(new_n750), .B(KEYINPUT95), .Z(new_n751));
  NOR2_X1   g0551(.A1(new_n639), .A2(new_n749), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(G330), .B2(new_n638), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n751), .A2(new_n753), .ZN(G396));
  NAND2_X1  g0554(.A1(new_n447), .A2(new_n628), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n460), .B1(new_n456), .B2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n460), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n628), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n681), .B(new_n759), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(new_n680), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n748), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n267), .A2(new_n707), .B1(new_n708), .B2(new_n207), .ZN(new_n763));
  INV_X1    g0563(.A(G311), .ZN(new_n764));
  OAI221_X1 g0564(.A(new_n311), .B1(new_n692), .B2(new_n764), .C1(new_n728), .C2(new_n206), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n763), .B(new_n765), .C1(G283), .C2(new_n711), .ZN(new_n766));
  AOI22_X1  g0566(.A1(G294), .A2(new_n703), .B1(new_n704), .B2(G116), .ZN(new_n767));
  INV_X1    g0567(.A(new_n697), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n766), .B(new_n767), .C1(new_n709), .C2(new_n768), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT96), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n704), .A2(G159), .B1(G137), .B2(new_n697), .ZN(new_n771));
  INV_X1    g0571(.A(G150), .ZN(new_n772));
  INV_X1    g0572(.A(new_n711), .ZN(new_n773));
  INV_X1    g0573(.A(G143), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n771), .B1(new_n772), .B2(new_n773), .C1(new_n725), .C2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT34), .ZN(new_n776));
  OR2_X1    g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n693), .A2(G132), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n775), .A2(new_n776), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n728), .A2(new_n202), .B1(new_n707), .B2(new_n203), .ZN(new_n780));
  INV_X1    g0580(.A(new_n708), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n311), .B(new_n780), .C1(G50), .C2(new_n781), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n777), .A2(new_n778), .A3(new_n779), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n770), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n748), .B1(new_n784), .B2(new_n731), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n731), .A2(new_n741), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n741), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n785), .B1(G77), .B2(new_n787), .C1(new_n788), .C2(new_n759), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n762), .A2(new_n789), .ZN(G384));
  INV_X1    g0590(.A(KEYINPUT101), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n678), .B(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n677), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n428), .A2(new_n629), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n434), .B(KEYINPUT73), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n794), .B1(new_n795), .B2(new_n466), .ZN(new_n796));
  INV_X1    g0596(.A(new_n794), .ZN(new_n797));
  INV_X1    g0597(.A(new_n466), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n434), .B(new_n797), .C1(new_n798), .C2(new_n428), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR4_X1   g0601(.A1(new_n793), .A2(new_n801), .A3(new_n758), .A4(new_n756), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n509), .A2(new_n510), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n803), .A2(new_n626), .B1(new_n484), .B2(new_n505), .ZN(new_n804));
  AND3_X1   g0604(.A1(new_n484), .A2(new_n497), .A3(new_n505), .ZN(new_n805));
  OAI21_X1  g0605(.A(KEYINPUT37), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(KEYINPUT98), .ZN(new_n807));
  AND3_X1   g0607(.A1(new_n479), .A2(new_n327), .A3(new_n483), .ZN(new_n808));
  INV_X1    g0608(.A(new_n505), .ZN(new_n809));
  INV_X1    g0609(.A(new_n626), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n808), .A2(new_n809), .B1(new_n511), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT37), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n811), .A2(new_n812), .A3(new_n506), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(KEYINPUT99), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT98), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n815), .B(KEYINPUT37), .C1(new_n804), .C2(new_n805), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT99), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n811), .A2(new_n817), .A3(new_n812), .A4(new_n506), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n807), .A2(new_n814), .A3(new_n816), .A4(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n626), .B1(new_n484), .B2(new_n505), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT17), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n506), .B(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n820), .B1(new_n599), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT38), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n472), .A2(new_n478), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(KEYINPUT97), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT97), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n472), .A2(new_n829), .A3(new_n478), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n828), .A2(new_n482), .A3(new_n830), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n479), .A2(new_n327), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n833), .A2(new_n500), .B1(new_n803), .B2(new_n626), .ZN(new_n834));
  OAI21_X1  g0634(.A(KEYINPUT37), .B1(new_n834), .B2(new_n805), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(new_n813), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n514), .A2(new_n513), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n598), .ZN(new_n838));
  INV_X1    g0638(.A(new_n516), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n822), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n502), .B1(new_n831), .B2(new_n832), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n841), .A2(new_n626), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n836), .B(KEYINPUT38), .C1(new_n840), .C2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n826), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n802), .A2(KEYINPUT40), .A3(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n836), .B1(new_n840), .B2(new_n843), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(new_n825), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n844), .ZN(new_n850));
  AOI21_X1  g0650(.A(KEYINPUT40), .B1(new_n802), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  OR2_X1    g0652(.A1(new_n677), .A2(new_n792), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n518), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n852), .B(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(G330), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n683), .A2(new_n518), .A3(new_n685), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n857), .A2(new_n438), .A3(new_n607), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n856), .B(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT100), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n466), .A2(new_n427), .A3(new_n629), .ZN(new_n861));
  INV_X1    g0661(.A(new_n844), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n507), .B1(new_n515), .B2(new_n516), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n842), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT38), .B1(new_n864), .B2(new_n836), .ZN(new_n865));
  OAI21_X1  g0665(.A(KEYINPUT39), .B1(new_n862), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT39), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n826), .A2(new_n867), .A3(new_n844), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n861), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n862), .A2(new_n865), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n617), .A2(new_n629), .A3(new_n759), .ZN(new_n871));
  INV_X1    g0671(.A(new_n758), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n800), .ZN(new_n874));
  OAI22_X1  g0674(.A1(new_n870), .A2(new_n874), .B1(new_n600), .B2(new_n810), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n860), .B1(new_n869), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n861), .ZN(new_n877));
  AND3_X1   g0677(.A1(new_n826), .A2(new_n867), .A3(new_n844), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n867), .B1(new_n849), .B2(new_n844), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n758), .B1(new_n684), .B2(new_n759), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n801), .A2(new_n881), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n882), .A2(new_n850), .B1(new_n599), .B2(new_n626), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n880), .A2(new_n883), .A3(KEYINPUT100), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n876), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n859), .B(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n254), .B2(new_n622), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n323), .A2(new_n324), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT35), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n231), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n890), .B(G116), .C1(new_n889), .C2(new_n888), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n891), .B(KEYINPUT36), .ZN(new_n892));
  OAI21_X1  g0692(.A(G77), .B1(new_n202), .B2(new_n203), .ZN(new_n893));
  OAI22_X1  g0693(.A1(new_n893), .A2(new_n232), .B1(G50), .B2(new_n203), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n894), .A2(G1), .A3(new_n621), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n887), .A2(new_n892), .A3(new_n895), .ZN(G367));
  OAI221_X1 g0696(.A(new_n745), .B1(new_n228), .B2(new_n439), .C1(new_n734), .C2(new_n242), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n749), .A2(new_n897), .ZN(new_n898));
  XOR2_X1   g0698(.A(new_n898), .B(KEYINPUT106), .Z(new_n899));
  NOR2_X1   g0699(.A1(new_n629), .A2(new_n304), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n610), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n614), .B2(new_n900), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n708), .A2(new_n202), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n728), .A2(new_n203), .ZN(new_n904));
  AOI211_X1 g0704(.A(new_n903), .B(new_n904), .C1(G159), .C2(new_n711), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n697), .A2(G143), .ZN(new_n906));
  AOI22_X1  g0706(.A1(G150), .A2(new_n703), .B1(new_n704), .B2(G50), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n271), .B1(new_n707), .B2(new_n220), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(G137), .B2(new_n693), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n905), .A2(new_n906), .A3(new_n907), .A4(new_n909), .ZN(new_n910));
  OR2_X1    g0710(.A1(new_n725), .A2(new_n709), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n781), .A2(G116), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT46), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI211_X1 g0714(.A(new_n271), .B(new_n914), .C1(G317), .C2(new_n693), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n707), .A2(new_n206), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n912), .B2(new_n913), .ZN(new_n917));
  INV_X1    g0717(.A(G294), .ZN(new_n918));
  OAI22_X1  g0718(.A1(new_n773), .A2(new_n918), .B1(new_n728), .B2(new_n207), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(G283), .B2(new_n704), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n911), .A2(new_n915), .A3(new_n917), .A4(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n768), .A2(new_n764), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n910), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n923), .B(KEYINPUT47), .Z(new_n924));
  OAI221_X1 g0724(.A(new_n899), .B1(new_n743), .B2(new_n902), .C1(new_n924), .C2(new_n744), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n651), .B(KEYINPUT41), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n636), .B(new_n640), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n928), .A2(new_n687), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n347), .A2(new_n355), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n643), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT44), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n932), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n933), .A2(KEYINPUT104), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n930), .B1(new_n328), .B2(new_n629), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n611), .A2(new_n349), .A3(new_n628), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n643), .ZN(new_n939));
  XNOR2_X1  g0739(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n939), .B(new_n940), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n935), .B(new_n941), .C1(KEYINPUT104), .C2(new_n934), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n929), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n927), .B1(new_n943), .B2(new_n688), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT105), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n747), .A2(G1), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n641), .A2(new_n938), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n938), .A2(new_n564), .A3(new_n635), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT42), .Z(new_n949));
  OAI21_X1  g0749(.A(new_n355), .B1(new_n936), .B2(new_n563), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n629), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n949), .A2(new_n951), .B1(KEYINPUT43), .B2(new_n902), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n902), .A2(KEYINPUT43), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n952), .B(new_n953), .Z(new_n954));
  OAI22_X1  g0754(.A1(new_n945), .A2(new_n946), .B1(new_n947), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n947), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT102), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n925), .B1(new_n955), .B2(new_n957), .ZN(G387));
  INV_X1    g0758(.A(new_n743), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n734), .B1(new_n239), .B2(G45), .ZN(new_n960));
  INV_X1    g0760(.A(new_n655), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n960), .B1(new_n961), .B2(new_n738), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n360), .A2(new_n201), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT107), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT50), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n655), .B1(new_n203), .B2(new_n220), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  AOI211_X1 g0766(.A(G45), .B(new_n966), .C1(new_n965), .C2(new_n964), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n962), .A2(new_n967), .B1(G107), .B2(new_n228), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n633), .A2(new_n959), .B1(new_n745), .B2(new_n968), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n704), .A2(G303), .B1(G322), .B2(new_n697), .ZN(new_n970));
  INV_X1    g0770(.A(G317), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n970), .B1(new_n764), .B2(new_n773), .C1(new_n725), .C2(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT48), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n973), .B1(new_n706), .B2(new_n728), .C1(new_n918), .C2(new_n708), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n974), .A2(KEYINPUT108), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(KEYINPUT108), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT49), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n693), .A2(G326), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n975), .A2(KEYINPUT49), .A3(new_n976), .ZN(new_n981));
  INV_X1    g0781(.A(new_n707), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n271), .B1(new_n982), .B2(G116), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n979), .A2(new_n980), .A3(new_n981), .A4(new_n983), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n768), .A2(new_n474), .B1(new_n708), .B2(new_n220), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(new_n360), .B2(new_n711), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n715), .A2(new_n259), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G50), .A2(new_n703), .B1(new_n704), .B2(G68), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n311), .B(new_n916), .C1(G150), .C2(new_n693), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n986), .A2(new_n987), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n984), .A2(new_n990), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n749), .B(new_n969), .C1(new_n991), .C2(new_n744), .ZN(new_n992));
  INV_X1    g0792(.A(new_n946), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n928), .A2(new_n687), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n651), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n992), .B1(new_n993), .B2(new_n928), .C1(new_n929), .C2(new_n995), .ZN(G393));
  XNOR2_X1  g0796(.A(new_n642), .B(new_n942), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n943), .B(new_n651), .C1(new_n997), .C2(new_n929), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n946), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n704), .A2(G294), .B1(G303), .B2(new_n711), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n215), .B2(new_n728), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT109), .Z(new_n1002));
  AOI21_X1  g0802(.A(new_n271), .B1(new_n693), .B2(G322), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n764), .A2(new_n702), .B1(new_n768), .B2(new_n971), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT52), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n722), .B1(G283), .B2(new_n781), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n715), .A2(G77), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n203), .B2(new_n708), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n271), .B1(new_n692), .B2(new_n774), .C1(new_n267), .C2(new_n707), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n441), .B2(new_n726), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT51), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n474), .A2(new_n702), .B1(new_n768), .B2(new_n772), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1012), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1015), .B1(new_n1013), .B2(new_n1014), .C1(new_n201), .C2(new_n773), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1007), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n748), .B1(new_n1017), .B2(new_n731), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n745), .B1(new_n206), .B2(new_n228), .C1(new_n734), .C2(new_n249), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1018), .B(new_n1019), .C1(new_n743), .C2(new_n938), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n998), .A2(new_n999), .A3(new_n1020), .ZN(G390));
  INV_X1    g0821(.A(G330), .ZN(new_n1022));
  NOR3_X1   g0822(.A1(new_n756), .A2(new_n758), .A3(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n677), .B2(new_n679), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1024), .A2(new_n801), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT110), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1023), .B1(new_n677), .B2(new_n792), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1025), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n877), .B1(new_n873), .B2(new_n800), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(new_n866), .B2(new_n868), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n861), .B1(new_n801), .B2(new_n881), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1031), .A2(new_n845), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1028), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1031), .B1(new_n878), .B2(new_n879), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1029), .A2(new_n844), .A3(new_n826), .ZN(new_n1035));
  NOR3_X1   g0835(.A1(new_n1027), .A2(KEYINPUT110), .A3(new_n801), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1033), .A2(new_n1037), .A3(new_n946), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n866), .A2(new_n741), .A3(new_n868), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n704), .A2(G97), .B1(G283), .B2(new_n697), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n207), .B2(new_n773), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT113), .Z(new_n1042));
  NOR2_X1   g0842(.A1(new_n718), .A2(new_n271), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1008), .B1(new_n203), .B2(new_n707), .C1(new_n918), .C2(new_n692), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(G116), .B2(new_n703), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1042), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT114), .Z(new_n1047));
  XOR2_X1   g0847(.A(KEYINPUT54), .B(G143), .Z(new_n1048));
  NAND2_X1  g0848(.A1(new_n704), .A2(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n711), .A2(G137), .B1(G125), .B2(new_n693), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n715), .A2(G159), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(G128), .B2(new_n697), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n271), .B1(new_n707), .B2(new_n201), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT112), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(G132), .B2(new_n703), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n708), .A2(new_n772), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT53), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1053), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1047), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n748), .B1(new_n1060), .B2(new_n731), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1039), .B(new_n1061), .C1(new_n360), .C2(new_n787), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1038), .A2(new_n1062), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n518), .B(G330), .C1(new_n677), .C2(new_n792), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1064), .A2(new_n857), .A3(new_n438), .A4(new_n607), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n873), .A2(new_n801), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n881), .A2(new_n800), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1066), .A2(new_n853), .A3(new_n1023), .A4(new_n1067), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n873), .A2(new_n801), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n881), .A2(new_n800), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1024), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1065), .B1(new_n1068), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(new_n1033), .B2(new_n1037), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1033), .A2(new_n1037), .A3(new_n1072), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT111), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1033), .A2(new_n1037), .A3(new_n1072), .A4(KEYINPUT111), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1073), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1063), .B1(new_n1078), .B2(new_n651), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(G378));
  OR3_X1    g0880(.A1(new_n847), .A2(new_n1022), .A3(new_n851), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n407), .A2(new_n408), .A3(new_n438), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT118), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n376), .A2(new_n810), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1083), .B(new_n1084), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1085), .B(new_n1086), .ZN(new_n1087));
  AND3_X1   g0887(.A1(new_n876), .A2(new_n884), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1087), .B1(new_n876), .B2(new_n884), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1081), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1087), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n869), .A2(new_n875), .A3(new_n860), .ZN(new_n1092));
  AOI21_X1  g0892(.A(KEYINPUT100), .B1(new_n880), .B2(new_n883), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1091), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NOR3_X1   g0894(.A1(new_n847), .A2(new_n851), .A3(new_n1022), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n876), .A2(new_n884), .A3(new_n1087), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1090), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1065), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AND3_X1   g0901(.A1(new_n1098), .A2(new_n1101), .A3(KEYINPUT57), .ZN(new_n1102));
  AOI21_X1  g0902(.A(KEYINPUT57), .B1(new_n1098), .B2(new_n1101), .ZN(new_n1103));
  NOR3_X1   g0903(.A1(new_n1102), .A2(new_n1103), .A3(new_n652), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1087), .A2(new_n741), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n768), .A2(new_n215), .B1(new_n708), .B2(new_n220), .ZN(new_n1106));
  NOR3_X1   g0906(.A1(new_n904), .A2(G41), .A3(new_n271), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n706), .B2(new_n692), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n1106), .B(new_n1108), .C1(G97), .C2(new_n711), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n726), .A2(new_n439), .B1(new_n207), .B2(new_n702), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1109), .B(new_n1111), .C1(new_n202), .C2(new_n707), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1112), .B(KEYINPUT58), .Z(new_n1113));
  AOI22_X1  g0913(.A1(new_n711), .A2(G132), .B1(new_n697), .B2(G125), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1048), .ZN(new_n1115));
  OAI21_X1  g0915(.A(KEYINPUT116), .B1(new_n1115), .B2(new_n708), .ZN(new_n1116));
  OR3_X1    g0916(.A1(new_n1115), .A2(KEYINPUT116), .A3(new_n708), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n1114), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(G128), .A2(new_n703), .B1(new_n704), .B2(G137), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1118), .B(new_n1119), .C1(new_n772), .C2(new_n728), .ZN(new_n1120));
  OR2_X1    g0920(.A1(new_n1120), .A2(KEYINPUT59), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n693), .A2(G124), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1120), .A2(KEYINPUT59), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n275), .A2(new_n649), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT115), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(G159), .B2(new_n982), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .A4(new_n1126), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1125), .B(new_n201), .C1(G41), .C2(new_n271), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n731), .B1(new_n1113), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n748), .B1(new_n201), .B2(new_n786), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT117), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1105), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(new_n1098), .B2(new_n946), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1104), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(G375));
  NAND2_X1  g0938(.A1(new_n1071), .A2(new_n1068), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n801), .A2(new_n741), .ZN(new_n1140));
  INV_X1    g0940(.A(G128), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n271), .B1(new_n692), .B2(new_n1141), .C1(new_n202), .C2(new_n707), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n728), .A2(new_n201), .B1(new_n708), .B2(new_n474), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n1142), .B(new_n1143), .C1(G132), .C2(new_n697), .ZN(new_n1144));
  INV_X1    g0944(.A(G137), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n1144), .B1(new_n1145), .B2(new_n725), .C1(new_n772), .C2(new_n726), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(new_n711), .B2(new_n1048), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n711), .A2(G116), .B1(new_n715), .B2(new_n259), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n271), .B1(new_n982), .B2(G77), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1148), .B(new_n1149), .C1(new_n918), .C2(new_n768), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n704), .A2(G107), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT121), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n708), .A2(new_n206), .B1(new_n692), .B2(new_n709), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n1151), .B1(new_n1152), .B2(new_n1153), .C1(new_n706), .C2(new_n702), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n1150), .B(new_n1154), .C1(new_n1152), .C2(new_n1153), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n731), .B1(new_n1147), .B2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n787), .A2(G68), .ZN(new_n1157));
  OAI21_X1  g0957(.A(KEYINPUT120), .B1(new_n748), .B2(new_n1157), .ZN(new_n1158));
  OR3_X1    g0958(.A1(new_n748), .A2(KEYINPUT120), .A3(new_n1157), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1156), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  XOR2_X1   g0960(.A(new_n1160), .B(KEYINPUT122), .Z(new_n1161));
  AOI22_X1  g0961(.A1(new_n1139), .A2(new_n946), .B1(new_n1140), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1071), .A2(new_n1065), .A3(new_n1068), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT119), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1164), .B(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1167), .A2(new_n1072), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1163), .B1(new_n1168), .B2(new_n926), .ZN(new_n1169));
  XOR2_X1   g0969(.A(new_n1169), .B(KEYINPUT123), .Z(G381));
  NOR4_X1   g0970(.A1(G387), .A2(G381), .A3(G396), .A4(G393), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1137), .A2(new_n1079), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(G390), .A2(G384), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1171), .A2(new_n1173), .A3(new_n1174), .ZN(G407));
  OAI211_X1 g0975(.A(G407), .B(G213), .C1(G343), .C2(new_n1172), .ZN(G409));
  OAI21_X1  g0976(.A(G378), .B1(new_n1104), .B2(new_n1136), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1164), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(KEYINPUT60), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT60), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1072), .A2(new_n1180), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n651), .B(new_n1179), .C1(new_n1167), .C2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n1162), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1183), .A2(new_n762), .A3(new_n789), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1182), .A2(G384), .A3(new_n1162), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n627), .A2(G213), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1098), .A2(new_n946), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1189), .A2(new_n1079), .A3(new_n1133), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(KEYINPUT124), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT124), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1097), .A2(new_n1090), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n1135), .A2(new_n1192), .B1(new_n1193), .B2(new_n926), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1188), .B1(new_n1191), .B2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1177), .A2(new_n1186), .A3(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(KEYINPUT62), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT61), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1188), .A2(G2897), .ZN(new_n1199));
  AND3_X1   g0999(.A1(new_n1184), .A2(new_n1185), .A3(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1199), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1191), .A2(new_n1194), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n1187), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1103), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1193), .A2(KEYINPUT57), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1205), .A2(new_n651), .A3(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1079), .B1(new_n1207), .B2(new_n1135), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1202), .B1(new_n1204), .B2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT62), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1177), .A2(new_n1195), .A3(new_n1210), .A4(new_n1186), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1197), .A2(new_n1198), .A3(new_n1209), .A4(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(KEYINPUT125), .ZN(new_n1213));
  XOR2_X1   g1013(.A(G393), .B(G396), .Z(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(G390), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(G387), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1177), .A2(new_n1195), .ZN(new_n1217));
  AOI21_X1  g1017(.A(KEYINPUT61), .B1(new_n1217), .B2(new_n1202), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT125), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1218), .A2(new_n1197), .A3(new_n1219), .A4(new_n1211), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1213), .A2(new_n1216), .A3(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1209), .A2(KEYINPUT63), .ZN(new_n1222));
  AOI21_X1  g1022(.A(KEYINPUT61), .B1(new_n1222), .B2(new_n1196), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT63), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1196), .A2(new_n1224), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1216), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1223), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1221), .A2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(KEYINPUT126), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT126), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1221), .A2(new_n1230), .A3(new_n1227), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1229), .A2(new_n1231), .ZN(G405));
  NAND2_X1  g1032(.A1(new_n1172), .A2(new_n1177), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT127), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1186), .A2(new_n1234), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1233), .B(new_n1235), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(new_n1236), .B(new_n1216), .ZN(G402));
endmodule


