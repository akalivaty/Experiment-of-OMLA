

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582;

  XNOR2_X1 U321 ( .A(n393), .B(n338), .ZN(n571) );
  XNOR2_X2 U322 ( .A(n339), .B(n571), .ZN(n500) );
  XNOR2_X1 U323 ( .A(KEYINPUT48), .B(KEYINPUT116), .ZN(n387) );
  XOR2_X1 U324 ( .A(G99GAT), .B(G85GAT), .Z(n341) );
  XNOR2_X1 U325 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U326 ( .A(n349), .B(n348), .ZN(n353) );
  XNOR2_X1 U327 ( .A(n388), .B(n387), .ZN(n523) );
  NOR2_X1 U328 ( .A1(n526), .A2(n447), .ZN(n560) );
  XOR2_X1 U329 ( .A(n307), .B(n306), .Z(n526) );
  XNOR2_X1 U330 ( .A(n448), .B(G190GAT), .ZN(n449) );
  XNOR2_X1 U331 ( .A(n450), .B(n449), .ZN(G1351GAT) );
  XOR2_X1 U332 ( .A(KEYINPUT83), .B(KEYINPUT84), .Z(n290) );
  XNOR2_X1 U333 ( .A(G169GAT), .B(KEYINPUT20), .ZN(n289) );
  XNOR2_X1 U334 ( .A(n290), .B(n289), .ZN(n307) );
  XOR2_X1 U335 ( .A(G190GAT), .B(G134GAT), .Z(n292) );
  XNOR2_X1 U336 ( .A(G43GAT), .B(G99GAT), .ZN(n291) );
  XNOR2_X1 U337 ( .A(n292), .B(n291), .ZN(n296) );
  XOR2_X1 U338 ( .A(G176GAT), .B(G127GAT), .Z(n294) );
  XNOR2_X1 U339 ( .A(G15GAT), .B(G120GAT), .ZN(n293) );
  XNOR2_X1 U340 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U341 ( .A(n296), .B(n295), .Z(n305) );
  XOR2_X1 U342 ( .A(KEYINPUT82), .B(KEYINPUT17), .Z(n298) );
  XNOR2_X1 U343 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n297) );
  XNOR2_X1 U344 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U345 ( .A(KEYINPUT19), .B(n299), .Z(n403) );
  XNOR2_X1 U346 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n300) );
  XNOR2_X1 U347 ( .A(n300), .B(KEYINPUT81), .ZN(n415) );
  XOR2_X1 U348 ( .A(n415), .B(G71GAT), .Z(n302) );
  NAND2_X1 U349 ( .A1(G227GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U351 ( .A(n403), .B(n303), .ZN(n304) );
  XNOR2_X1 U352 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U353 ( .A(G1GAT), .B(G113GAT), .Z(n309) );
  XNOR2_X1 U354 ( .A(G197GAT), .B(G141GAT), .ZN(n308) );
  XNOR2_X1 U355 ( .A(n309), .B(n308), .ZN(n324) );
  XOR2_X1 U356 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n311) );
  XNOR2_X1 U357 ( .A(KEYINPUT29), .B(KEYINPUT67), .ZN(n310) );
  XNOR2_X1 U358 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U359 ( .A(G36GAT), .B(G29GAT), .Z(n313) );
  XOR2_X1 U360 ( .A(G22GAT), .B(G15GAT), .Z(n361) );
  XOR2_X1 U361 ( .A(G169GAT), .B(G8GAT), .Z(n397) );
  XNOR2_X1 U362 ( .A(n361), .B(n397), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U364 ( .A(n315), .B(n314), .Z(n317) );
  NAND2_X1 U365 ( .A1(G229GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U366 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U367 ( .A(n318), .B(KEYINPUT69), .Z(n322) );
  XOR2_X1 U368 ( .A(G43GAT), .B(G50GAT), .Z(n320) );
  XNOR2_X1 U369 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n319) );
  XNOR2_X1 U370 ( .A(n320), .B(n319), .ZN(n355) );
  XNOR2_X1 U371 ( .A(n355), .B(KEYINPUT70), .ZN(n321) );
  XNOR2_X1 U372 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U373 ( .A(n324), .B(n323), .ZN(n541) );
  INV_X1 U374 ( .A(n541), .ZN(n567) );
  XOR2_X1 U375 ( .A(KEYINPUT41), .B(KEYINPUT64), .Z(n339) );
  XOR2_X1 U376 ( .A(G92GAT), .B(G64GAT), .Z(n326) );
  XNOR2_X1 U377 ( .A(G204GAT), .B(KEYINPUT73), .ZN(n325) );
  XNOR2_X1 U378 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U379 ( .A(G176GAT), .B(n327), .Z(n393) );
  XNOR2_X1 U380 ( .A(G71GAT), .B(KEYINPUT71), .ZN(n328) );
  XNOR2_X1 U381 ( .A(n328), .B(KEYINPUT13), .ZN(n364) );
  XOR2_X1 U382 ( .A(n341), .B(n364), .Z(n330) );
  NAND2_X1 U383 ( .A1(G230GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U384 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U385 ( .A(n331), .B(KEYINPUT33), .ZN(n334) );
  XNOR2_X1 U386 ( .A(G120GAT), .B(G148GAT), .ZN(n332) );
  XNOR2_X1 U387 ( .A(n332), .B(G57GAT), .ZN(n422) );
  XOR2_X1 U388 ( .A(n422), .B(KEYINPUT31), .Z(n333) );
  XNOR2_X1 U389 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U390 ( .A(n335), .B(KEYINPUT32), .Z(n337) );
  XOR2_X1 U391 ( .A(G106GAT), .B(G78GAT), .Z(n437) );
  XNOR2_X1 U392 ( .A(n437), .B(KEYINPUT72), .ZN(n336) );
  XOR2_X1 U393 ( .A(n337), .B(n336), .Z(n338) );
  NAND2_X1 U394 ( .A1(n567), .A2(n500), .ZN(n340) );
  XNOR2_X1 U395 ( .A(KEYINPUT46), .B(n340), .ZN(n378) );
  XOR2_X1 U396 ( .A(KEYINPUT65), .B(n341), .Z(n343) );
  XOR2_X1 U397 ( .A(G29GAT), .B(G134GAT), .Z(n425) );
  XNOR2_X1 U398 ( .A(G218GAT), .B(n425), .ZN(n342) );
  XNOR2_X1 U399 ( .A(n343), .B(n342), .ZN(n349) );
  XOR2_X1 U400 ( .A(KEYINPUT66), .B(KEYINPUT75), .Z(n345) );
  XNOR2_X1 U401 ( .A(G106GAT), .B(KEYINPUT9), .ZN(n344) );
  XOR2_X1 U402 ( .A(n345), .B(n344), .Z(n347) );
  NAND2_X1 U403 ( .A1(G232GAT), .A2(G233GAT), .ZN(n346) );
  XOR2_X1 U404 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n351) );
  XNOR2_X1 U405 ( .A(G162GAT), .B(G92GAT), .ZN(n350) );
  XOR2_X1 U406 ( .A(n351), .B(n350), .Z(n352) );
  XNOR2_X1 U407 ( .A(n353), .B(n352), .ZN(n357) );
  XNOR2_X1 U408 ( .A(G36GAT), .B(G190GAT), .ZN(n354) );
  XNOR2_X1 U409 ( .A(n354), .B(KEYINPUT76), .ZN(n389) );
  XNOR2_X1 U410 ( .A(n355), .B(n389), .ZN(n356) );
  XOR2_X1 U411 ( .A(n357), .B(n356), .Z(n552) );
  INV_X1 U412 ( .A(n552), .ZN(n535) );
  XOR2_X1 U413 ( .A(G64GAT), .B(G57GAT), .Z(n359) );
  XNOR2_X1 U414 ( .A(G211GAT), .B(G155GAT), .ZN(n358) );
  XNOR2_X1 U415 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U416 ( .A(n360), .B(G78GAT), .Z(n363) );
  XNOR2_X1 U417 ( .A(n361), .B(G183GAT), .ZN(n362) );
  XNOR2_X1 U418 ( .A(n363), .B(n362), .ZN(n368) );
  XOR2_X1 U419 ( .A(G1GAT), .B(G127GAT), .Z(n424) );
  XOR2_X1 U420 ( .A(n364), .B(n424), .Z(n366) );
  NAND2_X1 U421 ( .A1(G231GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U422 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U423 ( .A(n368), .B(n367), .Z(n376) );
  XOR2_X1 U424 ( .A(KEYINPUT15), .B(KEYINPUT79), .Z(n370) );
  XNOR2_X1 U425 ( .A(G8GAT), .B(KEYINPUT80), .ZN(n369) );
  XNOR2_X1 U426 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U427 ( .A(KEYINPUT77), .B(KEYINPUT78), .Z(n372) );
  XNOR2_X1 U428 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n371) );
  XNOR2_X1 U429 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U430 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U431 ( .A(n376), .B(n375), .Z(n549) );
  INV_X1 U432 ( .A(n549), .ZN(n575) );
  NOR2_X1 U433 ( .A1(n535), .A2(n575), .ZN(n377) );
  NAND2_X1 U434 ( .A1(n378), .A2(n377), .ZN(n379) );
  XNOR2_X1 U435 ( .A(n379), .B(KEYINPUT47), .ZN(n386) );
  XNOR2_X1 U436 ( .A(KEYINPUT36), .B(KEYINPUT107), .ZN(n380) );
  XOR2_X1 U437 ( .A(n552), .B(n380), .Z(n579) );
  NOR2_X1 U438 ( .A1(n579), .A2(n549), .ZN(n381) );
  XOR2_X1 U439 ( .A(KEYINPUT45), .B(n381), .Z(n382) );
  NOR2_X1 U440 ( .A1(n571), .A2(n382), .ZN(n383) );
  XNOR2_X1 U441 ( .A(KEYINPUT115), .B(n383), .ZN(n384) );
  NOR2_X1 U442 ( .A1(n384), .A2(n567), .ZN(n385) );
  NOR2_X1 U443 ( .A1(n386), .A2(n385), .ZN(n388) );
  XOR2_X1 U444 ( .A(n389), .B(KEYINPUT96), .Z(n391) );
  NAND2_X1 U445 ( .A1(G226GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U446 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U447 ( .A(n393), .B(n392), .ZN(n401) );
  XOR2_X1 U448 ( .A(KEYINPUT95), .B(KEYINPUT77), .Z(n399) );
  XOR2_X1 U449 ( .A(KEYINPUT87), .B(G218GAT), .Z(n395) );
  XNOR2_X1 U450 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n394) );
  XNOR2_X1 U451 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U452 ( .A(G197GAT), .B(n396), .Z(n441) );
  XNOR2_X1 U453 ( .A(n397), .B(n441), .ZN(n398) );
  XNOR2_X1 U454 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U455 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U456 ( .A(n403), .B(n402), .ZN(n516) );
  NOR2_X1 U457 ( .A1(n523), .A2(n516), .ZN(n404) );
  XNOR2_X1 U458 ( .A(n404), .B(KEYINPUT54), .ZN(n563) );
  XOR2_X1 U459 ( .A(KEYINPUT90), .B(KEYINPUT5), .Z(n406) );
  XNOR2_X1 U460 ( .A(G85GAT), .B(KEYINPUT1), .ZN(n405) );
  XNOR2_X1 U461 ( .A(n406), .B(n405), .ZN(n410) );
  XOR2_X1 U462 ( .A(KEYINPUT4), .B(KEYINPUT92), .Z(n408) );
  XNOR2_X1 U463 ( .A(KEYINPUT93), .B(KEYINPUT6), .ZN(n407) );
  XNOR2_X1 U464 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U465 ( .A(n410), .B(n409), .Z(n421) );
  XOR2_X1 U466 ( .A(KEYINPUT2), .B(KEYINPUT88), .Z(n412) );
  XNOR2_X1 U467 ( .A(G141GAT), .B(G155GAT), .ZN(n411) );
  XNOR2_X1 U468 ( .A(n412), .B(n411), .ZN(n414) );
  XOR2_X1 U469 ( .A(G162GAT), .B(KEYINPUT3), .Z(n413) );
  XOR2_X1 U470 ( .A(n414), .B(n413), .Z(n442) );
  INV_X1 U471 ( .A(n442), .ZN(n419) );
  XOR2_X1 U472 ( .A(n415), .B(KEYINPUT91), .Z(n417) );
  NAND2_X1 U473 ( .A1(G225GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U474 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U475 ( .A(n419), .B(n418), .Z(n420) );
  XNOR2_X1 U476 ( .A(n421), .B(n420), .ZN(n423) );
  XOR2_X1 U477 ( .A(n423), .B(n422), .Z(n427) );
  XNOR2_X1 U478 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U479 ( .A(n427), .B(n426), .ZN(n467) );
  XNOR2_X1 U480 ( .A(KEYINPUT94), .B(n467), .ZN(n562) );
  XOR2_X1 U481 ( .A(G204GAT), .B(KEYINPUT24), .Z(n429) );
  XNOR2_X1 U482 ( .A(G50GAT), .B(KEYINPUT23), .ZN(n428) );
  XNOR2_X1 U483 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U484 ( .A(KEYINPUT85), .B(KEYINPUT86), .Z(n431) );
  XNOR2_X1 U485 ( .A(G22GAT), .B(G148GAT), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U487 ( .A(n433), .B(n432), .Z(n439) );
  XOR2_X1 U488 ( .A(KEYINPUT22), .B(KEYINPUT89), .Z(n435) );
  NAND2_X1 U489 ( .A1(G228GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U490 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U492 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U493 ( .A(n441), .B(n440), .ZN(n443) );
  XOR2_X1 U494 ( .A(n443), .B(n442), .Z(n462) );
  INV_X1 U495 ( .A(n462), .ZN(n444) );
  AND2_X1 U496 ( .A1(n562), .A2(n444), .ZN(n445) );
  AND2_X1 U497 ( .A1(n563), .A2(n445), .ZN(n446) );
  XNOR2_X1 U498 ( .A(n446), .B(KEYINPUT55), .ZN(n447) );
  NAND2_X1 U499 ( .A1(n560), .A2(n535), .ZN(n450) );
  XOR2_X1 U500 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n448) );
  NOR2_X1 U501 ( .A1(n535), .A2(n549), .ZN(n451) );
  XNOR2_X1 U502 ( .A(KEYINPUT16), .B(n451), .ZN(n472) );
  XOR2_X1 U503 ( .A(KEYINPUT28), .B(n462), .Z(n524) );
  INV_X1 U504 ( .A(n524), .ZN(n454) );
  XOR2_X1 U505 ( .A(KEYINPUT27), .B(n516), .Z(n460) );
  INV_X1 U506 ( .A(n460), .ZN(n452) );
  NOR2_X1 U507 ( .A1(n562), .A2(n452), .ZN(n453) );
  XNOR2_X1 U508 ( .A(n453), .B(KEYINPUT97), .ZN(n522) );
  NOR2_X1 U509 ( .A1(n454), .A2(n522), .ZN(n455) );
  NAND2_X1 U510 ( .A1(n526), .A2(n455), .ZN(n456) );
  XNOR2_X1 U511 ( .A(n456), .B(KEYINPUT98), .ZN(n470) );
  XOR2_X1 U512 ( .A(KEYINPUT100), .B(KEYINPUT26), .Z(n458) );
  NAND2_X1 U513 ( .A1(n526), .A2(n462), .ZN(n457) );
  XNOR2_X1 U514 ( .A(n458), .B(n457), .ZN(n459) );
  XOR2_X1 U515 ( .A(KEYINPUT99), .B(n459), .Z(n564) );
  NAND2_X1 U516 ( .A1(n460), .A2(n564), .ZN(n466) );
  NOR2_X1 U517 ( .A1(n526), .A2(n516), .ZN(n461) );
  NOR2_X1 U518 ( .A1(n462), .A2(n461), .ZN(n463) );
  XOR2_X1 U519 ( .A(n463), .B(KEYINPUT25), .Z(n464) );
  XNOR2_X1 U520 ( .A(KEYINPUT101), .B(n464), .ZN(n465) );
  NAND2_X1 U521 ( .A1(n466), .A2(n465), .ZN(n468) );
  NAND2_X1 U522 ( .A1(n468), .A2(n467), .ZN(n469) );
  NAND2_X1 U523 ( .A1(n470), .A2(n469), .ZN(n471) );
  XNOR2_X1 U524 ( .A(KEYINPUT102), .B(n471), .ZN(n486) );
  NAND2_X1 U525 ( .A1(n472), .A2(n486), .ZN(n473) );
  XNOR2_X1 U526 ( .A(n473), .B(KEYINPUT103), .ZN(n502) );
  OR2_X1 U527 ( .A1(n571), .A2(n541), .ZN(n474) );
  XOR2_X1 U528 ( .A(KEYINPUT74), .B(n474), .Z(n489) );
  NAND2_X1 U529 ( .A1(n502), .A2(n489), .ZN(n483) );
  NOR2_X1 U530 ( .A1(n562), .A2(n483), .ZN(n476) );
  XNOR2_X1 U531 ( .A(KEYINPUT34), .B(KEYINPUT104), .ZN(n475) );
  XNOR2_X1 U532 ( .A(n476), .B(n475), .ZN(n477) );
  XOR2_X1 U533 ( .A(G1GAT), .B(n477), .Z(G1324GAT) );
  NOR2_X1 U534 ( .A1(n516), .A2(n483), .ZN(n479) );
  XNOR2_X1 U535 ( .A(G8GAT), .B(KEYINPUT105), .ZN(n478) );
  XNOR2_X1 U536 ( .A(n479), .B(n478), .ZN(G1325GAT) );
  NOR2_X1 U537 ( .A1(n526), .A2(n483), .ZN(n481) );
  XNOR2_X1 U538 ( .A(KEYINPUT106), .B(KEYINPUT35), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U540 ( .A(G15GAT), .B(n482), .ZN(G1326GAT) );
  NOR2_X1 U541 ( .A1(n524), .A2(n483), .ZN(n484) );
  XOR2_X1 U542 ( .A(G22GAT), .B(n484), .Z(G1327GAT) );
  NOR2_X1 U543 ( .A1(n579), .A2(n575), .ZN(n485) );
  NAND2_X1 U544 ( .A1(n486), .A2(n485), .ZN(n487) );
  XNOR2_X1 U545 ( .A(KEYINPUT37), .B(n487), .ZN(n488) );
  XNOR2_X1 U546 ( .A(KEYINPUT108), .B(n488), .ZN(n512) );
  NAND2_X1 U547 ( .A1(n512), .A2(n489), .ZN(n490) );
  XNOR2_X1 U548 ( .A(KEYINPUT38), .B(n490), .ZN(n498) );
  NOR2_X1 U549 ( .A1(n498), .A2(n562), .ZN(n492) );
  XNOR2_X1 U550 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n491) );
  XNOR2_X1 U551 ( .A(n492), .B(n491), .ZN(G1328GAT) );
  NOR2_X1 U552 ( .A1(n498), .A2(n516), .ZN(n493) );
  XOR2_X1 U553 ( .A(G36GAT), .B(n493), .Z(G1329GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT40), .B(KEYINPUT110), .Z(n495) );
  XNOR2_X1 U555 ( .A(G43GAT), .B(KEYINPUT109), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n495), .B(n494), .ZN(n497) );
  NOR2_X1 U557 ( .A1(n526), .A2(n498), .ZN(n496) );
  XOR2_X1 U558 ( .A(n497), .B(n496), .Z(G1330GAT) );
  NOR2_X1 U559 ( .A1(n498), .A2(n524), .ZN(n499) );
  XOR2_X1 U560 ( .A(G50GAT), .B(n499), .Z(G1331GAT) );
  NAND2_X1 U561 ( .A1(n500), .A2(n541), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n501), .B(KEYINPUT111), .ZN(n513) );
  NAND2_X1 U563 ( .A1(n502), .A2(n513), .ZN(n509) );
  NOR2_X1 U564 ( .A1(n562), .A2(n509), .ZN(n503) );
  XOR2_X1 U565 ( .A(KEYINPUT42), .B(n503), .Z(n504) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(n504), .ZN(G1332GAT) );
  NOR2_X1 U567 ( .A1(n516), .A2(n509), .ZN(n505) );
  XOR2_X1 U568 ( .A(KEYINPUT112), .B(n505), .Z(n506) );
  XNOR2_X1 U569 ( .A(G64GAT), .B(n506), .ZN(G1333GAT) );
  NOR2_X1 U570 ( .A1(n526), .A2(n509), .ZN(n508) );
  XNOR2_X1 U571 ( .A(G71GAT), .B(KEYINPUT113), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n508), .B(n507), .ZN(G1334GAT) );
  NOR2_X1 U573 ( .A1(n524), .A2(n509), .ZN(n511) );
  XNOR2_X1 U574 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n511), .B(n510), .ZN(G1335GAT) );
  NAND2_X1 U576 ( .A1(n513), .A2(n512), .ZN(n519) );
  NOR2_X1 U577 ( .A1(n562), .A2(n519), .ZN(n514) );
  XOR2_X1 U578 ( .A(G85GAT), .B(n514), .Z(n515) );
  XNOR2_X1 U579 ( .A(KEYINPUT114), .B(n515), .ZN(G1336GAT) );
  NOR2_X1 U580 ( .A1(n516), .A2(n519), .ZN(n517) );
  XOR2_X1 U581 ( .A(G92GAT), .B(n517), .Z(G1337GAT) );
  NOR2_X1 U582 ( .A1(n526), .A2(n519), .ZN(n518) );
  XOR2_X1 U583 ( .A(G99GAT), .B(n518), .Z(G1338GAT) );
  NOR2_X1 U584 ( .A1(n524), .A2(n519), .ZN(n520) );
  XOR2_X1 U585 ( .A(KEYINPUT44), .B(n520), .Z(n521) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(n521), .ZN(G1339GAT) );
  NOR2_X1 U587 ( .A1(n523), .A2(n522), .ZN(n540) );
  NAND2_X1 U588 ( .A1(n540), .A2(n524), .ZN(n525) );
  NOR2_X1 U589 ( .A1(n526), .A2(n525), .ZN(n536) );
  NAND2_X1 U590 ( .A1(n567), .A2(n536), .ZN(n527) );
  XNOR2_X1 U591 ( .A(G113GAT), .B(n527), .ZN(G1340GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n529) );
  NAND2_X1 U593 ( .A1(n536), .A2(n500), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U595 ( .A(G120GAT), .B(n530), .Z(G1341GAT) );
  XNOR2_X1 U596 ( .A(G127GAT), .B(KEYINPUT119), .ZN(n534) );
  XOR2_X1 U597 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n532) );
  NAND2_X1 U598 ( .A1(n536), .A2(n575), .ZN(n531) );
  XNOR2_X1 U599 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(G1342GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT51), .B(KEYINPUT120), .Z(n538) );
  NAND2_X1 U602 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U604 ( .A(G134GAT), .B(n539), .ZN(G1343GAT) );
  NAND2_X1 U605 ( .A1(n564), .A2(n540), .ZN(n551) );
  NOR2_X1 U606 ( .A1(n541), .A2(n551), .ZN(n543) );
  XNOR2_X1 U607 ( .A(G141GAT), .B(KEYINPUT121), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(G1344GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT122), .B(KEYINPUT52), .Z(n545) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n548) );
  INV_X1 U612 ( .A(n500), .ZN(n546) );
  NOR2_X1 U613 ( .A1(n546), .A2(n551), .ZN(n547) );
  XOR2_X1 U614 ( .A(n548), .B(n547), .Z(G1345GAT) );
  NOR2_X1 U615 ( .A1(n549), .A2(n551), .ZN(n550) );
  XOR2_X1 U616 ( .A(G155GAT), .B(n550), .Z(G1346GAT) );
  NOR2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n554) );
  XNOR2_X1 U618 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U620 ( .A(G162GAT), .B(n555), .ZN(G1347GAT) );
  NAND2_X1 U621 ( .A1(n567), .A2(n560), .ZN(n556) );
  XNOR2_X1 U622 ( .A(G169GAT), .B(n556), .ZN(G1348GAT) );
  NAND2_X1 U623 ( .A1(n560), .A2(n500), .ZN(n558) );
  XOR2_X1 U624 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(G176GAT), .B(n559), .ZN(G1349GAT) );
  NAND2_X1 U627 ( .A1(n560), .A2(n575), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n569) );
  NAND2_X1 U630 ( .A1(n563), .A2(n562), .ZN(n566) );
  INV_X1 U631 ( .A(n564), .ZN(n565) );
  NOR2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n577) );
  NAND2_X1 U633 ( .A1(n577), .A2(n567), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(n570), .ZN(G1352GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n573) );
  NAND2_X1 U637 ( .A1(n577), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(G204GAT), .B(n574), .ZN(G1353GAT) );
  NAND2_X1 U640 ( .A1(n577), .A2(n575), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U642 ( .A(n577), .ZN(n578) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n581) );
  XNOR2_X1 U644 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

