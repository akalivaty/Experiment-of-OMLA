//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 0 0 1 0 0 0 1 0 0 1 0 0 1 0 1 1 0 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 0 1 1 1 0 1 0 1 1 0 1 1 1 0 1 1 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT69), .B(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(G210), .A3(new_n189), .ZN(new_n190));
  XOR2_X1   g004(.A(new_n190), .B(KEYINPUT27), .Z(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT26), .B(G101), .ZN(new_n192));
  XOR2_X1   g006(.A(new_n191), .B(new_n192), .Z(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT1), .B1(new_n194), .B2(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G128), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G143), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n194), .A2(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n196), .A2(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(G143), .B(G146), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(G128), .A3(new_n195), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G134), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT64), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G134), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n206), .A2(new_n208), .A3(G137), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n210));
  INV_X1    g024(.A(G137), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(KEYINPUT65), .A2(G137), .ZN(new_n213));
  AND2_X1   g027(.A1(KEYINPUT11), .A2(G134), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(G137), .B1(new_n206), .B2(new_n208), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n209), .B(new_n215), .C1(new_n216), .C2(KEYINPUT11), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n204), .B1(new_n217), .B2(G131), .ZN(new_n218));
  INV_X1    g032(.A(G131), .ZN(new_n219));
  AOI21_X1  g033(.A(G134), .B1(new_n212), .B2(new_n213), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n206), .A2(new_n208), .ZN(new_n221));
  AOI22_X1  g035(.A1(new_n220), .A2(KEYINPUT66), .B1(new_n221), .B2(new_n211), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT65), .B(G137), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(new_n205), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n219), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT67), .B1(new_n218), .B2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n223), .A2(KEYINPUT66), .A3(new_n205), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n221), .A2(new_n211), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n220), .A2(KEYINPUT66), .ZN(new_n232));
  OAI21_X1  g046(.A(G131), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT67), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT11), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT64), .B(G134), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n235), .B1(new_n236), .B2(G137), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n237), .A2(new_n219), .A3(new_n209), .A4(new_n215), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n233), .A2(new_n234), .A3(new_n238), .A4(new_n204), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT11), .B1(new_n221), .B2(new_n211), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n209), .A2(new_n215), .ZN(new_n241));
  OAI21_X1  g055(.A(G131), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n238), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n202), .A2(KEYINPUT0), .A3(G128), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT0), .B(G128), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n244), .B1(new_n202), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G119), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G116), .ZN(new_n250));
  INV_X1    g064(.A(G116), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G119), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT2), .B(G113), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n253), .A2(new_n255), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n228), .A2(new_n239), .A3(new_n248), .A4(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n228), .A2(new_n239), .A3(new_n248), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT30), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n218), .A2(new_n227), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n246), .B1(new_n242), .B2(new_n238), .ZN(new_n267));
  OR3_X1    g081(.A1(new_n266), .A2(new_n267), .A3(KEYINPUT30), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n263), .B1(new_n269), .B2(new_n259), .ZN(new_n270));
  AOI211_X1 g084(.A(new_n262), .B(new_n260), .C1(new_n265), .C2(new_n268), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n193), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT31), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI211_X1 g088(.A(KEYINPUT31), .B(new_n193), .C1(new_n270), .C2(new_n271), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n266), .A2(new_n267), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT28), .B1(new_n277), .B2(new_n260), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n259), .B1(new_n266), .B2(new_n267), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n261), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT28), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n278), .B1(new_n281), .B2(KEYINPUT70), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT70), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n280), .A2(new_n283), .A3(KEYINPUT28), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n193), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT71), .B1(new_n276), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT71), .ZN(new_n288));
  AOI211_X1 g102(.A(new_n288), .B(new_n285), .C1(new_n274), .C2(new_n275), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n187), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT32), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI211_X1 g106(.A(KEYINPUT32), .B(new_n187), .C1(new_n287), .C2(new_n289), .ZN(new_n293));
  INV_X1    g107(.A(new_n270), .ZN(new_n294));
  INV_X1    g108(.A(new_n271), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(KEYINPUT72), .B1(new_n296), .B2(new_n193), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT29), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT72), .ZN(new_n299));
  INV_X1    g113(.A(new_n193), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n294), .A2(new_n299), .A3(new_n300), .A4(new_n295), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n282), .A2(new_n193), .A3(new_n284), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n297), .A2(new_n298), .A3(new_n301), .A4(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n264), .A2(new_n259), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n261), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n278), .B1(new_n305), .B2(KEYINPUT28), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n300), .A2(new_n298), .ZN(new_n307));
  AOI21_X1  g121(.A(G902), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G472), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n292), .A2(new_n293), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT86), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT81), .ZN(new_n313));
  INV_X1    g127(.A(G107), .ZN(new_n314));
  OAI22_X1  g128(.A1(new_n313), .A2(KEYINPUT3), .B1(new_n314), .B2(G104), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT3), .ZN(new_n316));
  INV_X1    g130(.A(G104), .ZN(new_n317));
  OAI22_X1  g131(.A1(KEYINPUT81), .A2(new_n316), .B1(new_n317), .B2(G107), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n313), .A2(new_n314), .A3(KEYINPUT3), .A4(G104), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n315), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(KEYINPUT4), .B1(new_n321), .B2(G101), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G101), .ZN(new_n324));
  AOI22_X1  g138(.A1(KEYINPUT81), .A2(new_n316), .B1(new_n317), .B2(G107), .ZN(new_n325));
  AND4_X1   g139(.A1(new_n313), .A2(new_n314), .A3(KEYINPUT3), .A4(G104), .ZN(new_n326));
  AOI22_X1  g140(.A1(new_n313), .A2(KEYINPUT3), .B1(new_n314), .B2(G104), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n324), .B(new_n325), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT82), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n320), .A2(KEYINPUT82), .A3(new_n324), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n330), .A2(new_n331), .B1(G101), .B2(new_n321), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT4), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n323), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(new_n247), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT83), .B1(new_n317), .B2(G107), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n336), .B1(new_n317), .B2(G107), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n317), .A2(G107), .ZN(new_n338));
  OAI21_X1  g152(.A(G101), .B1(new_n338), .B2(KEYINPUT83), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT1), .ZN(new_n341));
  AND4_X1   g155(.A1(new_n341), .A2(new_n198), .A3(new_n199), .A4(G128), .ZN(new_n342));
  AOI22_X1  g156(.A1(new_n195), .A2(G128), .B1(new_n198), .B2(new_n199), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI211_X1 g158(.A(new_n340), .B(new_n344), .C1(new_n330), .C2(new_n331), .ZN(new_n345));
  OAI21_X1  g159(.A(KEYINPUT10), .B1(new_n345), .B2(KEYINPUT84), .ZN(new_n346));
  INV_X1    g160(.A(new_n243), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n330), .A2(new_n331), .ZN(new_n348));
  INV_X1    g162(.A(new_n340), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(new_n204), .A3(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT84), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT10), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n335), .A2(new_n346), .A3(new_n347), .A4(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(G110), .B(G140), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n189), .A2(G227), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n355), .B(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n335), .A2(new_n346), .A3(new_n353), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n243), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  AND4_X1   g176(.A1(new_n347), .A2(new_n335), .A3(new_n346), .A4(new_n353), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT12), .ZN(new_n364));
  AOI21_X1  g178(.A(KEYINPUT82), .B1(new_n320), .B2(new_n324), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n318), .A2(new_n319), .ZN(new_n366));
  AND4_X1   g180(.A1(KEYINPUT82), .A2(new_n366), .A3(new_n324), .A4(new_n325), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n349), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n344), .ZN(new_n369));
  AOI211_X1 g183(.A(new_n364), .B(new_n347), .C1(new_n369), .C2(new_n350), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT85), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n204), .B1(new_n348), .B2(new_n349), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n243), .B1(new_n345), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n364), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n370), .B1(new_n371), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n373), .A2(KEYINPUT85), .A3(new_n364), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n363), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n312), .B(new_n362), .C1(new_n377), .C2(new_n358), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n347), .B1(new_n369), .B2(new_n350), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n371), .B1(new_n379), .B2(KEYINPUT12), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(KEYINPUT12), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n376), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n358), .B1(new_n382), .B2(new_n354), .ZN(new_n383));
  AND3_X1   g197(.A1(new_n361), .A2(new_n354), .A3(new_n358), .ZN(new_n384));
  OAI21_X1  g198(.A(KEYINPUT86), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n378), .A2(new_n385), .A3(G469), .ZN(new_n386));
  INV_X1    g200(.A(G469), .ZN(new_n387));
  INV_X1    g201(.A(G902), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n359), .A2(new_n382), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n340), .B1(new_n330), .B2(new_n331), .ZN(new_n391));
  AOI211_X1 g205(.A(KEYINPUT84), .B(KEYINPUT10), .C1(new_n391), .C2(new_n204), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n352), .B1(new_n350), .B2(new_n351), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n347), .B1(new_n394), .B2(new_n335), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n357), .B1(new_n395), .B2(new_n363), .ZN(new_n396));
  AOI21_X1  g210(.A(G902), .B1(new_n390), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n389), .B1(new_n397), .B2(new_n387), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n386), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G221), .ZN(new_n400));
  XNOR2_X1  g214(.A(KEYINPUT9), .B(G234), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n400), .B1(new_n402), .B2(new_n388), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n403), .B(KEYINPUT80), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n399), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(KEYINPUT87), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT87), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n399), .A2(new_n408), .A3(new_n405), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(G125), .B(G140), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT16), .ZN(new_n412));
  INV_X1    g226(.A(G125), .ZN(new_n413));
  OR3_X1    g227(.A1(new_n413), .A2(KEYINPUT16), .A3(G140), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n197), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n412), .A2(G146), .A3(new_n414), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  XOR2_X1   g232(.A(KEYINPUT24), .B(G110), .Z(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(KEYINPUT75), .ZN(new_n420));
  OR3_X1    g234(.A1(new_n249), .A2(KEYINPUT74), .A3(G128), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n249), .A2(G128), .ZN(new_n422));
  OAI21_X1  g236(.A(KEYINPUT74), .B1(new_n249), .B2(G128), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n418), .B1(new_n420), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT23), .ZN(new_n426));
  OR3_X1    g240(.A1(new_n426), .A2(new_n249), .A3(G128), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n426), .B1(new_n249), .B2(G128), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n428), .A3(new_n422), .ZN(new_n429));
  OR2_X1    g243(.A1(new_n429), .A2(KEYINPUT76), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(KEYINPUT76), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n430), .A2(new_n431), .A3(G110), .ZN(new_n432));
  OR2_X1    g246(.A1(new_n425), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n429), .ZN(new_n434));
  XOR2_X1   g248(.A(KEYINPUT77), .B(G110), .Z(new_n435));
  AOI22_X1  g249(.A1(new_n420), .A2(new_n424), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n411), .A2(new_n197), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n417), .A2(new_n437), .ZN(new_n438));
  OR2_X1    g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n433), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(KEYINPUT78), .ZN(new_n441));
  XNOR2_X1  g255(.A(KEYINPUT22), .B(G137), .ZN(new_n442));
  INV_X1    g256(.A(G234), .ZN(new_n443));
  NOR3_X1   g257(.A1(new_n400), .A2(new_n443), .A3(G953), .ZN(new_n444));
  XOR2_X1   g258(.A(new_n442), .B(new_n444), .Z(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT78), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n433), .A2(new_n447), .A3(new_n439), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n441), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(KEYINPUT79), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT79), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n441), .A2(new_n451), .A3(new_n446), .A4(new_n448), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n433), .A2(new_n445), .A3(new_n439), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n450), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NOR3_X1   g268(.A1(new_n454), .A2(KEYINPUT25), .A3(G902), .ZN(new_n455));
  OAI21_X1  g269(.A(G217), .B1(new_n443), .B2(G902), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n456), .B(KEYINPUT73), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(KEYINPUT25), .B1(new_n454), .B2(G902), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n457), .A2(new_n388), .ZN(new_n461));
  OR2_X1    g275(.A1(new_n454), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n247), .A2(G125), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n204), .A2(new_n413), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G224), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(G953), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT7), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OR3_X1    g285(.A1(new_n467), .A2(KEYINPUT92), .A3(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(KEYINPUT92), .B1(new_n467), .B2(new_n471), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n470), .B1(new_n469), .B2(KEYINPUT93), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n467), .B(new_n474), .C1(KEYINPUT93), .C2(new_n469), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n472), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(G113), .B1(new_n250), .B2(KEYINPUT5), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n254), .A2(KEYINPUT5), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n477), .B1(new_n478), .B2(KEYINPUT90), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n479), .B1(KEYINPUT90), .B2(new_n478), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n257), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(KEYINPUT91), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n391), .ZN(new_n483));
  XNOR2_X1  g297(.A(G110), .B(G122), .ZN(new_n484));
  XOR2_X1   g298(.A(new_n484), .B(KEYINPUT8), .Z(new_n485));
  INV_X1    g299(.A(new_n477), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n478), .A2(new_n486), .B1(new_n254), .B2(new_n256), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n485), .B1(new_n368), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n476), .B1(new_n483), .B2(new_n488), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n334), .A2(new_n259), .B1(new_n391), .B2(new_n487), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n484), .ZN(new_n491));
  AOI21_X1  g305(.A(G902), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n391), .A2(new_n487), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n321), .A2(G101), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n348), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n322), .B1(new_n495), .B2(KEYINPUT4), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n493), .B1(new_n496), .B2(new_n260), .ZN(new_n497));
  INV_X1    g311(.A(new_n484), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n497), .A2(KEYINPUT88), .A3(KEYINPUT6), .A4(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT6), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n500), .B1(new_n490), .B2(new_n484), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n498), .A2(KEYINPUT88), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n490), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n499), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT89), .ZN(new_n505));
  XOR2_X1   g319(.A(new_n467), .B(new_n469), .Z(new_n506));
  AND3_X1   g320(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n505), .B1(new_n504), .B2(new_n506), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n492), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(G210), .B1(G237), .B2(G902), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n510), .B(new_n492), .C1(new_n507), .C2(new_n508), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(G475), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n188), .A2(G214), .A3(new_n189), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n194), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n188), .A2(G143), .A3(G214), .A4(new_n189), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(KEYINPUT18), .A3(G131), .ZN(new_n521));
  NAND2_X1  g335(.A1(KEYINPUT18), .A2(G131), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n518), .A2(new_n519), .A3(new_n522), .ZN(new_n523));
  OR2_X1    g337(.A1(new_n411), .A2(KEYINPUT94), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n411), .A2(KEYINPUT94), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n525), .A3(G146), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n437), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n521), .A2(new_n523), .A3(new_n527), .ZN(new_n528));
  OR2_X1    g342(.A1(new_n418), .A2(KEYINPUT97), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n219), .B1(new_n518), .B2(new_n519), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT17), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n418), .A2(KEYINPUT97), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n529), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n520), .A2(G131), .ZN(new_n534));
  NOR3_X1   g348(.A1(new_n534), .A2(new_n530), .A3(KEYINPUT17), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n528), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  XNOR2_X1  g350(.A(G113), .B(G122), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT95), .B(G104), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n537), .B(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n539), .B(new_n528), .C1(new_n533), .C2(new_n535), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n516), .B1(new_n543), .B2(new_n388), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT19), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n546), .B1(new_n524), .B2(new_n525), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n411), .A2(KEYINPUT19), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n197), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n549), .B(new_n417), .C1(new_n534), .C2(new_n530), .ZN(new_n550));
  AOI211_X1 g364(.A(KEYINPUT96), .B(new_n539), .C1(new_n550), .C2(new_n528), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT96), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(new_n528), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n552), .B1(new_n553), .B2(new_n540), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n551), .B1(new_n554), .B2(new_n542), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT20), .ZN(new_n556));
  NOR2_X1   g370(.A1(G475), .A2(G902), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n556), .B1(new_n555), .B2(new_n557), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n545), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(G234), .A2(G237), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n562), .A2(G952), .A3(new_n189), .ZN(new_n563));
  XNOR2_X1  g377(.A(KEYINPUT21), .B(G898), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n562), .A2(G902), .A3(G953), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n563), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(KEYINPUT100), .ZN(new_n568));
  XNOR2_X1  g382(.A(G116), .B(G122), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(new_n314), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT13), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n571), .A2(new_n194), .A3(G128), .ZN(new_n572));
  XNOR2_X1  g386(.A(G128), .B(G143), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  OAI211_X1 g388(.A(G134), .B(new_n572), .C1(new_n574), .C2(new_n571), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n570), .B(new_n575), .C1(new_n221), .C2(new_n574), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n251), .A2(KEYINPUT14), .A3(G122), .ZN(new_n577));
  INV_X1    g391(.A(new_n569), .ZN(new_n578));
  OAI211_X1 g392(.A(G107), .B(new_n577), .C1(new_n578), .C2(KEYINPUT14), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n569), .A2(new_n314), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n574), .A2(new_n221), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n236), .A2(new_n573), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n579), .B(new_n580), .C1(new_n581), .C2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n576), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n402), .A2(G217), .A3(new_n189), .ZN(new_n585));
  OR2_X1    g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT98), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n584), .A2(new_n585), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n584), .A2(KEYINPUT98), .A3(new_n585), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n589), .A2(KEYINPUT99), .A3(new_n388), .A4(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(G478), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n592), .A2(KEYINPUT15), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n591), .B(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n561), .A2(new_n568), .A3(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(G214), .B1(G237), .B2(G902), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n515), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n311), .A2(new_n410), .A3(new_n464), .A4(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(G101), .ZN(G3));
  OAI21_X1  g415(.A(new_n388), .B1(new_n287), .B2(new_n289), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(G472), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n603), .A2(new_n290), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n604), .A2(new_n464), .A3(new_n410), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(KEYINPUT101), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n512), .A2(KEYINPUT102), .A3(new_n513), .ZN(new_n607));
  OR2_X1    g421(.A1(new_n507), .A2(new_n508), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT102), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n608), .A2(new_n609), .A3(new_n510), .A4(new_n492), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n607), .A2(new_n597), .A3(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT33), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT103), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n588), .A2(new_n614), .ZN(new_n615));
  OR2_X1    g429(.A1(new_n615), .A2(new_n586), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n586), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n613), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(KEYINPUT33), .B1(new_n589), .B2(new_n590), .ZN(new_n619));
  OAI211_X1 g433(.A(G478), .B(new_n388), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n589), .A2(new_n388), .A3(new_n590), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n592), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n560), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n568), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n606), .A2(new_n612), .A3(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT34), .B(G104), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G6));
  OAI211_X1 g443(.A(new_n545), .B(new_n594), .C1(new_n559), .C2(new_n558), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n606), .A2(new_n568), .A3(new_n612), .A4(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(KEYINPUT104), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT35), .B(G107), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G9));
  INV_X1    g449(.A(new_n461), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n441), .A2(new_n448), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n446), .A2(KEYINPUT36), .ZN(new_n638));
  XOR2_X1   g452(.A(new_n637), .B(new_n638), .Z(new_n639));
  AOI22_X1  g453(.A1(new_n458), .A2(new_n459), .B1(new_n636), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n604), .A2(new_n410), .A3(new_n599), .A4(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT37), .B(G110), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G12));
  OR2_X1    g458(.A1(new_n566), .A2(G900), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n563), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n631), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n647), .B1(new_n407), .B2(new_n409), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n611), .A2(new_n640), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n311), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(KEYINPUT105), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT105), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n311), .A2(new_n648), .A3(new_n649), .A4(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G128), .ZN(G30));
  AND2_X1   g469(.A1(new_n292), .A2(new_n293), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n296), .A2(new_n300), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n388), .B1(new_n305), .B2(new_n193), .ZN(new_n658));
  OAI21_X1  g472(.A(G472), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n514), .B(KEYINPUT38), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n560), .A2(new_n594), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n641), .A2(new_n598), .A3(new_n662), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n660), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n646), .B(KEYINPUT39), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n410), .A2(new_n665), .ZN(new_n666));
  OR2_X1    g480(.A1(new_n666), .A2(KEYINPUT40), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(KEYINPUT40), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n664), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(new_n194), .ZN(G45));
  INV_X1    g484(.A(new_n646), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n624), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n673), .B1(new_n407), .B2(new_n409), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n311), .A2(new_n674), .A3(new_n649), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G146), .ZN(G48));
  AND2_X1   g490(.A1(new_n390), .A2(new_n396), .ZN(new_n677));
  OAI21_X1  g491(.A(G469), .B1(new_n677), .B2(G902), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n397), .A2(new_n387), .ZN(new_n679));
  INV_X1    g493(.A(new_n403), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(KEYINPUT106), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT106), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n678), .A2(new_n683), .A3(new_n679), .A4(new_n680), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n611), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n311), .A2(new_n686), .A3(new_n464), .A4(new_n626), .ZN(new_n687));
  XOR2_X1   g501(.A(new_n687), .B(KEYINPUT107), .Z(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT41), .B(G113), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G15));
  INV_X1    g504(.A(new_n311), .ZN(new_n691));
  INV_X1    g505(.A(new_n686), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n463), .A2(new_n625), .A3(new_n630), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G116), .ZN(G18));
  NOR2_X1   g510(.A1(new_n640), .A2(new_n596), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G119), .ZN(G21));
  NOR2_X1   g513(.A1(new_n611), .A2(new_n662), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n685), .A2(new_n625), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n276), .B1(new_n193), .B2(new_n306), .ZN(new_n702));
  AOI22_X1  g516(.A1(new_n602), .A2(G472), .B1(new_n187), .B2(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n700), .A2(new_n701), .A3(new_n464), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G122), .ZN(G24));
  NAND4_X1  g519(.A1(new_n686), .A2(new_n641), .A3(new_n672), .A4(new_n703), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G125), .ZN(G27));
  OR2_X1    g521(.A1(new_n292), .A2(KEYINPUT109), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n292), .A2(KEYINPUT109), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n708), .A2(new_n293), .A3(new_n310), .A4(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n515), .A2(new_n597), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT42), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n362), .B1(new_n377), .B2(new_n358), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n398), .B1(new_n387), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n680), .ZN(new_n715));
  NOR4_X1   g529(.A1(new_n711), .A2(new_n712), .A3(new_n673), .A4(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n710), .A2(new_n464), .A3(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n711), .A2(new_n715), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n718), .A2(new_n311), .A3(new_n464), .A4(new_n672), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n719), .A2(new_n720), .A3(new_n712), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n720), .B1(new_n719), .B2(new_n712), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n717), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G131), .ZN(G33));
  INV_X1    g538(.A(new_n647), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n718), .A2(new_n311), .A3(new_n464), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G134), .ZN(G36));
  NAND2_X1  g541(.A1(new_n378), .A2(new_n385), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT45), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n730), .B(G469), .C1(new_n729), .C2(new_n713), .ZN(new_n731));
  INV_X1    g545(.A(new_n389), .ZN(new_n732));
  AOI21_X1  g546(.A(KEYINPUT46), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n733), .B1(new_n387), .B2(new_n397), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n731), .A2(KEYINPUT46), .A3(new_n732), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n403), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n736), .A2(new_n665), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n603), .A2(new_n290), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n561), .A2(new_n623), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT110), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n740), .A2(KEYINPUT43), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n740), .A2(KEYINPUT43), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n739), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n743), .B1(new_n739), .B2(new_n742), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n738), .A2(new_n641), .A3(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT44), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n711), .B1(new_n745), .B2(new_n746), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n737), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G137), .ZN(G39));
  NAND2_X1  g564(.A1(KEYINPUT111), .A2(KEYINPUT47), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n736), .A2(new_n751), .ZN(new_n752));
  XOR2_X1   g566(.A(KEYINPUT111), .B(KEYINPUT47), .Z(new_n753));
  OAI21_X1  g567(.A(new_n752), .B1(new_n736), .B2(new_n753), .ZN(new_n754));
  NOR4_X1   g568(.A1(new_n311), .A2(new_n464), .A3(new_n673), .A4(new_n711), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  OR2_X1    g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  XOR2_X1   g571(.A(KEYINPUT112), .B(G140), .Z(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(G42));
  INV_X1    g573(.A(new_n711), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n760), .A2(KEYINPUT116), .A3(new_n684), .A4(new_n682), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT116), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n762), .B1(new_n711), .B2(new_n685), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n563), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n744), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(KEYINPUT117), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n768), .A2(new_n641), .A3(new_n703), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n656), .A2(new_n464), .A3(new_n659), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n764), .A2(new_n770), .A3(new_n563), .ZN(new_n771));
  AND4_X1   g585(.A1(new_n561), .A2(new_n771), .A3(new_n622), .A4(new_n620), .ZN(new_n772));
  OR3_X1    g586(.A1(new_n769), .A2(KEYINPUT118), .A3(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n678), .A2(new_n679), .A3(new_n404), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n754), .A2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT119), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n754), .A2(KEYINPUT119), .A3(new_n774), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n703), .A2(new_n464), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(new_n766), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n781), .A2(new_n711), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n777), .A2(new_n778), .A3(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(KEYINPUT118), .B1(new_n769), .B2(new_n772), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT50), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n661), .A2(new_n597), .A3(new_n685), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n786), .B1(new_n781), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n780), .A2(KEYINPUT50), .A3(new_n787), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n785), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n773), .A2(new_n783), .A3(new_n784), .A4(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n769), .A2(new_n772), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n789), .A2(new_n790), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n775), .A2(new_n782), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT48), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n710), .A2(new_n464), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n768), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n797), .B1(new_n768), .B2(new_n798), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT120), .ZN(new_n802));
  OAI211_X1 g616(.A(G952), .B(new_n189), .C1(new_n781), .C2(new_n692), .ZN(new_n803));
  INV_X1    g617(.A(new_n624), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n803), .B1(new_n771), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n801), .A2(new_n802), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n802), .B1(new_n801), .B2(new_n805), .ZN(new_n808));
  OAI221_X1 g622(.A(new_n792), .B1(new_n796), .B2(KEYINPUT51), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n598), .B1(new_n512), .B2(new_n513), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n624), .A2(new_n630), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n810), .A2(new_n568), .A3(new_n811), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n630), .A2(KEYINPUT113), .A3(new_n625), .ZN(new_n813));
  AOI22_X1  g627(.A1(new_n812), .A2(KEYINPUT113), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n814), .A2(new_n604), .A3(new_n464), .A4(new_n410), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n311), .B(new_n686), .C1(new_n694), .C2(new_n697), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n815), .A2(new_n816), .A3(new_n704), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n642), .A2(new_n600), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR4_X1   g633(.A1(new_n640), .A2(new_n594), .A3(new_n560), .A4(new_n671), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n820), .A2(new_n410), .A3(new_n760), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n726), .B1(new_n821), .B2(new_n691), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n718), .A2(new_n641), .A3(new_n672), .A4(new_n703), .ZN(new_n823));
  OR2_X1    g637(.A1(new_n823), .A2(KEYINPUT114), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(KEYINPUT114), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n822), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AND4_X1   g640(.A1(new_n688), .A2(new_n723), .A3(new_n819), .A4(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n706), .A2(new_n675), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n829), .B1(new_n653), .B2(new_n651), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n641), .A2(new_n671), .A3(new_n715), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n660), .A2(new_n700), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n828), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n706), .A2(new_n675), .ZN(new_n834));
  AND4_X1   g648(.A1(new_n828), .A2(new_n654), .A3(new_n834), .A4(new_n832), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(KEYINPUT53), .B1(new_n827), .B2(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n723), .A2(new_n826), .A3(new_n688), .A4(new_n819), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n839), .B1(new_n833), .B2(new_n835), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n654), .A2(new_n834), .A3(new_n832), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(KEYINPUT52), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n830), .A2(new_n828), .A3(new_n832), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n842), .A2(new_n843), .A3(KEYINPUT115), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n838), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n837), .B1(new_n845), .B2(KEYINPUT53), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n827), .A2(new_n836), .A3(KEYINPUT53), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n849), .B1(new_n845), .B2(KEYINPUT53), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT54), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  OAI22_X1  g666(.A1(new_n809), .A2(new_n852), .B1(G952), .B2(G953), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n678), .A2(new_n679), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n854), .A2(KEYINPUT49), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n739), .A2(new_n404), .A3(new_n598), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n854), .A2(KEYINPUT49), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OR4_X1    g672(.A1(new_n661), .A2(new_n770), .A3(new_n855), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n853), .A2(new_n859), .ZN(G75));
  XOR2_X1   g674(.A(KEYINPUT121), .B(KEYINPUT55), .Z(new_n861));
  XOR2_X1   g675(.A(new_n504), .B(new_n506), .Z(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n842), .A2(new_n843), .A3(KEYINPUT115), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT115), .B1(new_n842), .B2(new_n843), .ZN(new_n865));
  OAI211_X1 g679(.A(KEYINPUT53), .B(new_n827), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n842), .A2(new_n843), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n867), .B1(new_n868), .B2(new_n838), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n388), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  AOI211_X1 g684(.A(KEYINPUT56), .B(new_n863), .C1(new_n870), .C2(G210), .ZN(new_n871));
  AOI211_X1 g685(.A(new_n867), .B(new_n838), .C1(new_n840), .C2(new_n844), .ZN(new_n872));
  OAI211_X1 g686(.A(G210), .B(G902), .C1(new_n872), .C2(new_n837), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT56), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n862), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n861), .B1(new_n871), .B2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(G210), .ZN(new_n877));
  AOI211_X1 g691(.A(new_n877), .B(new_n388), .C1(new_n866), .C2(new_n869), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n863), .B1(new_n878), .B2(KEYINPUT56), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n873), .A2(new_n874), .A3(new_n862), .ZN(new_n880));
  INV_X1    g694(.A(new_n861), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n189), .A2(G952), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n876), .A2(new_n882), .A3(new_n884), .ZN(G51));
  XNOR2_X1  g699(.A(new_n389), .B(KEYINPUT57), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT122), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n866), .A2(new_n887), .A3(new_n847), .A4(new_n869), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n888), .B1(new_n846), .B2(new_n847), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n887), .B1(new_n846), .B2(new_n847), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n886), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n677), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OR3_X1    g707(.A1(new_n846), .A2(new_n388), .A3(new_n731), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n883), .B1(new_n893), .B2(new_n894), .ZN(G54));
  AND3_X1   g709(.A1(new_n870), .A2(KEYINPUT58), .A3(G475), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n884), .B1(new_n896), .B2(new_n555), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n897), .B1(new_n555), .B2(new_n896), .ZN(G60));
  NOR2_X1   g712(.A1(new_n889), .A2(new_n890), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n618), .A2(new_n619), .ZN(new_n900));
  NAND2_X1  g714(.A1(G478), .A2(G902), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT59), .Z(new_n902));
  NOR3_X1   g716(.A1(new_n899), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n902), .B1(new_n848), .B2(new_n851), .ZN(new_n904));
  INV_X1    g718(.A(new_n900), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n884), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n903), .A2(new_n906), .ZN(G63));
  NAND2_X1  g721(.A1(G217), .A2(G902), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(KEYINPUT123), .Z(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT60), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n846), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n639), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n454), .B1(new_n846), .B2(new_n910), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n912), .A2(new_n884), .A3(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT61), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n912), .A2(KEYINPUT61), .A3(new_n884), .A4(new_n913), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(G66));
  OAI21_X1  g732(.A(G953), .B1(new_n564), .B2(new_n468), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n688), .A2(new_n819), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n919), .B1(new_n920), .B2(G953), .ZN(new_n921));
  INV_X1    g735(.A(new_n504), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n922), .B1(G898), .B2(new_n189), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n921), .B(new_n923), .ZN(G69));
  AOI21_X1  g738(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n749), .A2(new_n830), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT126), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n737), .A2(new_n798), .A3(new_n700), .ZN(new_n928));
  AND4_X1   g742(.A1(new_n723), .A2(new_n757), .A3(new_n726), .A4(new_n928), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n189), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n547), .A2(new_n548), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n269), .B(new_n932), .Z(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n934), .B1(G900), .B2(G953), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n760), .A2(new_n811), .ZN(new_n938));
  OR4_X1    g752(.A1(new_n691), .A2(new_n938), .A3(new_n666), .A4(new_n463), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n749), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT124), .ZN(new_n941));
  INV_X1    g755(.A(new_n757), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n669), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n830), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT62), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(G953), .B1(new_n943), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(KEYINPUT125), .B1(new_n948), .B2(new_n933), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n925), .B1(new_n937), .B2(new_n949), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n948), .A2(new_n933), .ZN(new_n951));
  INV_X1    g765(.A(new_n925), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n951), .A2(KEYINPUT125), .A3(new_n952), .A4(new_n936), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n950), .A2(new_n953), .ZN(G72));
  NAND3_X1  g768(.A1(new_n943), .A2(new_n920), .A3(new_n947), .ZN(new_n955));
  NAND2_X1  g769(.A1(G472), .A2(G902), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT63), .Z(new_n957));
  NAND2_X1  g771(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n883), .B1(new_n958), .B2(new_n657), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n930), .A2(new_n920), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n957), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n961), .A2(new_n300), .A3(new_n296), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n297), .A2(new_n272), .A3(new_n301), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n850), .A2(new_n963), .A3(new_n957), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n959), .A2(new_n962), .A3(new_n964), .ZN(G57));
endmodule


