//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 0 0 0 0 0 1 1 0 1 1 0 0 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:54 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(new_n202), .A2(G50), .ZN(new_n205));
  NAND2_X1  g0005(.A1(G1), .A2(G13), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  NOR3_X1   g0010(.A1(new_n210), .A2(new_n207), .A3(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(KEYINPUT0), .ZN(new_n213));
  OAI22_X1  g0013(.A1(new_n205), .A2(new_n209), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n215));
  INV_X1    g0015(.A(G116), .ZN(new_n216));
  INV_X1    g0016(.A(G270), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n219));
  INV_X1    g0019(.A(G50), .ZN(new_n220));
  INV_X1    g0020(.A(G226), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI211_X1 g0024(.A(new_n218), .B(new_n224), .C1(G97), .C2(G257), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(G1), .B2(G20), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT1), .Z(new_n227));
  AOI211_X1 g0027(.A(new_n214), .B(new_n227), .C1(new_n213), .C2(new_n212), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G68), .B(G77), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G50), .B(G58), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G87), .B(G116), .ZN(new_n240));
  INV_X1    g0040(.A(G107), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(G97), .ZN(new_n242));
  INV_X1    g0042(.A(G97), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G107), .ZN(new_n244));
  NAND3_X1  g0044(.A1(new_n240), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G97), .B(G107), .ZN(new_n246));
  OAI21_X1  g0046(.A(new_n245), .B1(new_n240), .B2(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n239), .B(new_n247), .ZN(G351));
  OAI21_X1  g0048(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n249));
  INV_X1    g0049(.A(G274), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(KEYINPUT72), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT72), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n253), .B1(new_n257), .B2(G33), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(G226), .A3(G1698), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT75), .ZN(new_n260));
  INV_X1    g0060(.A(G1698), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n258), .A2(G223), .A3(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT75), .ZN(new_n263));
  NAND4_X1  g0063(.A1(new_n258), .A2(new_n263), .A3(G226), .A4(G1698), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G87), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n260), .A2(new_n262), .A3(new_n264), .A4(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  INV_X1    g0067(.A(G41), .ZN(new_n268));
  OAI211_X1 g0068(.A(G1), .B(G13), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n251), .B1(new_n266), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n249), .ZN(new_n272));
  INV_X1    g0072(.A(G232), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G169), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n271), .A2(G179), .A3(new_n275), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(KEYINPUT7), .A2(G20), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT73), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n257), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n267), .A2(KEYINPUT3), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n267), .B1(new_n254), .B2(new_n256), .ZN(new_n285));
  NOR3_X1   g0085(.A1(new_n285), .A2(KEYINPUT73), .A3(new_n253), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n280), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(KEYINPUT7), .B1(new_n258), .B2(G20), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n287), .A2(G68), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G58), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n202), .B1(new_n290), .B2(new_n222), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G20), .A2(G33), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n291), .A2(G20), .B1(G159), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n289), .A2(KEYINPUT16), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n206), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n267), .A2(KEYINPUT3), .ZN(new_n297));
  XNOR2_X1  g0097(.A(KEYINPUT72), .B(KEYINPUT3), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n297), .B1(new_n298), .B2(new_n267), .ZN(new_n299));
  OAI21_X1  g0099(.A(KEYINPUT7), .B1(new_n299), .B2(G20), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n252), .A2(G33), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n283), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n280), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n300), .A2(G68), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(new_n293), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT16), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n294), .A2(new_n296), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G13), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n309), .A2(G1), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G20), .ZN(new_n311));
  INV_X1    g0111(.A(new_n296), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n311), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  OR2_X1    g0114(.A1(new_n314), .A2(KEYINPUT67), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n210), .A2(G20), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(KEYINPUT67), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  XNOR2_X1  g0118(.A(KEYINPUT8), .B(G58), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT65), .ZN(new_n320));
  OR3_X1    g0120(.A1(new_n290), .A2(KEYINPUT65), .A3(KEYINPUT8), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  MUX2_X1   g0123(.A(new_n311), .B(new_n318), .S(new_n323), .Z(new_n324));
  AND3_X1   g0124(.A1(new_n308), .A2(KEYINPUT74), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(KEYINPUT74), .B1(new_n308), .B2(new_n324), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n279), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT18), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n308), .A2(new_n324), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(G200), .B2(new_n276), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT77), .ZN(new_n331));
  OR2_X1    g0131(.A1(KEYINPUT76), .A2(G190), .ZN(new_n332));
  NAND2_X1  g0132(.A1(KEYINPUT76), .A2(G190), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n271), .A2(new_n335), .A3(new_n275), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n330), .A2(new_n331), .A3(KEYINPUT17), .A4(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n276), .A2(G200), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n338), .A2(new_n308), .A3(new_n324), .A4(new_n336), .ZN(new_n339));
  OR2_X1    g0139(.A1(new_n331), .A2(KEYINPUT17), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n331), .A2(KEYINPUT17), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT18), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n279), .B(new_n343), .C1(new_n325), .C2(new_n326), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n328), .A2(new_n337), .A3(new_n342), .A4(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n253), .A2(new_n297), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n273), .A2(G1698), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n347), .B(new_n348), .C1(G226), .C2(G1698), .ZN(new_n349));
  NAND2_X1  g0149(.A1(G33), .A2(G97), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT70), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT70), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n349), .A2(new_n353), .A3(new_n350), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n352), .A2(new_n270), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT13), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n272), .A2(new_n223), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n357), .A2(new_n251), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n355), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n356), .B1(new_n355), .B2(new_n358), .ZN(new_n361));
  OAI21_X1  g0161(.A(G169), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(KEYINPUT14), .ZN(new_n363));
  INV_X1    g0163(.A(new_n361), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n359), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT14), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n365), .A2(new_n366), .A3(G169), .ZN(new_n367));
  INV_X1    g0167(.A(G179), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n363), .B(new_n367), .C1(new_n365), .C2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n222), .A2(G20), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n207), .A2(G33), .ZN(new_n371));
  INV_X1    g0171(.A(G77), .ZN(new_n372));
  INV_X1    g0172(.A(new_n292), .ZN(new_n373));
  OAI221_X1 g0173(.A(new_n370), .B1(new_n371), .B2(new_n372), .C1(new_n373), .C2(new_n220), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n296), .ZN(new_n375));
  XOR2_X1   g0175(.A(new_n375), .B(KEYINPUT71), .Z(new_n376));
  OR2_X1    g0176(.A1(new_n376), .A2(KEYINPUT11), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(KEYINPUT11), .ZN(new_n378));
  NOR3_X1   g0178(.A1(new_n370), .A2(G1), .A3(new_n309), .ZN(new_n379));
  OR2_X1    g0179(.A1(new_n379), .A2(KEYINPUT12), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n296), .B1(new_n210), .B2(G20), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n381), .A2(G68), .B1(KEYINPUT12), .B2(new_n379), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n377), .A2(new_n378), .A3(new_n380), .A4(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n369), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n383), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n365), .A2(G200), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n364), .A2(new_n359), .A3(G190), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(G238), .A2(G1698), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n347), .B(new_n389), .C1(new_n273), .C2(G1698), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n390), .B(new_n270), .C1(G107), .C2(new_n347), .ZN(new_n391));
  INV_X1    g0191(.A(new_n251), .ZN(new_n392));
  INV_X1    g0192(.A(G244), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n391), .B(new_n392), .C1(new_n393), .C2(new_n272), .ZN(new_n394));
  OR2_X1    g0194(.A1(new_n394), .A2(G179), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G20), .A2(G77), .ZN(new_n396));
  XNOR2_X1  g0196(.A(KEYINPUT15), .B(G87), .ZN(new_n397));
  XOR2_X1   g0197(.A(new_n292), .B(KEYINPUT69), .Z(new_n398));
  OAI221_X1 g0198(.A(new_n396), .B1(new_n397), .B2(new_n371), .C1(new_n398), .C2(new_n319), .ZN(new_n399));
  INV_X1    g0199(.A(new_n311), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n399), .A2(new_n296), .B1(new_n372), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n381), .A2(G77), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(G169), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n394), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n395), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n346), .A2(new_n384), .A3(new_n388), .A4(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n302), .B1(G222), .B2(new_n261), .ZN(new_n408));
  INV_X1    g0208(.A(G223), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n408), .B1(new_n409), .B2(new_n261), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n410), .B(new_n270), .C1(G77), .C2(new_n347), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n411), .B(new_n392), .C1(new_n221), .C2(new_n272), .ZN(new_n412));
  INV_X1    g0212(.A(G190), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n415));
  INV_X1    g0215(.A(G150), .ZN(new_n416));
  OAI221_X1 g0216(.A(new_n415), .B1(new_n416), .B2(new_n373), .C1(new_n322), .C2(new_n371), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n296), .ZN(new_n418));
  OR2_X1    g0218(.A1(new_n418), .A2(KEYINPUT66), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n418), .A2(KEYINPUT66), .B1(new_n220), .B2(new_n400), .ZN(new_n420));
  OR2_X1    g0220(.A1(new_n318), .A2(new_n220), .ZN(new_n421));
  AND3_X1   g0221(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n414), .B1(new_n422), .B2(KEYINPUT9), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n412), .A2(G200), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT9), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n423), .A2(new_n424), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT10), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT10), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n423), .A2(new_n430), .A3(new_n424), .A4(new_n427), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n412), .A2(new_n404), .ZN(new_n433));
  OR2_X1    g0233(.A1(new_n412), .A2(G179), .ZN(new_n434));
  AND3_X1   g0234(.A1(new_n425), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n394), .A2(G200), .ZN(new_n438));
  INV_X1    g0238(.A(new_n403), .ZN(new_n439));
  OR2_X1    g0239(.A1(new_n394), .A2(new_n413), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n440), .A2(KEYINPUT68), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(KEYINPUT68), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n438), .B(new_n439), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NOR3_X1   g0244(.A1(new_n407), .A2(new_n437), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT90), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n261), .B(new_n283), .C1(new_n298), .C2(new_n267), .ZN(new_n448));
  INV_X1    g0248(.A(G257), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n258), .A2(KEYINPUT90), .A3(G257), .A4(new_n261), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n302), .A2(G303), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n258), .A2(G264), .A3(G1698), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n450), .A2(new_n451), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n270), .ZN(new_n455));
  INV_X1    g0255(.A(G45), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(G1), .ZN(new_n457));
  AND2_X1   g0257(.A1(KEYINPUT5), .A2(G41), .ZN(new_n458));
  NOR2_X1   g0258(.A1(KEYINPUT5), .A2(G41), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OR2_X1    g0260(.A1(new_n460), .A2(new_n250), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n269), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n462), .A2(new_n217), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n455), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G200), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n400), .A2(new_n216), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n312), .B(new_n311), .C1(G1), .C2(new_n267), .ZN(new_n468));
  AOI21_X1  g0268(.A(G20), .B1(G33), .B2(G283), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n469), .B1(G33), .B2(new_n243), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n470), .B(new_n296), .C1(new_n207), .C2(G116), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT20), .ZN(new_n472));
  AND2_X1   g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n471), .A2(new_n472), .ZN(new_n474));
  OAI221_X1 g0274(.A(new_n467), .B1(new_n216), .B2(new_n468), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n463), .B1(new_n454), .B2(new_n270), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n477), .A2(new_n461), .A3(new_n335), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n466), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  NOR3_X1   g0279(.A1(new_n465), .A2(new_n476), .A3(new_n368), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n465), .A2(G169), .A3(new_n475), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(KEYINPUT21), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT21), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n404), .B1(new_n477), .B2(new_n461), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n484), .B1(new_n485), .B2(new_n475), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n479), .B(new_n481), .C1(new_n483), .C2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(G87), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n488), .A2(G20), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n282), .A2(KEYINPUT22), .A3(new_n283), .A4(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(G33), .A2(G116), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n207), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT22), .ZN(new_n494));
  INV_X1    g0294(.A(new_n489), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n494), .B1(new_n302), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT91), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI211_X1 g0299(.A(KEYINPUT91), .B(KEYINPUT23), .C1(new_n207), .C2(G107), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT23), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n207), .A2(G107), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n499), .A2(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n490), .A2(new_n493), .A3(new_n496), .A4(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT24), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n499), .A2(new_n500), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n502), .A2(new_n501), .ZN(new_n507));
  AND3_X1   g0307(.A1(new_n496), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT24), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n508), .A2(new_n509), .A3(new_n493), .A4(new_n490), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n296), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n310), .A2(new_n502), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT25), .ZN(new_n514));
  OAI22_X1  g0314(.A1(new_n468), .A2(new_n241), .B1(KEYINPUT25), .B2(new_n513), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n512), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(G264), .ZN(new_n518));
  OAI21_X1  g0318(.A(KEYINPUT93), .B1(new_n462), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT93), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n460), .A2(new_n520), .A3(G264), .A4(new_n269), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(G294), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n267), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(G250), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n261), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n283), .B(new_n527), .C1(new_n298), .C2(new_n267), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n261), .A2(G257), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n525), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n270), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n522), .B1(new_n531), .B2(KEYINPUT92), .ZN(new_n532));
  INV_X1    g0332(.A(new_n529), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n282), .A2(new_n533), .A3(new_n283), .A4(new_n527), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n269), .B1(new_n534), .B2(new_n525), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT92), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n461), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(G169), .B1(new_n532), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n519), .A2(KEYINPUT94), .A3(new_n521), .ZN(new_n539));
  AND2_X1   g0339(.A1(new_n539), .A2(new_n461), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT94), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n522), .A2(new_n541), .B1(new_n270), .B2(new_n530), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(new_n542), .A3(G179), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n538), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n517), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n515), .B1(new_n511), .B2(new_n296), .ZN(new_n546));
  NOR3_X1   g0346(.A1(new_n532), .A2(new_n537), .A3(G190), .ZN(new_n547));
  AOI21_X1  g0347(.A(G200), .B1(new_n540), .B2(new_n542), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n514), .B(new_n546), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT86), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n223), .A2(new_n261), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n393), .A2(G1698), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NOR3_X1   g0353(.A1(new_n285), .A2(new_n253), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n550), .B1(new_n554), .B2(new_n492), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n283), .B1(new_n298), .B2(new_n267), .ZN(new_n556));
  OAI211_X1 g0356(.A(KEYINPUT86), .B(new_n491), .C1(new_n556), .C2(new_n553), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n555), .A2(new_n270), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n210), .A2(G45), .ZN(new_n559));
  AND2_X1   g0359(.A1(G33), .A2(G41), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n559), .B(G250), .C1(new_n560), .C2(new_n206), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT84), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT84), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n269), .A2(new_n563), .A3(G250), .A4(new_n559), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n457), .A2(G274), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n562), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT85), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT85), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n562), .A2(new_n564), .A3(new_n568), .A4(new_n565), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n558), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G200), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT19), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n350), .B2(G20), .ZN(new_n574));
  NOR2_X1   g0374(.A1(G97), .A2(G107), .ZN(new_n575));
  AND2_X1   g0375(.A1(KEYINPUT88), .A2(G87), .ZN(new_n576));
  NOR2_X1   g0376(.A1(KEYINPUT88), .A2(G87), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n350), .A2(new_n207), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n578), .A2(KEYINPUT19), .A3(new_n579), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n207), .B(new_n283), .C1(new_n298), .C2(new_n267), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n574), .B(new_n580), .C1(new_n581), .C2(new_n222), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n582), .A2(new_n296), .B1(new_n400), .B2(new_n397), .ZN(new_n583));
  OR2_X1    g0383(.A1(new_n468), .A2(new_n488), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n558), .A2(new_n570), .A3(G190), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n572), .A2(new_n583), .A3(new_n584), .A4(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT87), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(new_n571), .B2(G179), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n571), .A2(new_n404), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n468), .A2(new_n397), .ZN(new_n590));
  XNOR2_X1  g0390(.A(new_n590), .B(KEYINPUT89), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n583), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n558), .A2(new_n570), .A3(KEYINPUT87), .A4(new_n368), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n588), .A2(new_n589), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n545), .A2(new_n549), .A3(new_n586), .A4(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n487), .A2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT83), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n393), .A2(G1698), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n283), .B(new_n598), .C1(new_n298), .C2(new_n267), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT80), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n282), .A2(KEYINPUT80), .A3(new_n283), .A4(new_n598), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT4), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(KEYINPUT81), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n598), .A2(KEYINPUT4), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n526), .B2(new_n261), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n607), .A2(new_n347), .B1(G33), .B2(G283), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT81), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n601), .A2(new_n602), .A3(new_n609), .A4(new_n603), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n605), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n270), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n461), .B1(new_n449), .B2(new_n462), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT82), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n612), .A2(KEYINPUT82), .A3(new_n614), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n413), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n400), .A2(new_n243), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(new_n468), .B2(new_n243), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n254), .A2(new_n256), .A3(new_n267), .ZN(new_n622));
  AOI21_X1  g0422(.A(G20), .B1(new_n622), .B2(new_n301), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT7), .ZN(new_n624));
  OAI211_X1 g0424(.A(G107), .B(new_n303), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(KEYINPUT78), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT78), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n300), .A2(new_n627), .A3(G107), .A4(new_n303), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT6), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n246), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n629), .B2(new_n242), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n631), .A2(G20), .B1(G77), .B2(new_n292), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n626), .A2(new_n628), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n296), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(KEYINPUT79), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT79), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n633), .A2(new_n636), .A3(new_n296), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n621), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n615), .A2(G200), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n597), .B1(new_n619), .B2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n617), .A2(new_n404), .A3(new_n618), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n612), .A2(new_n368), .A3(new_n614), .ZN(new_n643));
  INV_X1    g0443(.A(new_n621), .ZN(new_n644));
  INV_X1    g0444(.A(new_n637), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n636), .B1(new_n633), .B2(new_n296), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n642), .A2(new_n643), .A3(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(G200), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n649), .B1(new_n612), .B2(new_n614), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(KEYINPUT82), .B1(new_n612), .B2(new_n614), .ZN(new_n652));
  AOI211_X1 g0452(.A(new_n616), .B(new_n613), .C1(new_n611), .C2(new_n270), .ZN(new_n653));
  OAI21_X1  g0453(.A(G190), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n651), .A2(new_n654), .A3(KEYINPUT83), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n596), .A2(new_n641), .A3(new_n648), .A4(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n446), .A2(new_n656), .ZN(G372));
  NAND2_X1  g0457(.A1(new_n279), .A2(new_n329), .ZN(new_n658));
  XNOR2_X1  g0458(.A(new_n658), .B(new_n343), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n341), .B1(new_n339), .B2(new_n340), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n406), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n369), .A2(new_n383), .B1(new_n388), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n659), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n435), .B1(new_n666), .B2(new_n432), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n594), .A2(new_n586), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT26), .B1(new_n648), .B2(new_n668), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n589), .B(new_n592), .C1(G179), .C2(new_n571), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n652), .A2(new_n653), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n638), .B1(new_n671), .B2(new_n404), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT26), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT95), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n583), .A2(new_n674), .A3(new_n584), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n674), .B1(new_n583), .B2(new_n584), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n572), .B(new_n585), .C1(new_n675), .C2(new_n676), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n670), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n672), .A2(new_n673), .A3(new_n643), .A4(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n669), .A2(new_n670), .A3(new_n679), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n619), .A2(new_n640), .A3(new_n597), .ZN(new_n681));
  AOI21_X1  g0481(.A(KEYINPUT83), .B1(new_n651), .B2(new_n654), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT96), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n532), .A2(new_n537), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n522), .A2(new_n541), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n686), .A2(new_n531), .A3(new_n461), .A4(new_n539), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n685), .A2(new_n413), .B1(new_n687), .B2(new_n649), .ZN(new_n688));
  OAI211_X1 g0488(.A(new_n670), .B(new_n677), .C1(new_n688), .C2(new_n517), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n482), .A2(KEYINPUT21), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n485), .A2(new_n484), .A3(new_n475), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n480), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n689), .B1(new_n692), .B2(new_n545), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n683), .A2(new_n684), .A3(new_n648), .A4(new_n693), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n641), .A2(new_n693), .A3(new_n648), .A4(new_n655), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(KEYINPUT96), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n680), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n667), .B1(new_n446), .B2(new_n697), .ZN(G369));
  INV_X1    g0498(.A(new_n692), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n309), .A2(G20), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n210), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n701), .A2(KEYINPUT27), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(KEYINPUT27), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(G213), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(G343), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n476), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n699), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n487), .B2(new_n708), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G330), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n545), .A2(new_n549), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n517), .A2(new_n706), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n715), .B1(new_n545), .B2(new_n707), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n545), .A2(new_n706), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n692), .A2(new_n706), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n718), .B1(new_n719), .B2(new_n713), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n717), .A2(new_n720), .ZN(G399));
  INV_X1    g0521(.A(KEYINPUT97), .ZN(new_n722));
  INV_X1    g0522(.A(new_n211), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n722), .B1(new_n723), .B2(G41), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n211), .A2(KEYINPUT97), .A3(new_n268), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G1), .ZN(new_n727));
  OR2_X1    g0527(.A1(new_n576), .A2(new_n577), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n728), .A2(new_n216), .A3(new_n575), .ZN(new_n729));
  OAI22_X1  g0529(.A1(new_n727), .A2(new_n729), .B1(new_n205), .B2(new_n726), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT28), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n617), .A2(new_n618), .ZN(new_n732));
  INV_X1    g0532(.A(new_n571), .ZN(new_n733));
  INV_X1    g0533(.A(new_n477), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n543), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n732), .A2(KEYINPUT30), .A3(new_n733), .A4(new_n735), .ZN(new_n736));
  OAI211_X1 g0536(.A(new_n733), .B(new_n735), .C1(new_n652), .C2(new_n653), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT30), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n571), .B(KEYINPUT98), .ZN(new_n740));
  AOI21_X1  g0540(.A(G179), .B1(new_n540), .B2(new_n542), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n740), .A2(new_n465), .A3(new_n615), .A4(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n736), .A2(new_n739), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n706), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n744), .B(KEYINPUT31), .C1(new_n656), .C2(new_n706), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT31), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n743), .A2(new_n746), .A3(new_n706), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(G330), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n680), .ZN(new_n751));
  AND2_X1   g0551(.A1(new_n695), .A2(KEYINPUT96), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n695), .A2(KEYINPUT96), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n707), .ZN(new_n755));
  XOR2_X1   g0555(.A(KEYINPUT99), .B(KEYINPUT29), .Z(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OR3_X1    g0557(.A1(new_n648), .A2(KEYINPUT26), .A3(new_n668), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n670), .A2(new_n677), .ZN(new_n759));
  OAI21_X1  g0559(.A(KEYINPUT26), .B1(new_n648), .B2(new_n759), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n758), .A2(new_n695), .A3(new_n670), .A4(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n761), .A2(KEYINPUT29), .A3(new_n707), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n750), .B1(new_n757), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n731), .B1(new_n763), .B2(G1), .ZN(G364));
  OR2_X1    g0564(.A1(new_n710), .A2(G330), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n700), .B(KEYINPUT100), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n210), .B1(new_n766), .B2(G45), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n726), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n765), .A2(new_n711), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT101), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n207), .A2(G179), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n774), .A2(G190), .A3(G200), .ZN(new_n775));
  INV_X1    g0575(.A(G303), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n207), .A2(new_n368), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G200), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(G190), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G317), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n782), .A2(KEYINPUT33), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(KEYINPUT33), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n781), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n779), .A2(new_n334), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n777), .B(new_n785), .C1(G326), .C2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G190), .A2(G200), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n774), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G329), .ZN(new_n790));
  INV_X1    g0590(.A(G283), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n774), .A2(new_n413), .A3(G200), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n302), .B1(new_n789), .B2(new_n790), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n413), .A2(G179), .A3(G200), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n207), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n793), .B1(G294), .B2(new_n796), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n787), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G311), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n778), .A2(new_n788), .ZN(new_n800));
  INV_X1    g0600(.A(G322), .ZN(new_n801));
  NOR4_X1   g0601(.A1(new_n334), .A2(new_n207), .A3(new_n368), .A4(G200), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT102), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n802), .A2(new_n803), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n798), .B1(new_n799), .B2(new_n800), .C1(new_n801), .C2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n795), .A2(new_n243), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n728), .A2(new_n775), .B1(new_n800), .B2(new_n372), .ZN(new_n809));
  INV_X1    g0609(.A(new_n806), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n809), .B1(new_n810), .B2(G58), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n347), .B1(new_n792), .B2(new_n241), .ZN(new_n812));
  INV_X1    g0612(.A(G159), .ZN(new_n813));
  OAI21_X1  g0613(.A(KEYINPUT32), .B1(new_n789), .B2(new_n813), .ZN(new_n814));
  OR3_X1    g0614(.A1(new_n789), .A2(KEYINPUT32), .A3(new_n813), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n814), .B(new_n815), .C1(new_n781), .C2(new_n222), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n812), .B(new_n816), .C1(G50), .C2(new_n786), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n811), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n807), .B1(new_n808), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n206), .B1(G20), .B2(new_n404), .ZN(new_n820));
  NOR2_X1   g0620(.A1(G13), .A2(G33), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(G20), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n823), .A2(new_n820), .ZN(new_n824));
  INV_X1    g0624(.A(new_n284), .ZN(new_n825));
  INV_X1    g0625(.A(new_n286), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(new_n723), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n239), .A2(G45), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n829), .B(new_n830), .C1(G45), .C2(new_n205), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n347), .A2(G355), .A3(new_n211), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n831), .B(new_n832), .C1(G116), .C2(new_n211), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n819), .A2(new_n820), .B1(new_n824), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n823), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n834), .B1(new_n710), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n773), .B1(new_n771), .B2(new_n836), .ZN(G396));
  NAND2_X1  g0637(.A1(new_n403), .A2(new_n706), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n443), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n406), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n664), .A2(new_n707), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n754), .A2(new_n707), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(KEYINPUT104), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n755), .B(new_n842), .C1(new_n749), .C2(new_n748), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n694), .A2(new_n696), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n706), .B1(new_n847), .B2(new_n751), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n750), .B1(new_n848), .B2(new_n843), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n845), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n846), .A2(new_n845), .A3(new_n849), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n770), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n820), .ZN(new_n854));
  AOI22_X1  g0654(.A1(G137), .A2(new_n786), .B1(new_n780), .B2(G150), .ZN(new_n855));
  INV_X1    g0655(.A(G143), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n855), .B1(new_n813), .B2(new_n800), .C1(new_n806), .C2(new_n856), .ZN(new_n857));
  XOR2_X1   g0657(.A(KEYINPUT103), .B(KEYINPUT34), .Z(new_n858));
  XNOR2_X1  g0658(.A(new_n857), .B(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n792), .A2(new_n222), .ZN(new_n860));
  INV_X1    g0660(.A(G132), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n795), .A2(new_n290), .B1(new_n861), .B2(new_n789), .ZN(new_n862));
  INV_X1    g0662(.A(new_n775), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n860), .B(new_n862), .C1(G50), .C2(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n859), .A2(new_n828), .A3(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n786), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n866), .A2(new_n776), .B1(new_n488), .B2(new_n792), .ZN(new_n867));
  INV_X1    g0667(.A(new_n789), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n347), .B(new_n867), .C1(G311), .C2(new_n868), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n781), .A2(new_n791), .B1(new_n775), .B2(new_n241), .ZN(new_n870));
  INV_X1    g0670(.A(new_n800), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n808), .B(new_n870), .C1(G116), .C2(new_n871), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n869), .B(new_n872), .C1(new_n523), .C2(new_n806), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n854), .B1(new_n865), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(new_n842), .B2(new_n821), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n820), .A2(new_n821), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n372), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n771), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT105), .B1(new_n853), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n852), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n771), .B1(new_n880), .B2(new_n850), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT105), .ZN(new_n882));
  INV_X1    g0682(.A(new_n878), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n879), .A2(new_n884), .ZN(G384));
  INV_X1    g0685(.A(KEYINPUT38), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n294), .A2(new_n296), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT16), .B1(new_n289), .B2(new_n293), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n324), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n704), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT74), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n329), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n308), .A2(KEYINPUT74), .A3(new_n324), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n343), .B1(new_n895), .B2(new_n279), .ZN(new_n896));
  INV_X1    g0696(.A(new_n344), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n891), .B1(new_n898), .B2(new_n662), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n895), .B1(new_n279), .B2(new_n890), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT37), .B1(new_n330), .B2(new_n336), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n279), .A2(new_n889), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(new_n339), .A3(new_n891), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT37), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n886), .B1(new_n899), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n891), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n345), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n902), .A2(new_n905), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n909), .A2(KEYINPUT38), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n907), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n383), .A2(new_n706), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n384), .A2(new_n388), .A3(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n388), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n383), .B(new_n706), .C1(new_n915), .C2(new_n369), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n842), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  AND3_X1   g0717(.A1(new_n745), .A2(new_n747), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n912), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g0719(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT40), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n895), .A2(new_n890), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n922), .B1(new_n659), .B2(new_n662), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n922), .A2(new_n339), .A3(new_n658), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n924), .A2(KEYINPUT37), .B1(new_n901), .B2(new_n900), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n886), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n921), .B1(new_n926), .B2(new_n911), .ZN(new_n927));
  AOI22_X1  g0727(.A1(new_n919), .A2(new_n920), .B1(new_n918), .B2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n748), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n445), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n928), .B(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(G330), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT106), .ZN(new_n933));
  INV_X1    g0733(.A(new_n756), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n445), .B(new_n762), .C1(new_n848), .C2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n667), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n933), .B(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n914), .A2(new_n916), .ZN(new_n938));
  NOR3_X1   g0738(.A1(new_n697), .A2(new_n706), .A3(new_n842), .ZN(new_n939));
  INV_X1    g0739(.A(new_n841), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n912), .B(new_n938), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n659), .A2(new_n890), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n384), .A2(new_n706), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n907), .A2(KEYINPUT39), .A3(new_n911), .ZN(new_n944));
  AND2_X1   g0744(.A1(new_n926), .A2(new_n911), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n943), .B(new_n944), .C1(new_n945), .C2(KEYINPUT39), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n941), .A2(new_n942), .A3(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n937), .B(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n210), .B2(new_n766), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n216), .B1(new_n631), .B2(KEYINPUT35), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n950), .B(new_n208), .C1(KEYINPUT35), .C2(new_n631), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT36), .ZN(new_n952));
  OAI21_X1  g0752(.A(G77), .B1(new_n290), .B2(new_n222), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n205), .A2(new_n953), .B1(G50), .B2(new_n222), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n954), .A2(G1), .A3(new_n309), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n949), .A2(new_n952), .A3(new_n955), .ZN(G367));
  NAND2_X1  g0756(.A1(new_n647), .A2(new_n706), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n641), .A2(new_n648), .A3(new_n655), .A4(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n719), .A2(new_n713), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(KEYINPUT42), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n648), .B1(new_n958), .B2(new_n545), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n707), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT109), .Z(new_n965));
  OR3_X1    g0765(.A1(new_n675), .A2(new_n676), .A3(new_n707), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n678), .A2(new_n966), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n967), .A2(KEYINPUT108), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(KEYINPUT108), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n968), .B(new_n969), .C1(new_n670), .C2(new_n966), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n960), .A2(KEYINPUT42), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n965), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT110), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n971), .B1(new_n965), .B2(new_n972), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n717), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n958), .B1(new_n648), .B2(new_n707), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n974), .A2(new_n979), .A3(new_n980), .A4(new_n977), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n726), .B(KEYINPUT41), .Z(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n959), .B1(new_n716), .B2(new_n719), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(new_n711), .Z(new_n987));
  AND2_X1   g0787(.A1(new_n763), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n980), .A2(new_n720), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT45), .ZN(new_n990));
  OR3_X1    g0790(.A1(new_n980), .A2(KEYINPUT44), .A3(new_n720), .ZN(new_n991));
  OAI21_X1  g0791(.A(KEYINPUT44), .B1(new_n980), .B2(new_n720), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n717), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n979), .B1(new_n990), .B2(new_n993), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n988), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n985), .B1(new_n997), .B2(new_n763), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n982), .B(new_n983), .C1(new_n768), .C2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n829), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n824), .B1(new_n211), .B2(new_n397), .C1(new_n1000), .C2(new_n235), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n290), .A2(new_n775), .B1(new_n800), .B2(new_n220), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(G143), .B2(new_n786), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n792), .A2(new_n372), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(G68), .B2(new_n796), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n302), .B1(new_n780), .B2(G159), .ZN(new_n1006));
  AND3_X1   g0806(.A1(new_n1003), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(G137), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1007), .B1(new_n1008), .B2(new_n789), .C1(new_n416), .C2(new_n806), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n828), .B1(G283), .B2(new_n871), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n810), .A2(G303), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n863), .A2(G116), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT46), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n781), .A2(new_n523), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(new_n1013), .B2(new_n1012), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n866), .A2(new_n799), .B1(new_n241), .B2(new_n795), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n792), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1016), .B1(G97), .B2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1010), .A2(new_n1011), .A3(new_n1015), .A4(new_n1018), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n789), .A2(new_n782), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1009), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT47), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n771), .B1(new_n1022), .B2(new_n820), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1001), .B(new_n1023), .C1(new_n970), .C2(new_n835), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n999), .A2(new_n1024), .ZN(G387));
  AOI22_X1  g0825(.A1(G311), .A2(new_n780), .B1(new_n786), .B2(G322), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n776), .B2(new_n800), .C1(new_n806), .C2(new_n782), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT48), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n791), .B2(new_n795), .C1(new_n523), .C2(new_n775), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT111), .Z(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(KEYINPUT49), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n828), .B1(G326), .B2(new_n868), .ZN(new_n1032));
  AND2_X1   g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1033), .B1(KEYINPUT49), .B2(new_n1030), .C1(new_n216), .C2(new_n792), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n827), .B1(new_n810), .B2(G50), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n781), .A2(new_n322), .B1(new_n243), .B2(new_n792), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n397), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n796), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n863), .A2(G77), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1038), .B(new_n1039), .C1(new_n866), .C2(new_n813), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1036), .B(new_n1040), .C1(G68), .C2(new_n871), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1035), .B(new_n1041), .C1(new_n416), .C2(new_n789), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n854), .B1(new_n1034), .B2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n319), .A2(G50), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT50), .Z(new_n1045));
  NOR2_X1   g0845(.A1(new_n222), .A2(new_n372), .ZN(new_n1046));
  NOR4_X1   g0846(.A1(new_n1045), .A2(G45), .A3(new_n1046), .A4(new_n729), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n829), .B1(new_n232), .B2(new_n456), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n729), .A2(new_n211), .A3(new_n347), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1047), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n211), .A2(G107), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n824), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n716), .B2(new_n835), .ZN(new_n1053));
  NOR3_X1   g0853(.A1(new_n1043), .A2(new_n771), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n768), .B2(new_n987), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n769), .B1(new_n763), .B2(new_n987), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1055), .B1(new_n988), .B2(new_n1056), .ZN(G393));
  OR2_X1    g0857(.A1(new_n995), .A2(KEYINPUT112), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n995), .A2(KEYINPUT112), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n996), .B(KEYINPUT113), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n769), .B(new_n997), .C1(new_n1062), .C2(new_n988), .ZN(new_n1063));
  OAI21_X1  g0863(.A(KEYINPUT114), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1061), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT114), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1065), .A2(new_n1066), .A3(new_n1059), .A4(new_n1058), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1064), .A2(new_n1067), .A3(new_n768), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n829), .A2(new_n247), .B1(G97), .B2(new_n723), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n824), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n806), .A2(new_n799), .B1(new_n782), .B2(new_n866), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT52), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n302), .B1(new_n789), .B2(new_n801), .C1(new_n241), .C2(new_n792), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n781), .A2(new_n776), .B1(new_n216), .B2(new_n795), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n1073), .B(new_n1074), .C1(G283), .C2(new_n863), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1072), .B(new_n1075), .C1(new_n523), .C2(new_n800), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n792), .A2(new_n488), .B1(new_n789), .B2(new_n856), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n222), .B2(new_n775), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n781), .A2(new_n220), .B1(new_n800), .B2(new_n319), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT115), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT51), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n806), .A2(new_n813), .B1(new_n416), .B2(new_n866), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1079), .B(new_n1081), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n1084), .B1(new_n1082), .B2(new_n1083), .C1(new_n372), .C2(new_n795), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1076), .B1(new_n1085), .B2(new_n827), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n771), .B1(new_n1086), .B2(new_n820), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1070), .B(new_n1087), .C1(new_n980), .C2(new_n835), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1063), .A2(new_n1068), .A3(new_n1088), .ZN(G390));
  NAND4_X1  g0889(.A1(new_n745), .A2(new_n747), .A3(G330), .A4(new_n843), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n938), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT118), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n745), .A2(new_n917), .A3(G330), .A4(new_n747), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n844), .A2(new_n841), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1090), .A2(KEYINPUT118), .A3(new_n1091), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n761), .A2(new_n707), .A3(new_n840), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT116), .ZN(new_n1100));
  AND3_X1   g0900(.A1(new_n1099), .A2(new_n1100), .A3(new_n841), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1100), .B1(new_n1099), .B2(new_n841), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1094), .B(new_n1092), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1098), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n445), .A2(new_n929), .A3(G330), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n935), .A2(new_n667), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1104), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT117), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1091), .B1(new_n844), .B2(new_n841), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1109), .B1(new_n1110), .B2(new_n943), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n944), .B1(new_n945), .B2(KEYINPUT39), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n943), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n940), .B1(new_n848), .B2(new_n843), .ZN(new_n1114));
  OAI211_X1 g0914(.A(KEYINPUT117), .B(new_n1113), .C1(new_n1114), .C2(new_n1091), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1111), .A2(new_n1112), .A3(new_n1115), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n945), .A2(new_n943), .ZN(new_n1117));
  OR2_X1    g0917(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1117), .B1(new_n1118), .B2(new_n1091), .ZN(new_n1119));
  AND3_X1   g0919(.A1(new_n1116), .A2(new_n1119), .A3(new_n1094), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1094), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1108), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1094), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1116), .A2(new_n1119), .A3(new_n1094), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1108), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1122), .A2(new_n1128), .A3(new_n769), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n241), .A2(new_n781), .B1(new_n866), .B2(new_n791), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n860), .B(new_n1130), .C1(G97), .C2(new_n871), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n795), .A2(new_n372), .B1(new_n775), .B2(new_n488), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n347), .B(new_n1132), .C1(G294), .C2(new_n868), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1131), .B(new_n1133), .C1(new_n216), .C2(new_n806), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n863), .A2(G150), .ZN(new_n1135));
  XOR2_X1   g0935(.A(new_n1135), .B(KEYINPUT53), .Z(new_n1136));
  AOI22_X1  g0936(.A1(new_n786), .A2(G128), .B1(new_n1017), .B2(G50), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n302), .B1(new_n796), .B2(G159), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(KEYINPUT54), .B(G143), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n781), .A2(new_n1008), .B1(new_n800), .B2(new_n1140), .ZN(new_n1141));
  XOR2_X1   g0941(.A(new_n1141), .B(KEYINPUT119), .Z(new_n1142));
  NAND2_X1  g0942(.A1(new_n868), .A2(G125), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n810), .A2(G132), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1139), .A2(new_n1142), .A3(new_n1143), .A4(new_n1144), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n1134), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n876), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n1146), .A2(new_n854), .B1(new_n323), .B2(new_n1147), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n771), .B(new_n1148), .C1(new_n1112), .C2(new_n821), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1149), .B1(new_n1150), .B2(new_n768), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1129), .A2(new_n1151), .ZN(G378));
  NAND2_X1  g0952(.A1(new_n437), .A2(KEYINPUT55), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT55), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n432), .A2(new_n1154), .A3(new_n436), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n425), .A2(new_n890), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n1156), .B(KEYINPUT56), .Z(new_n1157));
  NAND3_X1  g0957(.A1(new_n1153), .A2(new_n1155), .A3(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1157), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1154), .B1(new_n432), .B2(new_n436), .ZN(new_n1160));
  AOI211_X1 g0960(.A(KEYINPUT55), .B(new_n435), .C1(new_n429), .C2(new_n431), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1159), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n1158), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n928), .B2(G330), .ZN(new_n1164));
  AND3_X1   g0964(.A1(new_n909), .A2(KEYINPUT38), .A3(new_n910), .ZN(new_n1165));
  AOI21_X1  g0965(.A(KEYINPUT38), .B1(new_n909), .B2(new_n910), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n745), .A2(new_n917), .A3(new_n747), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n920), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n927), .A2(new_n918), .ZN(new_n1170));
  AND4_X1   g0970(.A1(G330), .A2(new_n1169), .A3(new_n1170), .A4(new_n1163), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n947), .B1(new_n1164), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1163), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1173), .B1(new_n1174), .B2(new_n749), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n941), .A2(new_n942), .A3(new_n946), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n928), .A2(G330), .A3(new_n1163), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT120), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1172), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n947), .B(KEYINPUT120), .C1(new_n1164), .C2(new_n1171), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NOR3_X1   g0982(.A1(new_n1120), .A2(new_n1121), .A3(new_n1108), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1182), .B1(new_n1183), .B2(new_n1106), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT57), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1128), .A2(new_n1107), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT121), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1172), .A2(new_n1178), .A3(new_n1188), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1175), .A2(new_n1177), .A3(KEYINPUT121), .A4(new_n1176), .ZN(new_n1190));
  AND3_X1   g0990(.A1(new_n1189), .A2(KEYINPUT57), .A3(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n726), .B1(new_n1187), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1186), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1182), .A2(new_n768), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n786), .A2(G125), .B1(new_n871), .B2(G137), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1195), .B1(new_n861), .B2(new_n781), .C1(new_n775), .C2(new_n1140), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(new_n810), .B2(G128), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n416), .B2(new_n795), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1198), .B(KEYINPUT59), .Z(new_n1199));
  AOI21_X1  g0999(.A(G41), .B1(new_n1017), .B2(G159), .ZN(new_n1200));
  AOI21_X1  g1000(.A(G33), .B1(new_n868), .B2(G124), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1017), .A2(G58), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n868), .A2(G283), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1039), .A2(new_n1203), .A3(new_n268), .A4(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n786), .A2(G116), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1206), .B1(new_n397), .B2(new_n800), .C1(new_n781), .C2(new_n243), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1205), .B(new_n1207), .C1(G68), .C2(new_n796), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1208), .B(new_n827), .C1(new_n241), .C2(new_n806), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT58), .ZN(new_n1210));
  AOI21_X1  g1010(.A(G41), .B1(new_n828), .B2(G33), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1202), .B(new_n1210), .C1(G50), .C2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n771), .B1(new_n1212), .B2(new_n820), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1213), .B1(G50), .B2(new_n1147), .C1(new_n1173), .C2(new_n822), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1194), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1193), .A2(new_n1216), .ZN(G375));
  AOI21_X1  g1017(.A(new_n767), .B1(new_n1098), .B2(new_n1103), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT124), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n828), .A2(new_n1203), .ZN(new_n1220));
  XOR2_X1   g1020(.A(new_n1220), .B(KEYINPUT122), .Z(new_n1221));
  AOI22_X1  g1021(.A1(G50), .A2(new_n796), .B1(new_n786), .B2(G132), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(G150), .A2(new_n871), .B1(new_n868), .B2(G128), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1222), .B(new_n1223), .C1(new_n813), .C2(new_n775), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n810), .B2(G137), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1221), .B(new_n1225), .C1(new_n781), .C2(new_n1140), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n216), .A2(new_n781), .B1(new_n866), .B2(new_n523), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n1004), .B(new_n1227), .C1(G107), .C2(new_n871), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1038), .B1(new_n243), .B2(new_n775), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n347), .B(new_n1229), .C1(G303), .C2(new_n868), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1228), .B(new_n1230), .C1(new_n791), .C2(new_n806), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n854), .B1(new_n1226), .B2(new_n1231), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n771), .B(new_n1232), .C1(new_n222), .C2(new_n876), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(KEYINPUT123), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(new_n821), .B2(new_n1091), .ZN(new_n1235));
  NOR3_X1   g1035(.A1(new_n1218), .A2(new_n1219), .A3(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1219), .B1(new_n1218), .B2(new_n1235), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1098), .A2(new_n1106), .A3(new_n1103), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1108), .A2(new_n984), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1239), .A2(new_n1241), .ZN(G381));
  AOI21_X1  g1042(.A(new_n1215), .B1(new_n1186), .B2(new_n1192), .ZN(new_n1243));
  INV_X1    g1043(.A(G378), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(G387), .A2(G381), .ZN(new_n1247));
  NOR4_X1   g1047(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1247), .A2(KEYINPUT125), .A3(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1246), .A2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT125), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1251));
  OR2_X1    g1051(.A1(new_n1250), .A2(new_n1251), .ZN(G407));
  OAI211_X1 g1052(.A(G407), .B(G213), .C1(G343), .C2(new_n1245), .ZN(G409));
  NAND2_X1  g1053(.A1(new_n705), .A2(G213), .ZN(new_n1254));
  AND3_X1   g1054(.A1(new_n1129), .A2(new_n1151), .A3(new_n1214), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1189), .A2(new_n768), .A3(new_n1190), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(new_n1128), .B2(new_n1107), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1256), .B1(new_n1258), .B2(new_n984), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1255), .A2(new_n1259), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1254), .B(new_n1260), .C1(new_n1243), .C2(new_n1244), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT60), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1240), .A2(new_n1262), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1098), .A2(new_n1106), .A3(KEYINPUT60), .A4(new_n1103), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1263), .A2(new_n1108), .A3(new_n769), .A4(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1238), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1265), .B1(new_n1266), .B2(new_n1236), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1267), .A2(G384), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n1239), .A2(new_n1265), .B1(new_n879), .B2(new_n884), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1254), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(G2897), .ZN(new_n1271));
  NOR3_X1   g1071(.A1(new_n1268), .A2(new_n1269), .A3(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT126), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1273), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1239), .A2(new_n879), .A3(new_n884), .A4(new_n1265), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1267), .A2(G384), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1275), .A2(new_n1276), .A3(KEYINPUT126), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1274), .A2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1272), .B1(new_n1278), .B2(new_n1271), .ZN(new_n1279));
  AOI21_X1  g1079(.A(KEYINPUT61), .B1(new_n1261), .B2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1270), .B1(new_n1255), .B2(new_n1259), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1281), .B(new_n1278), .C1(new_n1244), .C2(new_n1243), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(KEYINPUT62), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(G375), .A2(G378), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT62), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1284), .A2(new_n1285), .A3(new_n1281), .A4(new_n1278), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1280), .A2(new_n1283), .A3(new_n1286), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(G393), .B(G396), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n999), .A2(new_n1024), .A3(G390), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(G390), .B1(new_n999), .B2(new_n1024), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1288), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1291), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1288), .A2(KEYINPUT127), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1293), .A2(new_n1289), .A3(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1291), .A2(KEYINPUT127), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1292), .A2(new_n1295), .A3(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1287), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1297), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT63), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1282), .A2(new_n1300), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1284), .A2(KEYINPUT63), .A3(new_n1281), .A4(new_n1278), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1299), .A2(new_n1280), .A3(new_n1301), .A4(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1298), .A2(new_n1303), .ZN(G405));
  NOR2_X1   g1104(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1305), .B1(new_n1246), .B2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1284), .A2(new_n1245), .A3(new_n1278), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1307), .A2(new_n1297), .A3(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1297), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1309), .A2(new_n1310), .ZN(G402));
endmodule


