//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 0 1 0 0 1 1 0 0 1 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 1 0 0 1 0 1 0 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n835, new_n837, new_n838, new_n840, new_n841, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956;
  INV_X1    g000(.A(KEYINPUT14), .ZN(new_n202));
  INV_X1    g001(.A(G29gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n205));
  AOI21_X1  g004(.A(G36gat), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G36gat), .ZN(new_n207));
  NOR3_X1   g006(.A1(new_n202), .A2(new_n207), .A3(G29gat), .ZN(new_n208));
  OR3_X1    g007(.A1(new_n206), .A2(KEYINPUT15), .A3(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT15), .B1(new_n206), .B2(new_n208), .ZN(new_n210));
  XNOR2_X1  g009(.A(G43gat), .B(G50gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n212), .B1(new_n210), .B2(new_n211), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n213), .B(KEYINPUT91), .ZN(new_n214));
  XNOR2_X1  g013(.A(G15gat), .B(G22gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT16), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n215), .B1(new_n216), .B2(G1gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(G1gat), .B2(new_n215), .ZN(new_n218));
  INV_X1    g017(.A(G8gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n218), .B(new_n219), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n214), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(G229gat), .A2(G233gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n214), .A2(KEYINPUT17), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT17), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n213), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(new_n220), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n221), .B(new_n222), .C1(new_n223), .C2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT92), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT18), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT18), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n227), .A2(KEYINPUT92), .A3(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT91), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n213), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n233), .B(new_n220), .ZN(new_n234));
  XOR2_X1   g033(.A(new_n222), .B(KEYINPUT13), .Z(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  OR2_X1    g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n229), .A2(new_n231), .A3(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G113gat), .B(G141gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n239), .B(G197gat), .ZN(new_n240));
  XOR2_X1   g039(.A(KEYINPUT11), .B(G169gat), .Z(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g041(.A(new_n242), .B(KEYINPUT12), .Z(new_n243));
  NAND2_X1  g042(.A1(new_n238), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n243), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n229), .A2(new_n245), .A3(new_n231), .A4(new_n237), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n244), .A2(KEYINPUT93), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT93), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n238), .A2(new_n248), .A3(new_n243), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT94), .ZN(new_n252));
  INV_X1    g051(.A(G64gat), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n252), .B1(new_n253), .B2(G57gat), .ZN(new_n254));
  INV_X1    g053(.A(G57gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n255), .A2(KEYINPUT94), .A3(G64gat), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n254), .B(new_n256), .C1(new_n255), .C2(G64gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(G71gat), .A2(G78gat), .ZN(new_n258));
  OR2_X1    g057(.A1(G71gat), .A2(G78gat), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT9), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(KEYINPUT95), .ZN(new_n263));
  XNOR2_X1  g062(.A(G57gat), .B(G64gat), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n258), .B(new_n259), .C1(new_n264), .C2(new_n260), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT21), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(G231gat), .A2(G233gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G127gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  XOR2_X1   g071(.A(G183gat), .B(G211gat), .Z(new_n273));
  AND2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n220), .B1(new_n266), .B2(new_n267), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT96), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n275), .A2(KEYINPUT96), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n280));
  INV_X1    g079(.A(G155gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  XOR2_X1   g081(.A(new_n279), .B(new_n282), .Z(new_n283));
  NOR2_X1   g082(.A1(new_n272), .A2(new_n273), .ZN(new_n284));
  OR3_X1    g083(.A1(new_n274), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n283), .B1(new_n274), .B2(new_n284), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G190gat), .B(G218gat), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(G85gat), .A2(G92gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n290), .B(KEYINPUT7), .ZN(new_n291));
  NAND2_X1  g090(.A1(G99gat), .A2(G106gat), .ZN(new_n292));
  INV_X1    g091(.A(G85gat), .ZN(new_n293));
  INV_X1    g092(.A(G92gat), .ZN(new_n294));
  AOI22_X1  g093(.A1(KEYINPUT8), .A2(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  XOR2_X1   g095(.A(G99gat), .B(G106gat), .Z(new_n297));
  OR2_X1    g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n296), .A2(new_n297), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n225), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n223), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n300), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n233), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n289), .B1(new_n302), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n233), .A2(new_n224), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n308), .A2(new_n225), .A3(new_n300), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n309), .A2(new_n304), .A3(new_n305), .A4(new_n288), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n307), .A2(new_n310), .A3(KEYINPUT97), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT98), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n307), .A2(new_n310), .A3(KEYINPUT98), .ZN(new_n314));
  XNOR2_X1  g113(.A(G134gat), .B(G162gat), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n311), .A2(new_n312), .A3(new_n317), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n287), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(G230gat), .ZN(new_n323));
  INV_X1    g122(.A(G233gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT100), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n298), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(new_n299), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n296), .A2(new_n326), .A3(new_n297), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n328), .A2(new_n265), .A3(new_n263), .A4(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT10), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n266), .A2(new_n300), .ZN(new_n332));
  AND2_X1   g131(.A1(new_n332), .A2(KEYINPUT99), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(KEYINPUT99), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n330), .B(new_n331), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n303), .A2(KEYINPUT10), .A3(new_n265), .A4(new_n263), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n325), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n325), .ZN(new_n339));
  OR2_X1    g138(.A1(new_n333), .A2(new_n334), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n340), .A2(new_n330), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n338), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(G120gat), .B(G148gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(G176gat), .B(G204gat), .ZN(new_n344));
  XOR2_X1   g143(.A(new_n343), .B(new_n344), .Z(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n342), .A2(new_n346), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n251), .A2(new_n322), .A3(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G78gat), .B(G106gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(KEYINPUT31), .B(G50gat), .ZN(new_n354));
  XOR2_X1   g153(.A(new_n353), .B(new_n354), .Z(new_n355));
  INV_X1    g154(.A(G228gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n356), .A2(new_n324), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G211gat), .B(G218gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(KEYINPUT74), .ZN(new_n360));
  XNOR2_X1  g159(.A(G197gat), .B(G204gat), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT22), .ZN(new_n362));
  INV_X1    g161(.A(G211gat), .ZN(new_n363));
  INV_X1    g162(.A(G218gat), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n360), .A2(new_n366), .ZN(new_n367));
  OR2_X1    g166(.A1(new_n359), .A2(KEYINPUT74), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n359), .A2(KEYINPUT74), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n368), .A2(new_n365), .A3(new_n361), .A4(new_n369), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n367), .A2(KEYINPUT75), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT75), .B1(new_n367), .B2(new_n370), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(KEYINPUT77), .B(G155gat), .ZN(new_n374));
  INV_X1    g173(.A(G162gat), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT2), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OR2_X1    g175(.A1(G141gat), .A2(G148gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n375), .A2(G155gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n281), .A2(G162gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(G141gat), .A2(G148gat), .ZN(new_n380));
  AND4_X1   g179(.A1(new_n377), .A2(new_n378), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT2), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n377), .A2(new_n382), .A3(new_n380), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n378), .A2(new_n379), .ZN(new_n384));
  AOI22_X1  g183(.A1(new_n376), .A2(new_n381), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT3), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT29), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n373), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n367), .A2(new_n370), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT29), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n385), .B1(new_n391), .B2(new_n386), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n358), .B1(new_n388), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NOR3_X1   g193(.A1(new_n388), .A2(new_n358), .A3(new_n392), .ZN(new_n395));
  NOR3_X1   g194(.A1(new_n394), .A2(new_n395), .A3(G22gat), .ZN(new_n396));
  INV_X1    g195(.A(G22gat), .ZN(new_n397));
  INV_X1    g196(.A(new_n395), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n397), .B1(new_n398), .B2(new_n393), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n355), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT81), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT81), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n402), .B(new_n355), .C1(new_n396), .C2(new_n399), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n399), .A2(new_n355), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT82), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n396), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n398), .A2(new_n397), .A3(new_n393), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT82), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n404), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n401), .A2(new_n403), .A3(new_n409), .ZN(new_n410));
  XOR2_X1   g209(.A(G15gat), .B(G43gat), .Z(new_n411));
  XNOR2_X1  g210(.A(G71gat), .B(G99gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(G183gat), .A2(G190gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(G169gat), .A2(G176gat), .ZN(new_n416));
  INV_X1    g215(.A(G169gat), .ZN(new_n417));
  INV_X1    g216(.A(G176gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT26), .ZN(new_n420));
  NOR2_X1   g219(.A1(G169gat), .A2(G176gat), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT26), .ZN(new_n422));
  AND3_X1   g221(.A1(new_n421), .A2(KEYINPUT69), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT69), .B1(new_n421), .B2(new_n422), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n416), .B(new_n420), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT27), .B(G183gat), .ZN(new_n426));
  INV_X1    g225(.A(G190gat), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT67), .ZN(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT67), .B1(new_n426), .B2(new_n427), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n433), .A2(new_n430), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n415), .B(new_n425), .C1(new_n432), .C2(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n415), .A2(KEYINPUT24), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(G183gat), .B(G190gat), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT24), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT66), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT23), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n444), .A2(G169gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n418), .A2(KEYINPUT65), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT65), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(G176gat), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n445), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n416), .A2(KEYINPUT23), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n419), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n442), .B1(new_n443), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n449), .A2(new_n451), .A3(KEYINPUT66), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n437), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n451), .B(KEYINPUT25), .C1(new_n444), .C2(new_n419), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n456), .A2(new_n442), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n435), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  NOR2_X1   g257(.A1(G127gat), .A2(G134gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n271), .A2(KEYINPUT70), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT70), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(G127gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n459), .B1(new_n463), .B2(G134gat), .ZN(new_n464));
  INV_X1    g263(.A(G113gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(G120gat), .ZN(new_n466));
  INV_X1    g265(.A(G120gat), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(G113gat), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT71), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n466), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT1), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n469), .B1(new_n466), .B2(new_n468), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n464), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(KEYINPUT72), .B(G120gat), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n466), .B1(new_n475), .B2(new_n465), .ZN(new_n476));
  INV_X1    g275(.A(new_n459), .ZN(new_n477));
  NAND2_X1  g276(.A1(G127gat), .A2(G134gat), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT1), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n458), .A2(new_n474), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n474), .A2(new_n480), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n435), .B(new_n482), .C1(new_n455), .C2(new_n457), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n481), .A2(new_n483), .A3(G227gat), .A4(G233gat), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT33), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n414), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n481), .A2(new_n483), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT34), .ZN(new_n488));
  NAND2_X1  g287(.A1(G227gat), .A2(G233gat), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n488), .B1(new_n487), .B2(new_n489), .ZN(new_n491));
  NOR3_X1   g290(.A1(new_n486), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n484), .A2(KEYINPUT32), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n486), .B1(new_n490), .B2(new_n491), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n494), .ZN(new_n497));
  INV_X1    g296(.A(new_n495), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n497), .B1(new_n498), .B2(new_n492), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n452), .A2(new_n443), .ZN(new_n501));
  INV_X1    g300(.A(new_n440), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n438), .B1(new_n502), .B2(KEYINPUT24), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n501), .A2(new_n503), .A3(new_n454), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n457), .B1(new_n504), .B2(new_n436), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n425), .A2(new_n415), .ZN(new_n506));
  OR2_X1    g305(.A1(new_n433), .A2(new_n430), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n506), .B1(new_n431), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n390), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(G226gat), .A2(G233gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n510), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n512), .B1(new_n505), .B2(new_n508), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n373), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(KEYINPUT76), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT76), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n458), .A2(new_n516), .A3(new_n512), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n515), .A2(new_n517), .B1(new_n510), .B2(new_n509), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n514), .B1(new_n518), .B2(new_n373), .ZN(new_n519));
  XNOR2_X1  g318(.A(G8gat), .B(G36gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(G64gat), .B(G92gat), .ZN(new_n521));
  XOR2_X1   g320(.A(new_n520), .B(new_n521), .Z(new_n522));
  OR2_X1    g321(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n519), .A2(new_n522), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n523), .A2(KEYINPUT30), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT30), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n519), .A2(new_n526), .A3(new_n522), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  NOR3_X1   g328(.A1(new_n410), .A2(new_n500), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n385), .A2(new_n474), .A3(new_n480), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT4), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n377), .A2(new_n378), .A3(new_n379), .A4(new_n380), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n281), .A2(KEYINPUT77), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n281), .A2(KEYINPUT77), .ZN(new_n536));
  OAI21_X1  g335(.A(G162gat), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n534), .B1(new_n537), .B2(KEYINPUT2), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n383), .A2(new_n384), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT3), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n376), .A2(new_n381), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n542), .A2(new_n386), .A3(new_n539), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n541), .A2(new_n482), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(G225gat), .A2(G233gat), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n385), .A2(new_n474), .A3(KEYINPUT4), .A4(new_n480), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n533), .A2(new_n544), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT78), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT5), .ZN(new_n550));
  INV_X1    g349(.A(new_n385), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n482), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n531), .ZN(new_n553));
  INV_X1    g352(.A(new_n545), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n550), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n549), .A2(new_n555), .ZN(new_n556));
  AND3_X1   g355(.A1(new_n385), .A2(new_n474), .A3(new_n480), .ZN(new_n557));
  AOI22_X1  g356(.A1(new_n474), .A2(new_n480), .B1(new_n542), .B2(new_n539), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n554), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT5), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n560), .A2(new_n548), .A3(new_n547), .ZN(new_n561));
  XOR2_X1   g360(.A(G1gat), .B(G29gat), .Z(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G57gat), .B(G85gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n556), .A2(new_n561), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT84), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT6), .ZN(new_n571));
  INV_X1    g370(.A(new_n561), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n560), .B1(new_n548), .B2(new_n547), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n566), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n556), .A2(KEYINPUT84), .A3(new_n561), .A4(new_n567), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n570), .A2(new_n571), .A3(new_n574), .A4(new_n575), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n568), .A2(new_n571), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(KEYINPUT35), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n530), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n574), .A2(new_n571), .A3(new_n568), .ZN(new_n581));
  OR2_X1    g380(.A1(new_n581), .A2(KEYINPUT80), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n577), .B1(new_n581), .B2(KEYINPUT80), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NOR4_X1   g384(.A1(new_n410), .A2(new_n585), .A3(new_n529), .A4(new_n500), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT35), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n580), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT73), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT36), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(KEYINPUT73), .A2(KEYINPUT36), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n500), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n496), .A2(new_n499), .A3(new_n589), .A4(new_n590), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n401), .A2(new_n403), .A3(new_n409), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n596), .B1(new_n584), .B2(new_n528), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n533), .A2(new_n544), .A3(new_n546), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(new_n554), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n600), .B(KEYINPUT39), .C1(new_n554), .C2(new_n553), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n601), .B(new_n566), .C1(KEYINPUT39), .C2(new_n600), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT40), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n603), .A2(KEYINPUT83), .ZN(new_n604));
  OR2_X1    g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n602), .A2(new_n604), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n605), .A2(new_n570), .A3(new_n575), .A4(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n596), .B1(new_n607), .B2(new_n528), .ZN(new_n608));
  XOR2_X1   g407(.A(KEYINPUT86), .B(KEYINPUT38), .Z(new_n609));
  INV_X1    g408(.A(new_n519), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n522), .B1(new_n610), .B2(KEYINPUT37), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT37), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n519), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n609), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n576), .A2(new_n578), .A3(new_n524), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n511), .A2(KEYINPUT85), .A3(new_n513), .A4(new_n373), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n616), .B1(new_n518), .B2(new_n373), .ZN(new_n617));
  AND3_X1   g416(.A1(new_n511), .A2(new_n513), .A3(new_n373), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n618), .A2(KEYINPUT85), .ZN(new_n619));
  OAI21_X1  g418(.A(KEYINPUT37), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n609), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n522), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n623), .B1(new_n519), .B2(new_n612), .ZN(new_n624));
  AND3_X1   g423(.A1(new_n620), .A2(new_n624), .A3(KEYINPUT87), .ZN(new_n625));
  AOI21_X1  g424(.A(KEYINPUT87), .B1(new_n620), .B2(new_n624), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n615), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n614), .B1(new_n627), .B2(KEYINPUT88), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n576), .A2(new_n578), .A3(new_n524), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n620), .A2(new_n624), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT87), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n620), .A2(new_n624), .A3(KEYINPUT87), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n629), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT88), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n608), .B1(new_n628), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT89), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n598), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AOI211_X1 g438(.A(KEYINPUT89), .B(new_n608), .C1(new_n628), .C2(new_n636), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n588), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT90), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n528), .A2(new_n607), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n410), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n614), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n646), .B1(new_n634), .B2(new_n635), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n627), .A2(KEYINPUT88), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(KEYINPUT89), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n637), .A2(new_n638), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n650), .A2(new_n651), .A3(new_n598), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n652), .A2(KEYINPUT90), .A3(new_n588), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n352), .B1(new_n643), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(new_n585), .ZN(new_n655));
  XNOR2_X1  g454(.A(KEYINPUT101), .B(G1gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(G1324gat));
  INV_X1    g456(.A(new_n654), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n216), .A2(new_n219), .ZN(new_n659));
  NOR2_X1   g458(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n660));
  NOR4_X1   g459(.A1(new_n658), .A2(new_n528), .A3(new_n659), .A4(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n219), .B1(new_n654), .B2(new_n529), .ZN(new_n662));
  OAI21_X1  g461(.A(KEYINPUT42), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n663), .B1(KEYINPUT42), .B2(new_n661), .ZN(G1325gat));
  XNOR2_X1  g463(.A(new_n595), .B(KEYINPUT102), .ZN(new_n665));
  OAI21_X1  g464(.A(G15gat), .B1(new_n658), .B2(new_n665), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n500), .A2(G15gat), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n666), .B1(new_n658), .B2(new_n667), .ZN(G1326gat));
  NAND2_X1  g467(.A1(new_n654), .A2(new_n410), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT103), .ZN(new_n670));
  XNOR2_X1  g469(.A(KEYINPUT43), .B(G22gat), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n670), .B(new_n671), .Z(G1327gat));
  INV_X1    g471(.A(KEYINPUT45), .ZN(new_n673));
  INV_X1    g472(.A(new_n321), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n674), .B1(new_n643), .B2(new_n653), .ZN(new_n675));
  INV_X1    g474(.A(new_n287), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n250), .A2(new_n676), .A3(new_n350), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n585), .A2(new_n203), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n673), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OR3_X1    g479(.A1(new_n678), .A2(new_n673), .A3(new_n679), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT105), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT104), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n319), .A2(new_n684), .A3(new_n320), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n684), .B1(new_n319), .B2(new_n320), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n641), .A2(new_n683), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n689), .B1(new_n675), .B2(new_n683), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(new_n677), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n682), .B1(new_n691), .B2(new_n584), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(G29gat), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n691), .A2(new_n682), .A3(new_n584), .ZN(new_n694));
  OAI211_X1 g493(.A(new_n680), .B(new_n681), .C1(new_n693), .C2(new_n694), .ZN(G1328gat));
  OAI21_X1  g494(.A(G36gat), .B1(new_n691), .B2(new_n528), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n529), .A2(new_n207), .ZN(new_n697));
  OAI21_X1  g496(.A(KEYINPUT46), .B1(new_n678), .B2(new_n697), .ZN(new_n698));
  OR3_X1    g497(.A1(new_n678), .A2(KEYINPUT46), .A3(new_n697), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n696), .A2(new_n698), .A3(new_n699), .ZN(G1329gat));
  NAND3_X1  g499(.A1(new_n690), .A2(new_n595), .A3(new_n677), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n701), .A2(G43gat), .ZN(new_n702));
  INV_X1    g501(.A(G43gat), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n496), .A2(new_n703), .A3(new_n499), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT47), .B1(new_n678), .B2(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n678), .A2(new_n704), .ZN(new_n706));
  INV_X1    g505(.A(new_n665), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n690), .A2(new_n707), .A3(new_n677), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n706), .B1(new_n708), .B2(G43gat), .ZN(new_n709));
  OAI22_X1  g508(.A1(new_n702), .A2(new_n705), .B1(new_n709), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g509(.A1(new_n410), .A2(G50gat), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n678), .A2(new_n596), .ZN(new_n712));
  OAI22_X1  g511(.A1(new_n691), .A2(new_n711), .B1(new_n712), .B2(G50gat), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT48), .ZN(G1331gat));
  AND4_X1   g513(.A1(new_n641), .A2(new_n250), .A3(new_n350), .A4(new_n322), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n584), .B(KEYINPUT106), .Z(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g517(.A1(new_n715), .A2(new_n529), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n720));
  XOR2_X1   g519(.A(KEYINPUT49), .B(G64gat), .Z(new_n721));
  OAI21_X1  g520(.A(new_n720), .B1(new_n719), .B2(new_n721), .ZN(G1333gat));
  NAND2_X1  g521(.A1(new_n715), .A2(new_n707), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n500), .A2(G71gat), .ZN(new_n724));
  AOI22_X1  g523(.A1(new_n723), .A2(G71gat), .B1(new_n715), .B2(new_n724), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g525(.A1(new_n715), .A2(new_n410), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g527(.A1(new_n251), .A2(new_n676), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n350), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n641), .A2(new_n642), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT90), .B1(new_n652), .B2(new_n588), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n321), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(KEYINPUT44), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n730), .B1(new_n734), .B2(new_n689), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(G85gat), .B1(new_n736), .B2(new_n584), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n729), .A2(new_n321), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n641), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT51), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT51), .B1(new_n641), .B2(new_n739), .ZN(new_n743));
  OR2_X1    g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n350), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n585), .A2(new_n293), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n737), .B1(new_n745), .B2(new_n746), .ZN(G1336gat));
  INV_X1    g546(.A(new_n730), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n643), .A2(new_n653), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n683), .B1(new_n749), .B2(new_n321), .ZN(new_n750));
  INV_X1    g549(.A(new_n689), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n529), .B(new_n748), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT108), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n690), .A2(KEYINPUT108), .A3(new_n529), .A4(new_n748), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n754), .A2(G92gat), .A3(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n744), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n350), .A2(new_n294), .A3(new_n529), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n759), .A2(KEYINPUT52), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n294), .B1(new_n735), .B2(new_n529), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n758), .B(KEYINPUT107), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n757), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(KEYINPUT52), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n761), .A2(new_n765), .ZN(G1337gat));
  OAI21_X1  g565(.A(G99gat), .B1(new_n736), .B2(new_n665), .ZN(new_n767));
  OR2_X1    g566(.A1(new_n500), .A2(G99gat), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n767), .B1(new_n745), .B2(new_n768), .ZN(G1338gat));
  INV_X1    g568(.A(KEYINPUT53), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n596), .A2(G106gat), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n350), .B(new_n771), .C1(new_n742), .C2(new_n743), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n773), .B1(new_n735), .B2(new_n410), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n690), .A2(new_n773), .A3(new_n410), .A4(new_n748), .ZN(new_n775));
  XNOR2_X1  g574(.A(KEYINPUT109), .B(G106gat), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n770), .B(new_n772), .C1(new_n774), .C2(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n776), .B1(new_n735), .B2(new_n410), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n772), .B(KEYINPUT110), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT53), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n779), .A2(new_n782), .ZN(G1339gat));
  AND3_X1   g582(.A1(new_n335), .A2(new_n325), .A3(new_n336), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT54), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n784), .A2(new_n337), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n345), .B1(new_n337), .B2(new_n785), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT113), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT113), .ZN(new_n789));
  AOI211_X1 g588(.A(KEYINPUT54), .B(new_n325), .C1(new_n335), .C2(new_n336), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n789), .B1(new_n790), .B2(new_n345), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n786), .B1(new_n788), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n347), .B1(new_n792), .B2(KEYINPUT55), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n787), .A2(KEYINPUT113), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n790), .A2(new_n789), .A3(new_n345), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n794), .B1(new_n797), .B2(new_n786), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n793), .A2(new_n798), .A3(new_n247), .A4(new_n249), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n234), .A2(new_n236), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n308), .A2(new_n220), .A3(new_n225), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n222), .B1(new_n801), .B2(new_n221), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n242), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  OR2_X1    g602(.A1(new_n803), .A2(KEYINPUT114), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(KEYINPUT114), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n804), .A2(new_n246), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n350), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n688), .B1(new_n799), .B2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n687), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n685), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n806), .A2(new_n793), .A3(new_n798), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n287), .B1(new_n808), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n322), .A2(new_n250), .A3(new_n351), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(KEYINPUT112), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT112), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n322), .A2(new_n250), .A3(new_n816), .A4(new_n351), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n813), .A2(new_n818), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n819), .A2(new_n716), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n820), .A2(new_n530), .ZN(new_n821));
  AOI21_X1  g620(.A(G113gat), .B1(new_n821), .B2(new_n251), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n819), .A2(new_n596), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(KEYINPUT115), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT115), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n819), .A2(new_n825), .A3(new_n596), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n529), .A2(new_n500), .A3(new_n584), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n250), .A2(new_n465), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n822), .B1(new_n830), .B2(new_n831), .ZN(G1340gat));
  OAI21_X1  g631(.A(G120gat), .B1(new_n829), .B2(new_n351), .ZN(new_n833));
  INV_X1    g632(.A(new_n475), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n821), .A2(new_n834), .A3(new_n350), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(G1341gat));
  OAI21_X1  g635(.A(new_n463), .B1(new_n829), .B2(new_n287), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n821), .A2(new_n460), .A3(new_n462), .A4(new_n676), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(G1342gat));
  INV_X1    g638(.A(G134gat), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n821), .A2(new_n840), .A3(new_n321), .ZN(new_n841));
  XOR2_X1   g640(.A(new_n841), .B(KEYINPUT56), .Z(new_n842));
  OAI21_X1  g641(.A(G134gat), .B1(new_n829), .B2(new_n674), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(G1343gat));
  NOR3_X1   g643(.A1(new_n595), .A2(new_n584), .A3(new_n529), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT57), .B1(new_n819), .B2(new_n410), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n410), .A2(KEYINPUT57), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n321), .B1(new_n799), .B2(new_n807), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n287), .B1(new_n848), .B2(new_n812), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n847), .B1(new_n849), .B2(new_n818), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n251), .B(new_n845), .C1(new_n846), .C2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(G141gat), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n707), .A2(new_n529), .A3(new_n596), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n250), .A2(G141gat), .ZN(new_n854));
  AND4_X1   g653(.A1(new_n716), .A2(new_n819), .A3(new_n853), .A4(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(KEYINPUT117), .ZN(new_n858));
  AOI21_X1  g657(.A(KEYINPUT116), .B1(new_n851), .B2(G141gat), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT58), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT117), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n852), .A2(new_n856), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n858), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n862), .B1(new_n852), .B2(new_n856), .ZN(new_n865));
  AOI211_X1 g664(.A(KEYINPUT117), .B(new_n855), .C1(new_n851), .C2(G141gat), .ZN(new_n866));
  OAI22_X1  g665(.A1(new_n865), .A2(new_n866), .B1(new_n860), .B2(new_n859), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n864), .A2(new_n867), .ZN(G1344gat));
  AND2_X1   g667(.A1(new_n820), .A2(new_n853), .ZN(new_n869));
  INV_X1    g668(.A(G148gat), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n869), .A2(new_n870), .A3(new_n350), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n845), .B1(new_n846), .B2(new_n850), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n872), .A2(new_n351), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT59), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n873), .A2(new_n874), .A3(G148gat), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n819), .A2(KEYINPUT57), .A3(new_n410), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n811), .A2(new_n674), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n287), .B1(new_n848), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n596), .B1(new_n878), .B2(new_n814), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n876), .B1(new_n879), .B2(KEYINPUT57), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(new_n350), .A3(new_n845), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n874), .B1(new_n881), .B2(G148gat), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n871), .B1(new_n875), .B2(new_n882), .ZN(G1345gat));
  OAI22_X1  g682(.A1(new_n872), .A2(new_n287), .B1(new_n535), .B2(new_n536), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n869), .A2(new_n374), .A3(new_n676), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(G1346gat));
  NAND3_X1  g685(.A1(new_n869), .A2(new_n375), .A3(new_n321), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(KEYINPUT118), .ZN(new_n888));
  OAI21_X1  g687(.A(G162gat), .B1(new_n872), .B2(new_n810), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(G1347gat));
  NOR2_X1   g689(.A1(new_n716), .A2(new_n528), .ZN(new_n891));
  XOR2_X1   g690(.A(new_n891), .B(KEYINPUT119), .Z(new_n892));
  NAND3_X1  g691(.A1(new_n892), .A2(new_n496), .A3(new_n499), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n893), .B1(new_n824), .B2(new_n826), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(G169gat), .A3(new_n251), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n585), .B1(new_n813), .B2(new_n818), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n410), .A2(new_n500), .A3(new_n528), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n417), .B1(new_n898), .B2(new_n250), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n895), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT120), .ZN(G1348gat));
  INV_X1    g700(.A(new_n898), .ZN(new_n902));
  AOI21_X1  g701(.A(G176gat), .B1(new_n902), .B2(new_n350), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n351), .B1(new_n446), .B2(new_n448), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n903), .B1(new_n894), .B2(new_n904), .ZN(G1349gat));
  NAND2_X1  g704(.A1(new_n894), .A2(new_n676), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(G183gat), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n902), .A2(new_n426), .A3(new_n676), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT60), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT60), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n907), .A2(new_n911), .A3(new_n908), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(G1350gat));
  AOI21_X1  g712(.A(new_n427), .B1(new_n894), .B2(new_n321), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n914), .A2(KEYINPUT61), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(KEYINPUT61), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n902), .A2(new_n427), .A3(new_n688), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT121), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n915), .A2(new_n916), .A3(new_n918), .ZN(G1351gat));
  INV_X1    g718(.A(G197gat), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT123), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n665), .A2(new_n529), .A3(new_n410), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT122), .ZN(new_n923));
  INV_X1    g722(.A(new_n896), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n921), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n922), .B(new_n926), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n927), .A2(KEYINPUT123), .A3(new_n896), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n920), .B1(new_n929), .B2(new_n250), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n892), .A2(new_n665), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT124), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n931), .B(new_n932), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n933), .A2(G197gat), .A3(new_n251), .A4(new_n880), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n930), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(KEYINPUT125), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT125), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n930), .A2(new_n934), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(G1352gat));
  INV_X1    g738(.A(G204gat), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n933), .A2(new_n350), .A3(new_n880), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n940), .B1(new_n941), .B2(KEYINPUT126), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n942), .B1(KEYINPUT126), .B2(new_n941), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n927), .A2(new_n940), .A3(new_n350), .A4(new_n896), .ZN(new_n944));
  XOR2_X1   g743(.A(new_n944), .B(KEYINPUT62), .Z(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(new_n945), .ZN(G1353gat));
  NAND3_X1  g745(.A1(new_n933), .A2(new_n676), .A3(new_n880), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT63), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n948), .A2(KEYINPUT127), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n363), .B1(KEYINPUT127), .B2(new_n948), .ZN(new_n950));
  AND3_X1   g749(.A1(new_n947), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n949), .B1(new_n947), .B2(new_n950), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n676), .A2(new_n363), .ZN(new_n953));
  OAI22_X1  g752(.A1(new_n951), .A2(new_n952), .B1(new_n929), .B2(new_n953), .ZN(G1354gat));
  AND3_X1   g753(.A1(new_n933), .A2(new_n321), .A3(new_n880), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n688), .A2(new_n364), .ZN(new_n956));
  OAI22_X1  g755(.A1(new_n955), .A2(new_n364), .B1(new_n929), .B2(new_n956), .ZN(G1355gat));
endmodule


