//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 0 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0 1 0 0 1 1 0 1 1 0 1 0 1 1 1 1 0 1 0 0 0 1 0 1 1 1 0 0 0 1 0 0 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n818, new_n819, new_n820,
    new_n822, new_n823, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940;
  XNOR2_X1  g000(.A(G15gat), .B(G43gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT73), .ZN(new_n203));
  XNOR2_X1  g002(.A(G71gat), .B(G99gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G169gat), .ZN(new_n206));
  INV_X1    g005(.A(G176gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT23), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n209), .B1(G169gat), .B2(G176gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  AND3_X1   g010(.A1(new_n208), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  NAND3_X1  g011(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT66), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT24), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G183gat), .ZN(new_n219));
  INV_X1    g018(.A(G190gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n215), .A2(new_n218), .A3(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n213), .A2(new_n214), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n212), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n221), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n219), .A2(new_n220), .A3(KEYINPUT65), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n226), .A2(new_n213), .A3(new_n218), .A4(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n208), .A2(new_n210), .A3(new_n211), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n229), .A2(KEYINPUT25), .ZN(new_n230));
  AOI22_X1  g029(.A1(new_n224), .A2(KEYINPUT25), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT69), .ZN(new_n232));
  AOI22_X1  g031(.A1(new_n232), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT26), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n234), .A2(new_n206), .A3(new_n207), .A4(KEYINPUT69), .ZN(new_n235));
  AOI22_X1  g034(.A1(new_n233), .A2(new_n235), .B1(G183gat), .B2(G190gat), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT67), .ZN(new_n237));
  OAI21_X1  g036(.A(KEYINPUT27), .B1(new_n237), .B2(new_n219), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT27), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n239), .A2(KEYINPUT67), .A3(G183gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n220), .A3(new_n240), .ZN(new_n241));
  XOR2_X1   g040(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n242));
  AND2_X1   g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT27), .B(G183gat), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n220), .A2(KEYINPUT28), .ZN(new_n245));
  AND2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n236), .B1(new_n243), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G113gat), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT70), .B1(new_n249), .B2(G120gat), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT71), .ZN(new_n251));
  INV_X1    g050(.A(G120gat), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n251), .B1(new_n252), .B2(G113gat), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n254), .A2(new_n252), .A3(G113gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n249), .A2(KEYINPUT71), .A3(G120gat), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n250), .A2(new_n253), .A3(new_n255), .A4(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(G134gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(G127gat), .ZN(new_n259));
  INV_X1    g058(.A(G127gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G134gat), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT1), .ZN(new_n262));
  AND3_X1   g061(.A1(new_n259), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT72), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n257), .A2(KEYINPUT72), .A3(new_n263), .ZN(new_n267));
  XOR2_X1   g066(.A(G113gat), .B(G120gat), .Z(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(new_n262), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n259), .A2(new_n261), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n266), .A2(new_n267), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n248), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n269), .A2(new_n270), .ZN(new_n273));
  AND3_X1   g072(.A1(new_n257), .A2(KEYINPUT72), .A3(new_n263), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT72), .B1(new_n257), .B2(new_n263), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n276), .A2(new_n231), .A3(new_n247), .ZN(new_n277));
  INV_X1    g076(.A(G227gat), .ZN(new_n278));
  INV_X1    g077(.A(G233gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n280), .B(KEYINPUT64), .Z(new_n281));
  NAND3_X1  g080(.A1(new_n272), .A2(new_n277), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT33), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n205), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(KEYINPUT32), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n272), .A2(new_n277), .ZN(new_n287));
  INV_X1    g086(.A(new_n280), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n281), .A2(KEYINPUT34), .ZN(new_n290));
  AOI22_X1  g089(.A1(new_n289), .A2(KEYINPUT34), .B1(new_n287), .B2(new_n290), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n282), .B(KEYINPUT32), .C1(new_n283), .C2(new_n205), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n286), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n291), .B1(new_n286), .B2(new_n292), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT3), .ZN(new_n296));
  INV_X1    g095(.A(G197gat), .ZN(new_n297));
  INV_X1    g096(.A(G204gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(G197gat), .A2(G204gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(G211gat), .A2(G218gat), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n301), .B1(KEYINPUT22), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT82), .ZN(new_n305));
  XNOR2_X1  g104(.A(G211gat), .B(G218gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n304), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT22), .ZN(new_n309));
  AOI22_X1  g108(.A1(new_n299), .A2(new_n300), .B1(new_n309), .B2(new_n302), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(new_n306), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT82), .B1(new_n310), .B2(new_n306), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n308), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n296), .B1(new_n313), .B2(KEYINPUT29), .ZN(new_n314));
  INV_X1    g113(.A(G162gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G155gat), .ZN(new_n316));
  INV_X1    g115(.A(G155gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G162gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  OR2_X1    g118(.A1(KEYINPUT76), .A2(G148gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(KEYINPUT76), .A2(G148gat), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n320), .A2(G141gat), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(G141gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G148gat), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n319), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  AND2_X1   g124(.A1(KEYINPUT77), .A2(G155gat), .ZN(new_n326));
  NOR2_X1   g125(.A1(KEYINPUT77), .A2(G155gat), .ZN(new_n327));
  OAI21_X1  g126(.A(G162gat), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT2), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT2), .ZN(new_n331));
  INV_X1    g130(.A(new_n324), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n323), .A2(G148gat), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(new_n319), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT78), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n325), .A2(new_n329), .B1(new_n319), .B2(new_n334), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT78), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n314), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT83), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n304), .A2(new_n307), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n344), .A2(KEYINPUT75), .A3(new_n311), .ZN(new_n345));
  OR3_X1    g144(.A1(new_n310), .A2(KEYINPUT75), .A3(new_n306), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n336), .A2(KEYINPUT3), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n343), .B(new_n347), .C1(new_n348), .C2(KEYINPUT29), .ZN(new_n349));
  AND2_X1   g148(.A1(new_n345), .A2(new_n346), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT29), .B1(new_n339), .B2(new_n296), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT83), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n342), .A2(new_n349), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(G228gat), .A2(G233gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(KEYINPUT81), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  AND2_X1   g155(.A1(G228gat), .A2(G233gat), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT29), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT3), .B1(new_n350), .B2(new_n358), .ZN(new_n359));
  OAI221_X1 g158(.A(new_n357), .B1(new_n350), .B2(new_n351), .C1(new_n359), .C2(new_n339), .ZN(new_n360));
  XNOR2_X1  g159(.A(G78gat), .B(G106gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(KEYINPUT31), .B(G50gat), .ZN(new_n362));
  XOR2_X1   g161(.A(new_n361), .B(new_n362), .Z(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n356), .A2(new_n360), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n364), .B1(new_n356), .B2(new_n360), .ZN(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT84), .B(G22gat), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NOR3_X1   g168(.A1(new_n366), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n356), .A2(new_n360), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(new_n363), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n368), .B1(new_n372), .B2(new_n365), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n295), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G8gat), .B(G36gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(G64gat), .B(G92gat), .ZN(new_n376));
  XOR2_X1   g175(.A(new_n375), .B(new_n376), .Z(new_n377));
  NAND2_X1  g176(.A1(new_n224), .A2(KEYINPUT25), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n230), .A2(new_n228), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n233), .A2(new_n235), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(new_n216), .ZN(new_n382));
  AOI22_X1  g181(.A1(new_n241), .A2(new_n242), .B1(new_n244), .B2(new_n245), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n358), .B1(new_n380), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G226gat), .A2(G233gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n386), .B1(new_n231), .B2(new_n247), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n347), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n386), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n391), .B1(new_n248), .B2(new_n358), .ZN(new_n392));
  NOR3_X1   g191(.A1(new_n392), .A2(new_n350), .A3(new_n388), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n377), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n387), .A2(new_n347), .A3(new_n389), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n350), .B1(new_n392), .B2(new_n388), .ZN(new_n396));
  INV_X1    g195(.A(new_n377), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n394), .A2(KEYINPUT30), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT30), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n400), .B(new_n377), .C1(new_n390), .C2(new_n393), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  XOR2_X1   g201(.A(G1gat), .B(G29gat), .Z(new_n403));
  XNOR2_X1  g202(.A(new_n403), .B(KEYINPUT0), .ZN(new_n404));
  XNOR2_X1  g203(.A(G57gat), .B(G85gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n404), .B(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT6), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n406), .A2(KEYINPUT6), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n338), .A2(new_n271), .A3(KEYINPUT4), .A4(new_n340), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n339), .B(new_n273), .C1(new_n275), .C2(new_n274), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT4), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n336), .A2(KEYINPUT3), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n339), .A2(new_n296), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n415), .A2(new_n276), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(G225gat), .A2(G233gat), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n411), .A2(new_n414), .A3(new_n417), .A4(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n276), .A2(new_n336), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n412), .ZN(new_n421));
  INV_X1    g220(.A(new_n418), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT79), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT79), .ZN(new_n424));
  AOI211_X1 g223(.A(new_n424), .B(new_n418), .C1(new_n420), .C2(new_n412), .ZN(new_n425));
  OAI211_X1 g224(.A(KEYINPUT5), .B(new_n419), .C1(new_n423), .C2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n412), .A2(KEYINPUT4), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n338), .A2(new_n271), .A3(new_n340), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n427), .B1(new_n428), .B2(KEYINPUT4), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT5), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n429), .A2(new_n430), .A3(new_n418), .A4(new_n417), .ZN(new_n431));
  AOI211_X1 g230(.A(new_n409), .B(new_n410), .C1(new_n426), .C2(new_n431), .ZN(new_n432));
  AND4_X1   g231(.A1(new_n408), .A2(new_n426), .A3(new_n431), .A4(new_n407), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n402), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT80), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n426), .A2(new_n431), .ZN(new_n437));
  INV_X1    g236(.A(new_n409), .ZN(new_n438));
  INV_X1    g237(.A(new_n410), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n426), .A2(new_n408), .A3(new_n431), .A4(new_n407), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n442), .A2(KEYINPUT80), .A3(new_n402), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n374), .B1(new_n436), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT35), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT90), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n286), .A2(new_n292), .ZN(new_n447));
  INV_X1    g246(.A(new_n291), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n286), .A2(new_n291), .A3(new_n292), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n373), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n372), .A2(new_n368), .A3(new_n365), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AOI221_X4 g253(.A(new_n435), .B1(new_n399), .B2(new_n401), .C1(new_n440), .C2(new_n441), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT80), .B1(new_n442), .B2(new_n402), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT90), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n457), .A2(new_n458), .A3(KEYINPUT35), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT88), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n434), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n442), .A2(KEYINPUT88), .A3(new_n402), .ZN(new_n462));
  XOR2_X1   g261(.A(KEYINPUT89), .B(KEYINPUT35), .Z(new_n463));
  NAND4_X1  g262(.A1(new_n454), .A2(new_n461), .A3(new_n462), .A4(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n446), .A2(new_n459), .A3(new_n464), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n370), .A2(new_n373), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n436), .A2(new_n466), .A3(new_n443), .ZN(new_n467));
  AND2_X1   g266(.A1(KEYINPUT74), .A2(KEYINPUT36), .ZN(new_n468));
  OR2_X1    g267(.A1(new_n295), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g268(.A1(KEYINPUT74), .A2(KEYINPUT36), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n295), .B1(new_n470), .B2(new_n468), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n442), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n397), .A2(KEYINPUT37), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n398), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n395), .A2(new_n396), .A3(KEYINPUT37), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT86), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT38), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT86), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n395), .A2(new_n396), .A3(new_n479), .A4(KEYINPUT37), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n475), .A2(new_n477), .A3(new_n478), .A4(new_n480), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n473), .A2(KEYINPUT87), .A3(new_n394), .A4(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT87), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n481), .A2(new_n394), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n483), .B1(new_n484), .B2(new_n442), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n475), .A2(new_n476), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n482), .A2(new_n485), .B1(KEYINPUT38), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n466), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n418), .B1(new_n429), .B2(new_n417), .ZN(new_n489));
  XOR2_X1   g288(.A(KEYINPUT85), .B(KEYINPUT39), .Z(new_n490));
  AOI21_X1  g289(.A(new_n407), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT39), .B1(new_n421), .B2(new_n422), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n491), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  XOR2_X1   g292(.A(new_n493), .B(KEYINPUT40), .Z(new_n494));
  INV_X1    g293(.A(new_n402), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n437), .A2(new_n407), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n488), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n467), .B(new_n472), .C1(new_n487), .C2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n465), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G113gat), .B(G141gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n501), .B(KEYINPUT92), .ZN(new_n502));
  XNOR2_X1  g301(.A(G169gat), .B(G197gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n502), .B(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n504), .B(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(KEYINPUT12), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(G29gat), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n509), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n510));
  XOR2_X1   g309(.A(KEYINPUT14), .B(G29gat), .Z(new_n511));
  OAI21_X1  g310(.A(new_n510), .B1(new_n511), .B2(G36gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(G43gat), .B(G50gat), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n513), .A2(KEYINPUT15), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT15), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT93), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n516), .B1(new_n513), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n518), .B1(new_n517), .B2(new_n513), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n512), .B(new_n518), .C1(new_n517), .C2(new_n513), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G15gat), .B(G22gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT95), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(G8gat), .ZN(new_n525));
  INV_X1    g324(.A(G8gat), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n523), .A2(KEYINPUT95), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT16), .ZN(new_n529));
  AOI21_X1  g328(.A(G1gat), .B1(new_n523), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n525), .A2(new_n530), .A3(new_n527), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n522), .B(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(G229gat), .A2(G233gat), .ZN(new_n536));
  XOR2_X1   g335(.A(new_n536), .B(KEYINPUT13), .Z(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n536), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n522), .A2(new_n534), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT17), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n520), .A2(new_n541), .A3(new_n521), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT94), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n520), .A2(KEYINPUT94), .A3(new_n521), .A4(new_n541), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n522), .A2(KEYINPUT17), .B1(new_n532), .B2(new_n533), .ZN(new_n547));
  AOI211_X1 g346(.A(new_n539), .B(new_n540), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n538), .B1(new_n548), .B2(KEYINPUT18), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n540), .B1(new_n546), .B2(new_n547), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(new_n536), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT18), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n508), .B1(new_n549), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n551), .A2(new_n552), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n548), .A2(KEYINPUT18), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n555), .A2(new_n556), .A3(new_n507), .A4(new_n538), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n554), .A2(KEYINPUT96), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT96), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n559), .B(new_n508), .C1(new_n549), .C2(new_n553), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(G71gat), .B(G78gat), .Z(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT9), .ZN(new_n565));
  INV_X1    g364(.A(G71gat), .ZN(new_n566));
  INV_X1    g365(.A(G78gat), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(G57gat), .B(G64gat), .Z(new_n569));
  NAND3_X1  g368(.A1(new_n564), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n568), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(new_n563), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT21), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G231gat), .A2(G233gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(G127gat), .ZN(new_n578));
  AND3_X1   g377(.A1(new_n572), .A2(KEYINPUT97), .A3(new_n570), .ZN(new_n579));
  AOI21_X1  g378(.A(KEYINPUT97), .B1(new_n570), .B2(new_n572), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n534), .B1(new_n581), .B2(new_n574), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n578), .B(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(G155gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(G183gat), .B(G211gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n583), .B(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(G232gat), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n589), .A2(new_n279), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT41), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G190gat), .B(G218gat), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT99), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n593), .B(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G134gat), .B(G162gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(G85gat), .A2(G92gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n600), .B(new_n601), .Z(new_n602));
  NAND2_X1  g401(.A1(G99gat), .A2(G106gat), .ZN(new_n603));
  INV_X1    g402(.A(G85gat), .ZN(new_n604));
  INV_X1    g403(.A(G92gat), .ZN(new_n605));
  AOI22_X1  g404(.A1(KEYINPUT8), .A2(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(G99gat), .B(G106gat), .Z(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n608), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n602), .A2(new_n610), .A3(new_n606), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  OAI22_X1  g411(.A1(new_n522), .A2(new_n612), .B1(new_n592), .B2(new_n591), .ZN(new_n613));
  AOI22_X1  g412(.A1(new_n522), .A2(KEYINPUT17), .B1(new_n611), .B2(new_n609), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n613), .B1(new_n546), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n594), .A2(new_n595), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n599), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NOR3_X1   g417(.A1(new_n615), .A2(new_n616), .A3(new_n599), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n598), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n619), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n621), .A2(new_n617), .A3(new_n597), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n588), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(G230gat), .A2(G233gat), .ZN(new_n625));
  XOR2_X1   g424(.A(KEYINPUT101), .B(KEYINPUT10), .Z(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  AND3_X1   g426(.A1(new_n602), .A2(new_n610), .A3(new_n606), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n610), .B1(new_n602), .B2(new_n606), .ZN(new_n629));
  OAI21_X1  g428(.A(KEYINPUT100), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT100), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n609), .A2(new_n631), .A3(new_n611), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n630), .A2(new_n632), .A3(new_n573), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n612), .A2(KEYINPUT100), .A3(new_n572), .A4(new_n570), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n627), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n609), .A2(KEYINPUT10), .A3(new_n611), .ZN(new_n636));
  NOR3_X1   g435(.A1(new_n636), .A2(new_n579), .A3(new_n580), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n625), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT102), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI211_X1 g439(.A(KEYINPUT102), .B(new_n625), .C1(new_n635), .C2(new_n637), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n633), .A2(new_n634), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(new_n625), .ZN(new_n643));
  XOR2_X1   g442(.A(G120gat), .B(G148gat), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT103), .ZN(new_n645));
  XNOR2_X1  g444(.A(G176gat), .B(G204gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n643), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n640), .A2(new_n641), .A3(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n638), .B1(new_n625), .B2(new_n642), .ZN(new_n651));
  AND3_X1   g450(.A1(new_n651), .A2(KEYINPUT104), .A3(new_n648), .ZN(new_n652));
  AOI21_X1  g451(.A(KEYINPUT104), .B1(new_n651), .B2(new_n648), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n650), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n500), .A2(new_n562), .A3(new_n624), .A4(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT105), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n660), .A2(new_n442), .ZN(new_n661));
  INV_X1    g460(.A(G1gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(G1324gat));
  XOR2_X1   g462(.A(KEYINPUT16), .B(G8gat), .Z(new_n664));
  OAI211_X1 g463(.A(new_n495), .B(new_n664), .C1(new_n658), .C2(new_n659), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT106), .ZN(new_n666));
  AND3_X1   g465(.A1(new_n665), .A2(new_n666), .A3(KEYINPUT42), .ZN(new_n667));
  AOI21_X1  g466(.A(KEYINPUT42), .B1(new_n665), .B2(new_n666), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n495), .B1(new_n658), .B2(new_n659), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n669), .A2(KEYINPUT107), .A3(G8gat), .ZN(new_n670));
  AOI21_X1  g469(.A(KEYINPUT107), .B1(new_n669), .B2(G8gat), .ZN(new_n671));
  OAI22_X1  g470(.A1(new_n667), .A2(new_n668), .B1(new_n670), .B2(new_n671), .ZN(G1325gat));
  OR3_X1    g471(.A1(new_n660), .A2(G15gat), .A3(new_n451), .ZN(new_n673));
  OAI21_X1  g472(.A(G15gat), .B1(new_n660), .B2(new_n472), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(G1326gat));
  NOR2_X1   g474(.A1(new_n660), .A2(new_n488), .ZN(new_n676));
  XOR2_X1   g475(.A(KEYINPUT43), .B(G22gat), .Z(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(G1327gat));
  NAND2_X1  g477(.A1(new_n500), .A2(new_n562), .ZN(new_n679));
  INV_X1    g478(.A(new_n623), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n588), .A2(new_n655), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n682), .A2(new_n509), .A3(new_n473), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT45), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n685), .B1(new_n500), .B2(new_n623), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT108), .B(KEYINPUT44), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  AOI211_X1 g487(.A(new_n680), .B(new_n688), .C1(new_n465), .C2(new_n499), .ZN(new_n689));
  OR2_X1    g488(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n681), .A2(new_n561), .ZN(new_n691));
  AND3_X1   g490(.A1(new_n690), .A2(new_n473), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n684), .B1(new_n509), .B2(new_n692), .ZN(G1328gat));
  INV_X1    g492(.A(G36gat), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n682), .A2(new_n694), .A3(new_n495), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT46), .Z(new_n696));
  NAND3_X1  g495(.A1(new_n690), .A2(new_n495), .A3(new_n691), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT109), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n690), .A2(KEYINPUT109), .A3(new_n495), .A4(new_n691), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n699), .A2(G36gat), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n696), .A2(new_n701), .ZN(G1329gat));
  INV_X1    g501(.A(new_n472), .ZN(new_n703));
  OAI211_X1 g502(.A(new_n703), .B(new_n691), .C1(new_n686), .C2(new_n689), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(G43gat), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n451), .A2(G43gat), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT47), .ZN(new_n707));
  AOI22_X1  g506(.A1(new_n682), .A2(new_n706), .B1(KEYINPUT110), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  OR2_X1    g508(.A1(new_n707), .A2(KEYINPUT110), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1330gat));
  NAND2_X1  g510(.A1(new_n682), .A2(new_n466), .ZN(new_n712));
  INV_X1    g511(.A(G50gat), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n488), .A2(new_n713), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n690), .A2(new_n691), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g517(.A1(new_n624), .A2(new_n561), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n719), .B1(new_n465), .B2(new_n499), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n654), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n721), .A2(new_n442), .ZN(new_n722));
  XOR2_X1   g521(.A(KEYINPUT111), .B(G57gat), .Z(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1332gat));
  NAND2_X1  g523(.A1(new_n654), .A2(new_n495), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n720), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n728));
  AND2_X1   g527(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n727), .B2(new_n728), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT112), .ZN(G1333gat));
  OAI21_X1  g531(.A(G71gat), .B1(new_n721), .B2(new_n472), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n655), .A2(new_n451), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n720), .A2(new_n566), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  XOR2_X1   g535(.A(new_n736), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n488), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(new_n567), .ZN(G1335gat));
  AOI21_X1  g538(.A(new_n680), .B1(new_n465), .B2(new_n499), .ZN(new_n740));
  INV_X1    g539(.A(new_n588), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n562), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT51), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n740), .A2(KEYINPUT51), .A3(new_n742), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n747), .A2(new_n604), .A3(new_n473), .A4(new_n654), .ZN(new_n748));
  INV_X1    g547(.A(new_n742), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n749), .A2(new_n655), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n750), .B1(new_n686), .B2(new_n689), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT113), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT113), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n753), .B(new_n750), .C1(new_n686), .C2(new_n689), .ZN(new_n754));
  AND3_X1   g553(.A1(new_n752), .A2(new_n473), .A3(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n748), .B1(new_n755), .B2(new_n604), .ZN(G1336gat));
  AOI211_X1 g555(.A(G92gat), .B(new_n725), .C1(new_n745), .C2(new_n746), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(G92gat), .B1(new_n751), .B2(new_n402), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n752), .A2(new_n495), .A3(new_n754), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n757), .B1(new_n762), .B2(G92gat), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n761), .B1(new_n763), .B2(new_n760), .ZN(G1337gat));
  INV_X1    g563(.A(G99gat), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n747), .A2(new_n765), .A3(new_n734), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n752), .A2(new_n703), .A3(new_n754), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n766), .B1(new_n767), .B2(new_n765), .ZN(G1338gat));
  NOR2_X1   g567(.A1(new_n488), .A2(G106gat), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  AOI211_X1 g569(.A(new_n655), .B(new_n770), .C1(new_n745), .C2(new_n746), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  XOR2_X1   g571(.A(KEYINPUT114), .B(G106gat), .Z(new_n773));
  OAI21_X1  g572(.A(new_n773), .B1(new_n751), .B2(new_n488), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT53), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n772), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n752), .A2(new_n466), .A3(new_n754), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n771), .B1(new_n777), .B2(new_n773), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n776), .B1(new_n778), .B2(new_n775), .ZN(G1339gat));
  INV_X1    g578(.A(KEYINPUT54), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n637), .B1(new_n642), .B2(new_n626), .ZN(new_n781));
  INV_X1    g580(.A(new_n625), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n640), .A2(new_n783), .A3(new_n641), .ZN(new_n784));
  INV_X1    g583(.A(new_n638), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n647), .B1(new_n785), .B2(new_n780), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n784), .A2(new_n786), .A3(KEYINPUT55), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n789), .A2(new_n650), .A3(new_n790), .ZN(new_n791));
  OAI22_X1  g590(.A1(new_n550), .A2(new_n536), .B1(new_n535), .B2(new_n537), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n506), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n620), .A2(new_n622), .A3(new_n557), .A4(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(KEYINPUT115), .B1(new_n791), .B2(new_n794), .ZN(new_n795));
  AND4_X1   g594(.A1(new_n557), .A2(new_n620), .A3(new_n622), .A4(new_n793), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n797));
  INV_X1    g596(.A(new_n650), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n798), .B1(new_n787), .B2(new_n788), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n796), .A2(new_n797), .A3(new_n790), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n795), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n799), .A2(new_n558), .A3(new_n560), .A4(new_n790), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n654), .A2(new_n557), .A3(new_n793), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n623), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n588), .B1(new_n801), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n624), .A2(new_n561), .A3(new_n655), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n442), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n807), .A2(new_n402), .A3(new_n454), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n562), .A2(new_n249), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(KEYINPUT116), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n466), .B1(new_n805), .B2(new_n806), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n495), .A2(new_n442), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n812), .A2(new_n295), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(G113gat), .B1(new_n814), .B2(new_n561), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n811), .A2(new_n815), .ZN(G1340gat));
  NAND2_X1  g615(.A1(new_n654), .A2(new_n252), .ZN(new_n817));
  XOR2_X1   g616(.A(new_n817), .B(KEYINPUT117), .Z(new_n818));
  NAND2_X1  g617(.A1(new_n808), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(G120gat), .B1(new_n814), .B2(new_n655), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(G1341gat));
  NAND3_X1  g620(.A1(new_n808), .A2(new_n260), .A3(new_n741), .ZN(new_n822));
  OAI21_X1  g621(.A(G127gat), .B1(new_n814), .B2(new_n588), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(G1342gat));
  NOR2_X1   g623(.A1(new_n680), .A2(new_n495), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n807), .A2(new_n258), .A3(new_n454), .A4(new_n825), .ZN(new_n826));
  OR2_X1    g625(.A1(new_n826), .A2(KEYINPUT56), .ZN(new_n827));
  OAI21_X1  g626(.A(G134gat), .B1(new_n814), .B2(new_n680), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(KEYINPUT56), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(G1343gat));
  NOR2_X1   g629(.A1(new_n703), .A2(new_n488), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n807), .A2(new_n831), .ZN(new_n832));
  NOR4_X1   g631(.A1(new_n832), .A2(G141gat), .A3(new_n495), .A4(new_n561), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT119), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT58), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n472), .A2(new_n813), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n805), .A2(new_n806), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT57), .B1(new_n838), .B2(new_n466), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT57), .ZN(new_n840));
  AOI211_X1 g639(.A(new_n840), .B(new_n488), .C1(new_n805), .C2(new_n806), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n562), .B(new_n837), .C1(new_n839), .C2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(G141gat), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n835), .B(new_n843), .C1(new_n834), .C2(new_n833), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n842), .A2(new_n845), .A3(G141gat), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n845), .B1(new_n842), .B2(G141gat), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n846), .A2(new_n847), .A3(new_n833), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT58), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n844), .B1(new_n848), .B2(new_n849), .ZN(G1344gat));
  NAND2_X1  g649(.A1(new_n320), .A2(new_n321), .ZN(new_n851));
  OR4_X1    g650(.A1(new_n851), .A2(new_n832), .A3(new_n495), .A4(new_n655), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n839), .A2(new_n841), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n837), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n854), .B1(new_n857), .B2(new_n654), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n791), .A2(new_n794), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n588), .B1(new_n804), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n806), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT57), .B1(new_n861), .B2(new_n466), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n654), .B(new_n837), .C1(new_n841), .C2(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n853), .B1(new_n863), .B2(G148gat), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n852), .B1(new_n858), .B2(new_n864), .ZN(G1345gat));
  OR2_X1    g664(.A1(new_n326), .A2(new_n327), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n741), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n855), .A2(new_n837), .A3(new_n867), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n807), .A2(new_n402), .A3(new_n741), .A4(new_n831), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT120), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n870), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI211_X1 g672(.A(KEYINPUT121), .B(new_n868), .C1(new_n873), .C2(new_n866), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT121), .ZN(new_n875));
  INV_X1    g674(.A(new_n868), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n866), .B1(new_n871), .B2(new_n872), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n874), .A2(new_n878), .ZN(G1346gat));
  INV_X1    g678(.A(KEYINPUT122), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n880), .B1(new_n856), .B2(new_n680), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(G162gat), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n856), .A2(new_n880), .A3(new_n680), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n825), .A2(new_n315), .ZN(new_n884));
  OAI22_X1  g683(.A1(new_n882), .A2(new_n883), .B1(new_n832), .B2(new_n884), .ZN(G1347gat));
  NOR2_X1   g684(.A1(new_n473), .A2(new_n402), .ZN(new_n886));
  AND3_X1   g685(.A1(new_n812), .A2(new_n295), .A3(new_n886), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n561), .A2(new_n206), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n473), .B1(new_n805), .B2(new_n806), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n454), .A2(new_n495), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n890), .B(KEYINPUT123), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n889), .A2(new_n562), .A3(new_n891), .ZN(new_n892));
  AOI22_X1  g691(.A1(new_n887), .A2(new_n888), .B1(new_n892), .B2(new_n206), .ZN(G1348gat));
  NAND3_X1  g692(.A1(new_n887), .A2(G176gat), .A3(new_n654), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT124), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n889), .A2(new_n891), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n207), .B1(new_n897), .B2(new_n655), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n894), .A2(new_n895), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n896), .A2(new_n898), .A3(new_n899), .ZN(G1349gat));
  INV_X1    g699(.A(new_n244), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n897), .A2(new_n901), .A3(new_n588), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n741), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(new_n903), .B2(G183gat), .ZN(new_n904));
  XOR2_X1   g703(.A(new_n904), .B(KEYINPUT60), .Z(G1350gat));
  NOR3_X1   g704(.A1(new_n897), .A2(G190gat), .A3(new_n680), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT125), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n887), .A2(new_n623), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n908), .B2(G190gat), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT61), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n906), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OR2_X1    g710(.A1(new_n909), .A2(new_n910), .ZN(new_n912));
  AOI211_X1 g711(.A(KEYINPUT125), .B(new_n220), .C1(new_n887), .C2(new_n623), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(G1351gat));
  AND2_X1   g713(.A1(new_n472), .A2(new_n886), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n915), .B1(new_n841), .B2(new_n862), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n916), .A2(new_n297), .A3(new_n561), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n889), .A2(new_n831), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n495), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(new_n562), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n917), .B1(new_n297), .B2(new_n921), .ZN(G1352gat));
  OAI21_X1  g721(.A(G204gat), .B1(new_n916), .B2(new_n655), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n725), .A2(G204gat), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n838), .A2(new_n442), .A3(new_n831), .A4(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT126), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT62), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT126), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n889), .A2(new_n928), .A3(new_n831), .A4(new_n924), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n926), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n927), .B1(new_n926), .B2(new_n929), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n923), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT127), .ZN(G1353gat));
  OR3_X1    g732(.A1(new_n919), .A2(G211gat), .A3(new_n588), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n916), .A2(new_n588), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n935), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n936));
  AOI21_X1  g735(.A(KEYINPUT63), .B1(new_n935), .B2(G211gat), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(G1354gat));
  OAI21_X1  g737(.A(G218gat), .B1(new_n916), .B2(new_n680), .ZN(new_n939));
  OR2_X1    g738(.A1(new_n680), .A2(G218gat), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n919), .B2(new_n940), .ZN(G1355gat));
endmodule


