//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 1 0 1 1 1 1 0 1 0 1 0 0 1 0 1 1 0 1 0 0 0 1 0 0 1 1 0 0 1 1 0 1 0 0 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n804, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n876, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929;
  INV_X1    g000(.A(KEYINPUT5), .ZN(new_n202));
  XOR2_X1   g001(.A(G113gat), .B(G120gat), .Z(new_n203));
  INV_X1    g002(.A(KEYINPUT1), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G127gat), .B(G134gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n203), .A2(new_n204), .A3(new_n206), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT77), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G148gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G141gat), .ZN(new_n214));
  INV_X1    g013(.A(G141gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G148gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n214), .A2(new_n216), .B1(KEYINPUT2), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT74), .ZN(new_n219));
  XNOR2_X1  g018(.A(G155gat), .B(G162gat), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(new_n219), .B2(new_n220), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT75), .B(G141gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n214), .B1(new_n223), .B2(new_n213), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT76), .B(G162gat), .ZN(new_n225));
  INV_X1    g024(.A(G155gat), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT2), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n224), .A2(new_n227), .A3(new_n220), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n222), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT80), .ZN(new_n231));
  OR2_X1    g030(.A1(new_n229), .A2(new_n210), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT80), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n212), .A2(new_n233), .A3(new_n229), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n231), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(G225gat), .A2(G233gat), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n202), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n229), .A2(new_n210), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT4), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  XOR2_X1   g040(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n241), .A2(KEYINPUT79), .B1(new_n232), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT79), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n239), .A2(new_n245), .A3(new_n240), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  AND2_X1   g046(.A1(new_n222), .A2(new_n228), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n229), .A2(KEYINPUT3), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n250), .A2(new_n251), .A3(new_n212), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n253), .A2(new_n237), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n247), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n232), .A2(new_n240), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n239), .A2(new_n243), .ZN(new_n258));
  AND2_X1   g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n254), .A2(new_n202), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G1gat), .B(G29gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(KEYINPUT0), .ZN(new_n263));
  XNOR2_X1  g062(.A(G57gat), .B(G85gat), .ZN(new_n264));
  XOR2_X1   g063(.A(new_n263), .B(new_n264), .Z(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT6), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n256), .A2(new_n265), .A3(new_n260), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n261), .A2(KEYINPUT6), .A3(new_n266), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(G113gat), .B(G141gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n274), .B(KEYINPUT88), .ZN(new_n275));
  XOR2_X1   g074(.A(G169gat), .B(G197gat), .Z(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(KEYINPUT12), .ZN(new_n280));
  XNOR2_X1  g079(.A(G15gat), .B(G22gat), .ZN(new_n281));
  INV_X1    g080(.A(G1gat), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n281), .A2(KEYINPUT16), .A3(new_n282), .ZN(new_n283));
  OR2_X1    g082(.A1(KEYINPUT90), .A2(G8gat), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n283), .B(new_n284), .C1(new_n282), .C2(new_n281), .ZN(new_n285));
  NAND2_X1  g084(.A1(KEYINPUT90), .A2(G8gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  XOR2_X1   g087(.A(G43gat), .B(G50gat), .Z(new_n289));
  INV_X1    g088(.A(KEYINPUT15), .ZN(new_n290));
  OR2_X1    g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n292));
  OR3_X1    g091(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n293));
  AOI22_X1  g092(.A1(new_n289), .A2(new_n290), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(G29gat), .A2(G36gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n291), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT89), .ZN(new_n297));
  OR2_X1    g096(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n292), .A2(new_n297), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(new_n293), .A3(new_n299), .ZN(new_n300));
  AND2_X1   g099(.A1(new_n300), .A2(new_n295), .ZN(new_n301));
  OAI211_X1 g100(.A(KEYINPUT17), .B(new_n296), .C1(new_n301), .C2(new_n291), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n296), .B1(new_n301), .B2(new_n291), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT17), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n288), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(G229gat), .A2(G233gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n287), .A2(new_n303), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT18), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n287), .B(new_n303), .ZN(new_n311));
  XOR2_X1   g110(.A(new_n307), .B(KEYINPUT13), .Z(new_n312));
  AOI22_X1  g111(.A1(new_n309), .A2(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  AND2_X1   g112(.A1(new_n306), .A2(new_n308), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n314), .A2(KEYINPUT18), .A3(new_n307), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n280), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n313), .A2(new_n315), .A3(new_n280), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G211gat), .B(G218gat), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT69), .ZN(new_n322));
  OR2_X1    g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AND2_X1   g122(.A1(G211gat), .A2(G218gat), .ZN(new_n324));
  AND2_X1   g123(.A1(G197gat), .A2(G204gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(G197gat), .A2(G204gat), .ZN(new_n326));
  OAI22_X1  g125(.A1(KEYINPUT22), .A2(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n323), .B(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT70), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n330));
  INV_X1    g129(.A(G183gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT27), .ZN(new_n332));
  AOI21_X1  g131(.A(G190gat), .B1(new_n332), .B2(KEYINPUT64), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n333), .B1(KEYINPUT64), .B2(new_n332), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT27), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G183gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n336), .B(KEYINPUT65), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n330), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(G190gat), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n336), .A2(new_n332), .A3(KEYINPUT28), .A4(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(G169gat), .ZN(new_n342));
  INV_X1    g141(.A(G176gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(G169gat), .A2(G176gat), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n344), .B1(new_n346), .B2(KEYINPUT26), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT67), .ZN(new_n348));
  OR2_X1    g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n344), .A2(KEYINPUT26), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n350), .B1(new_n347), .B2(new_n348), .ZN(new_n351));
  AOI22_X1  g150(.A1(new_n349), .A2(new_n351), .B1(G183gat), .B2(G190gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n341), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(G169gat), .A2(G176gat), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT23), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n354), .B(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(G183gat), .A2(G190gat), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n357), .A2(KEYINPUT24), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n358), .A2(new_n346), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n331), .A2(new_n339), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(KEYINPUT24), .A3(new_n357), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n356), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT25), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n362), .B(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n353), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT29), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(G226gat), .ZN(new_n368));
  INV_X1    g167(.A(G233gat), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n368), .A2(new_n369), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n365), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n329), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT70), .B1(new_n365), .B2(new_n371), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n328), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  XOR2_X1   g174(.A(G8gat), .B(G36gat), .Z(new_n376));
  XNOR2_X1  g175(.A(new_n376), .B(KEYINPUT72), .ZN(new_n377));
  XNOR2_X1  g176(.A(G64gat), .B(G92gat), .ZN(new_n378));
  XOR2_X1   g177(.A(new_n377), .B(new_n378), .Z(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n328), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n372), .A2(KEYINPUT71), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n372), .A2(KEYINPUT71), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n381), .B(new_n370), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n375), .A2(new_n380), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT30), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n380), .B1(new_n375), .B2(new_n384), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n385), .A2(KEYINPUT73), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT73), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n375), .A2(new_n391), .A3(new_n380), .A4(new_n384), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n390), .A2(new_n386), .A3(new_n392), .ZN(new_n393));
  AND2_X1   g192(.A1(new_n389), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT83), .ZN(new_n395));
  INV_X1    g194(.A(G22gat), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n381), .B1(new_n250), .B2(new_n366), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT81), .ZN(new_n398));
  AND2_X1   g197(.A1(new_n327), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n327), .A2(new_n398), .ZN(new_n400));
  OR3_X1    g199(.A1(new_n399), .A2(new_n400), .A3(new_n321), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n327), .A2(new_n398), .A3(new_n321), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(new_n366), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n248), .B1(new_n403), .B2(new_n249), .ZN(new_n404));
  INV_X1    g203(.A(G228gat), .ZN(new_n405));
  OAI22_X1  g204(.A1(new_n397), .A2(new_n404), .B1(new_n405), .B2(new_n369), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n249), .B1(new_n328), .B2(KEYINPUT29), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n229), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n408), .A2(G228gat), .A3(G233gat), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT82), .ZN(new_n410));
  NOR3_X1   g209(.A1(new_n409), .A2(new_n397), .A3(new_n410), .ZN(new_n411));
  AOI211_X1 g210(.A(new_n405), .B(new_n369), .C1(new_n407), .C2(new_n229), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n229), .A2(KEYINPUT3), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n328), .B1(new_n413), .B2(KEYINPUT29), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT82), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n396), .B(new_n406), .C1(new_n411), .C2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n410), .B1(new_n409), .B2(new_n397), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n412), .A2(KEYINPUT82), .A3(new_n414), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n396), .B1(new_n420), .B2(new_n406), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n395), .B1(new_n417), .B2(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(G78gat), .B(G106gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n423), .B(KEYINPUT31), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n424), .B(G50gat), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n406), .B1(new_n411), .B2(new_n415), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(G22gat), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n428), .A2(KEYINPUT83), .A3(new_n416), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n422), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n395), .B(new_n425), .C1(new_n417), .C2(new_n421), .ZN(new_n431));
  AND2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n365), .B(new_n210), .ZN(new_n433));
  NAND2_X1  g232(.A1(G227gat), .A2(G233gat), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT34), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT68), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n436), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  OR3_X1    g237(.A1(new_n433), .A2(new_n435), .A3(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n438), .B1(new_n433), .B2(new_n435), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT33), .B1(new_n433), .B2(new_n435), .ZN(new_n442));
  XNOR2_X1  g241(.A(G15gat), .B(G43gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(G71gat), .B(G99gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n443), .B(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n441), .A2(new_n446), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n439), .B(new_n440), .C1(new_n442), .C2(new_n445), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n435), .ZN(new_n449));
  AND2_X1   g248(.A1(new_n449), .A2(KEYINPUT32), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n447), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n450), .B1(new_n447), .B2(new_n448), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n394), .A2(new_n432), .A3(new_n272), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT35), .ZN(new_n456));
  INV_X1    g255(.A(new_n453), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n451), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n430), .A2(new_n431), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT35), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n460), .A2(new_n461), .A3(new_n272), .A4(new_n394), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n456), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n272), .A2(new_n393), .A3(new_n389), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n457), .A2(KEYINPUT36), .A3(new_n451), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT36), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n466), .B1(new_n452), .B2(new_n453), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n464), .A2(new_n459), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  AND2_X1   g267(.A1(new_n390), .A2(new_n392), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT37), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n375), .A2(new_n470), .A3(new_n384), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n381), .B1(new_n373), .B2(new_n374), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n328), .B(new_n370), .C1(new_n382), .C2(new_n383), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(KEYINPUT37), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT38), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n471), .A2(new_n474), .A3(new_n475), .A4(new_n379), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n469), .A2(new_n270), .A3(new_n271), .A4(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n375), .A2(new_n384), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT37), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n479), .A2(new_n379), .A3(new_n471), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT86), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(new_n481), .A3(KEYINPUT38), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n481), .B1(new_n480), .B2(KEYINPUT38), .ZN(new_n484));
  NOR3_X1   g283(.A1(new_n477), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n236), .B1(new_n259), .B2(new_n252), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT39), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n266), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n257), .A2(new_n258), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n237), .B1(new_n489), .B2(new_n253), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n490), .B(KEYINPUT39), .C1(new_n237), .C2(new_n235), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n488), .A2(KEYINPUT40), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT85), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT85), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n488), .A2(new_n494), .A3(new_n491), .A4(KEYINPUT40), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n488), .A2(new_n491), .ZN(new_n497));
  XNOR2_X1  g296(.A(KEYINPUT84), .B(KEYINPUT40), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n497), .A2(new_n498), .B1(new_n261), .B2(new_n266), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n432), .B1(new_n394), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n468), .B1(new_n485), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n320), .B1(new_n463), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT101), .ZN(new_n504));
  NAND2_X1  g303(.A1(G99gat), .A2(G106gat), .ZN(new_n505));
  OR2_X1    g304(.A1(G99gat), .A2(G106gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(G85gat), .A2(G92gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT7), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT7), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n509), .A2(G85gat), .A3(G92gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(G85gat), .ZN(new_n512));
  INV_X1    g311(.A(G92gat), .ZN(new_n513));
  AOI22_X1  g312(.A1(KEYINPUT8), .A2(new_n505), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI221_X4 g313(.A(KEYINPUT95), .B1(new_n505), .B2(new_n506), .C1(new_n511), .C2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT95), .ZN(new_n516));
  INV_X1    g315(.A(new_n505), .ZN(new_n517));
  NOR2_X1   g316(.A1(G99gat), .A2(G106gat), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n506), .A2(KEYINPUT95), .A3(new_n505), .ZN(new_n520));
  AND4_X1   g319(.A1(new_n519), .A2(new_n520), .A3(new_n511), .A4(new_n514), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n515), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n305), .A2(new_n302), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n520), .A2(new_n511), .A3(new_n514), .ZN(new_n524));
  INV_X1    g323(.A(new_n519), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n519), .A2(new_n520), .A3(new_n511), .A4(new_n514), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AND2_X1   g327(.A1(G232gat), .A2(G233gat), .ZN(new_n529));
  AOI22_X1  g328(.A1(new_n303), .A2(new_n528), .B1(KEYINPUT41), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n523), .A2(new_n530), .ZN(new_n531));
  XOR2_X1   g330(.A(G190gat), .B(G218gat), .Z(new_n532));
  AND2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n531), .A2(new_n532), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(G134gat), .B(G162gat), .Z(new_n536));
  NOR2_X1   g335(.A1(new_n529), .A2(KEYINPUT41), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n538), .A2(KEYINPUT96), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n538), .B(KEYINPUT96), .Z(new_n541));
  OAI21_X1  g340(.A(new_n541), .B1(new_n533), .B2(new_n534), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT21), .ZN(new_n544));
  INV_X1    g343(.A(G57gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(G64gat), .ZN(new_n546));
  INV_X1    g345(.A(G64gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(G57gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G71gat), .B(G78gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(G71gat), .A2(G78gat), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT9), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n549), .A2(new_n550), .A3(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(G71gat), .ZN(new_n555));
  INV_X1    g354(.A(G78gat), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n555), .A2(new_n556), .A3(KEYINPUT92), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n551), .A2(KEYINPUT91), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT92), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n559), .B1(G71gat), .B2(G78gat), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT91), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n561), .A2(G71gat), .A3(G78gat), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n557), .A2(new_n558), .A3(new_n560), .A4(new_n562), .ZN(new_n563));
  AOI22_X1  g362(.A1(new_n546), .A2(new_n548), .B1(new_n552), .B2(new_n551), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n554), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n288), .B1(new_n544), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n544), .ZN(new_n567));
  XNOR2_X1  g366(.A(G127gat), .B(G155gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n566), .B(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(G231gat), .A2(G233gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT93), .ZN(new_n572));
  XOR2_X1   g371(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(G183gat), .B(G211gat), .Z(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(KEYINPUT94), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n574), .B(new_n576), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n570), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n570), .A2(new_n577), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n543), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n565), .B1(new_n515), .B2(new_n521), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n549), .A2(new_n553), .ZN(new_n583));
  AND2_X1   g382(.A1(new_n558), .A2(new_n562), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n583), .A2(new_n584), .A3(new_n560), .A4(new_n557), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n526), .A2(new_n585), .A3(new_n554), .A4(new_n527), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT98), .ZN(new_n588));
  NAND2_X1  g387(.A1(G230gat), .A2(G233gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n587), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n582), .A2(new_n586), .A3(new_n590), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT98), .ZN(new_n593));
  XNOR2_X1  g392(.A(G120gat), .B(G148gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(G176gat), .B(G204gat), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n594), .B(new_n595), .Z(new_n596));
  NAND3_X1  g395(.A1(new_n591), .A2(new_n593), .A3(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT99), .ZN(new_n599));
  OAI211_X1 g398(.A(new_n554), .B(KEYINPUT10), .C1(new_n563), .C2(new_n564), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT97), .ZN(new_n602));
  AND3_X1   g401(.A1(new_n601), .A2(new_n528), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n602), .B1(new_n601), .B2(new_n528), .ZN(new_n604));
  OAI22_X1  g403(.A1(new_n587), .A2(KEYINPUT10), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n589), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n598), .A2(new_n599), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(KEYINPUT97), .B1(new_n522), .B2(new_n600), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n601), .A2(new_n528), .A3(new_n602), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n582), .A2(new_n586), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT10), .ZN(new_n611));
  AOI22_X1  g410(.A1(new_n608), .A2(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n612), .A2(new_n590), .ZN(new_n613));
  OAI21_X1  g412(.A(KEYINPUT99), .B1(new_n613), .B2(new_n597), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n607), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(KEYINPUT100), .B1(new_n612), .B2(new_n590), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT100), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n603), .A2(new_n604), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT10), .B1(new_n582), .B2(new_n586), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n618), .B(new_n589), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n596), .B1(new_n622), .B2(new_n592), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n616), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n581), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n503), .A2(new_n504), .A3(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n504), .B1(new_n503), .B2(new_n626), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n273), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(G1gat), .ZN(G1324gat));
  INV_X1    g430(.A(KEYINPUT42), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n463), .A2(new_n502), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n633), .A2(new_n319), .A3(new_n626), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(KEYINPUT101), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n394), .B1(new_n635), .B2(new_n627), .ZN(new_n636));
  XOR2_X1   g435(.A(KEYINPUT16), .B(G8gat), .Z(new_n637));
  AOI21_X1  g436(.A(new_n632), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n389), .A2(new_n393), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n639), .B1(new_n628), .B2(new_n629), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(G8gat), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT102), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n632), .A2(KEYINPUT102), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n643), .B1(new_n637), .B2(new_n644), .ZN(new_n645));
  AOI22_X1  g444(.A1(new_n638), .A2(new_n641), .B1(new_n636), .B2(new_n645), .ZN(G1325gat));
  NOR2_X1   g445(.A1(new_n628), .A2(new_n629), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n467), .A2(new_n465), .ZN(new_n648));
  OAI21_X1  g447(.A(G15gat), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OR2_X1    g448(.A1(new_n458), .A2(G15gat), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n649), .B1(new_n647), .B2(new_n650), .ZN(G1326gat));
  OAI21_X1  g450(.A(new_n459), .B1(new_n628), .B2(new_n629), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT43), .B(G22gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(G1327gat));
  INV_X1    g453(.A(KEYINPUT44), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n496), .A2(new_n499), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n459), .B1(new_n656), .B2(new_n639), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n273), .A2(new_n482), .A3(new_n476), .A4(new_n469), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n657), .B1(new_n658), .B2(new_n484), .ZN(new_n659));
  AOI22_X1  g458(.A1(new_n659), .A2(new_n468), .B1(new_n456), .B2(new_n462), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n655), .B1(new_n660), .B2(new_n543), .ZN(new_n661));
  INV_X1    g460(.A(new_n543), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n633), .A2(KEYINPUT44), .A3(new_n662), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n580), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(new_n624), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n317), .A2(KEYINPUT104), .A3(new_n318), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT104), .ZN(new_n669));
  INV_X1    g468(.A(new_n318), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n669), .B1(new_n670), .B2(new_n316), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n667), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT105), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n664), .A2(new_n273), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(G29gat), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n667), .A2(new_n662), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT103), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n633), .A2(new_n319), .A3(new_n678), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n679), .A2(G29gat), .A3(new_n272), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n680), .A2(KEYINPUT45), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(KEYINPUT45), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n676), .A2(new_n681), .A3(new_n682), .ZN(G1328gat));
  NOR3_X1   g482(.A1(new_n679), .A2(G36gat), .A3(new_n394), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT46), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n661), .A2(new_n663), .A3(new_n639), .A4(new_n674), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT106), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(G36gat), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n685), .B1(new_n688), .B2(new_n690), .ZN(G1329gat));
  INV_X1    g490(.A(new_n648), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n661), .A2(new_n663), .A3(new_n692), .A4(new_n674), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(G43gat), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n458), .A2(G43gat), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n503), .A2(new_n678), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g496(.A(KEYINPUT47), .B1(new_n696), .B2(KEYINPUT107), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI211_X1 g498(.A(new_n694), .B(new_n696), .C1(KEYINPUT107), .C2(KEYINPUT47), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(G1330gat));
  NAND4_X1  g500(.A1(new_n661), .A2(new_n663), .A3(new_n459), .A4(new_n674), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(G50gat), .ZN(new_n703));
  OR3_X1    g502(.A1(new_n679), .A2(G50gat), .A3(new_n432), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT48), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n703), .A2(KEYINPUT48), .A3(new_n704), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(G1331gat));
  NOR4_X1   g508(.A1(new_n672), .A2(new_n665), .A3(new_n662), .A4(new_n624), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n633), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n711), .A2(new_n272), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(new_n545), .ZN(G1332gat));
  AOI211_X1 g512(.A(new_n394), .B(new_n711), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n714));
  NOR2_X1   g513(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1333gat));
  AND2_X1   g515(.A1(new_n633), .A2(new_n710), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n555), .B1(new_n717), .B2(new_n692), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n711), .A2(G71gat), .A3(new_n458), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  XOR2_X1   g519(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(G1334gat));
  NOR2_X1   g521(.A1(new_n711), .A2(new_n432), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(new_n556), .ZN(G1335gat));
  NOR3_X1   g523(.A1(new_n272), .A2(G85gat), .A3(new_n624), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n672), .A2(new_n580), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n633), .A2(new_n662), .A3(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT110), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n728), .A2(KEYINPUT51), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n543), .B1(new_n463), .B2(new_n502), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n731), .B1(new_n732), .B2(new_n726), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n725), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n672), .A2(new_n580), .A3(new_n624), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n661), .A2(new_n663), .A3(new_n273), .A4(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT109), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(G85gat), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n736), .A2(new_n737), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n734), .B1(new_n739), .B2(new_n740), .ZN(G1336gat));
  NOR3_X1   g540(.A1(new_n394), .A2(G92gat), .A3(new_n624), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(new_n730), .B2(new_n733), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n661), .A2(new_n663), .A3(new_n639), .A4(new_n735), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(G92gat), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT52), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n743), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n727), .B(new_n748), .ZN(new_n749));
  AOI22_X1  g548(.A1(new_n749), .A2(new_n742), .B1(G92gat), .B2(new_n744), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n747), .B1(new_n750), .B2(new_n746), .ZN(G1337gat));
  NAND3_X1  g550(.A1(new_n664), .A2(new_n692), .A3(new_n735), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(G99gat), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n458), .A2(G99gat), .A3(new_n624), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n730), .B2(new_n733), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(G1338gat));
  NOR3_X1   g555(.A1(new_n432), .A2(G106gat), .A3(new_n624), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n757), .B1(new_n730), .B2(new_n733), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n661), .A2(new_n663), .A3(new_n459), .A4(new_n735), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G106gat), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT53), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n758), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  AOI22_X1  g561(.A1(new_n749), .A2(new_n757), .B1(G106gat), .B2(new_n759), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n762), .B1(new_n763), .B2(new_n761), .ZN(G1339gat));
  INV_X1    g563(.A(KEYINPUT54), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n617), .A2(new_n765), .A3(new_n621), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n612), .A2(new_n590), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n606), .A2(new_n767), .A3(KEYINPUT54), .ZN(new_n768));
  INV_X1    g567(.A(new_n596), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n766), .A2(KEYINPUT55), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n770), .A2(new_n615), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n765), .B1(new_n605), .B2(new_n589), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n596), .B1(new_n773), .B2(new_n767), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n766), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n772), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AOI211_X1 g576(.A(KEYINPUT113), .B(KEYINPUT55), .C1(new_n774), .C2(new_n766), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n771), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(KEYINPUT114), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT114), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n771), .B(new_n781), .C1(new_n777), .C2(new_n778), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n780), .A2(new_n672), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n624), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n311), .A2(new_n312), .ZN(new_n785));
  XOR2_X1   g584(.A(new_n785), .B(KEYINPUT115), .Z(new_n786));
  NOR2_X1   g585(.A1(new_n314), .A2(new_n307), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n279), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n784), .A2(new_n788), .A3(new_n318), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n662), .B1(new_n783), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n318), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n791), .A2(new_n543), .ZN(new_n792));
  AND3_X1   g591(.A1(new_n792), .A2(new_n780), .A3(new_n782), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n665), .B1(new_n790), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n625), .A2(new_n672), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(KEYINPUT112), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  AND4_X1   g596(.A1(new_n273), .A2(new_n797), .A3(new_n394), .A4(new_n460), .ZN(new_n798));
  AOI21_X1  g597(.A(G113gat), .B1(new_n798), .B2(new_n672), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n319), .A2(G113gat), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n799), .B1(new_n798), .B2(new_n800), .ZN(G1340gat));
  NAND2_X1  g600(.A1(new_n798), .A2(new_n784), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g602(.A1(new_n798), .A2(new_n580), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n804), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g604(.A1(new_n798), .A2(new_n662), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n806), .A2(G134gat), .ZN(new_n807));
  XOR2_X1   g606(.A(KEYINPUT116), .B(KEYINPUT56), .Z(new_n808));
  OR2_X1    g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n806), .A2(G134gat), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n807), .A2(new_n808), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(G1343gat));
  NAND3_X1  g611(.A1(new_n648), .A2(new_n273), .A3(new_n394), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(KEYINPUT117), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n432), .B1(new_n794), .B2(new_n796), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n815), .A2(KEYINPUT57), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n459), .A2(KEYINPUT57), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n775), .A2(new_n776), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n319), .A2(new_n771), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n662), .B1(new_n789), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n665), .B1(new_n793), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n817), .B1(new_n821), .B2(new_n796), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n814), .B1(new_n816), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n823), .A2(new_n320), .ZN(new_n824));
  INV_X1    g623(.A(new_n223), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT58), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n692), .A2(new_n272), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n815), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n815), .A2(KEYINPUT118), .A3(new_n828), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n831), .A2(new_n394), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n319), .A2(new_n215), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n827), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n829), .A2(new_n639), .A3(new_n834), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n814), .B(new_n672), .C1(new_n816), .C2(new_n822), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n836), .B1(new_n837), .B2(new_n223), .ZN(new_n838));
  OAI22_X1  g637(.A1(new_n826), .A2(new_n835), .B1(new_n838), .B2(new_n827), .ZN(G1344gat));
  OAI21_X1  g638(.A(KEYINPUT59), .B1(new_n833), .B2(new_n624), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n213), .ZN(new_n841));
  OR3_X1    g640(.A1(new_n823), .A2(KEYINPUT59), .A3(new_n624), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n817), .B1(new_n794), .B2(new_n796), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n791), .A2(new_n779), .A3(new_n543), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n665), .B1(new_n820), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n845), .B1(new_n319), .B2(new_n625), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT57), .B1(new_n846), .B2(new_n459), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n814), .A2(new_n784), .ZN(new_n849));
  OAI211_X1 g648(.A(KEYINPUT59), .B(G148gat), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n841), .A2(new_n842), .A3(new_n850), .ZN(G1345gat));
  OAI21_X1  g650(.A(G155gat), .B1(new_n823), .B2(new_n665), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n580), .A2(new_n226), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n852), .B1(new_n833), .B2(new_n853), .ZN(G1346gat));
  OAI211_X1 g653(.A(new_n814), .B(new_n662), .C1(new_n816), .C2(new_n822), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n225), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n858), .B1(new_n855), .B2(new_n856), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n662), .A2(new_n225), .ZN(new_n860));
  OAI22_X1  g659(.A1(new_n857), .A2(new_n859), .B1(new_n833), .B2(new_n860), .ZN(G1347gat));
  INV_X1    g660(.A(KEYINPUT121), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n460), .A2(new_n272), .A3(new_n639), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(KEYINPUT120), .B1(new_n797), .B2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT120), .ZN(new_n866));
  AOI211_X1 g665(.A(new_n866), .B(new_n863), .C1(new_n794), .C2(new_n796), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n319), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(G169gat), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n797), .A2(new_n342), .A3(new_n672), .A4(new_n864), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n862), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(new_n871), .ZN(new_n873));
  AOI211_X1 g672(.A(KEYINPUT121), .B(new_n873), .C1(new_n869), .C2(G169gat), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n872), .A2(new_n874), .ZN(G1348gat));
  NAND4_X1  g674(.A1(new_n797), .A2(new_n343), .A3(new_n784), .A4(new_n864), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n865), .A2(new_n867), .A3(new_n624), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n876), .B1(new_n877), .B2(new_n343), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n878), .B(KEYINPUT122), .ZN(G1349gat));
  INV_X1    g678(.A(KEYINPUT124), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(KEYINPUT60), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n880), .A2(KEYINPUT60), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n331), .B1(new_n868), .B2(new_n580), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n580), .A2(new_n336), .A3(new_n332), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n797), .A2(new_n864), .A3(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT123), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n885), .B(new_n886), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n881), .B(new_n882), .C1(new_n883), .C2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n797), .A2(new_n864), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n866), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n797), .A2(KEYINPUT120), .A3(new_n864), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n890), .A2(new_n580), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(G183gat), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n885), .B(KEYINPUT123), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n893), .A2(new_n880), .A3(KEYINPUT60), .A4(new_n894), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n888), .A2(new_n895), .ZN(G1350gat));
  INV_X1    g695(.A(KEYINPUT61), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n868), .A2(new_n662), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n897), .B1(new_n898), .B2(G190gat), .ZN(new_n899));
  AOI211_X1 g698(.A(KEYINPUT61), .B(new_n339), .C1(new_n868), .C2(new_n662), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n662), .A2(new_n339), .ZN(new_n901));
  OAI22_X1  g700(.A1(new_n899), .A2(new_n900), .B1(new_n889), .B2(new_n901), .ZN(G1351gat));
  NAND2_X1  g701(.A1(new_n639), .A2(new_n272), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n692), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n815), .A2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(G197gat), .B1(new_n906), .B2(new_n672), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n848), .A2(new_n692), .A3(new_n903), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n319), .A2(G197gat), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(G1352gat));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n784), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(G204gat), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n905), .A2(G204gat), .A3(new_n624), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n914), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n912), .A2(new_n915), .A3(new_n916), .ZN(G1353gat));
  OR3_X1    g716(.A1(new_n905), .A2(G211gat), .A3(new_n665), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n580), .B(new_n904), .C1(new_n843), .C2(new_n847), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n919), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n920));
  AOI21_X1  g719(.A(KEYINPUT63), .B1(new_n919), .B2(G211gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(G1354gat));
  INV_X1    g721(.A(G218gat), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n923), .B1(new_n905), .B2(new_n543), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n925), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n662), .A2(G218gat), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT126), .ZN(new_n929));
  AOI22_X1  g728(.A1(new_n926), .A2(new_n927), .B1(new_n908), .B2(new_n929), .ZN(G1355gat));
endmodule


