//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 1 0 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 0 0 0 1 1 1 1 0 1 1 0 1 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004;
  INV_X1    g000(.A(KEYINPUT4), .ZN(new_n187));
  INV_X1    g001(.A(G107), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT76), .B1(new_n188), .B2(G104), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT76), .ZN(new_n190));
  INV_X1    g004(.A(G104), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G107), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n189), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT3), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n194), .B1(new_n191), .B2(G107), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n188), .A2(KEYINPUT3), .A3(G104), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n193), .A2(new_n197), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n187), .B1(new_n198), .B2(G101), .ZN(new_n199));
  AOI22_X1  g013(.A1(new_n189), .A2(new_n192), .B1(new_n195), .B2(new_n196), .ZN(new_n200));
  INV_X1    g014(.A(G101), .ZN(new_n201));
  AOI21_X1  g015(.A(KEYINPUT77), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  AND4_X1   g016(.A1(KEYINPUT77), .A2(new_n193), .A3(new_n197), .A4(new_n201), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n199), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G119), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G116), .ZN(new_n206));
  INV_X1    g020(.A(G116), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G119), .ZN(new_n208));
  AND2_X1   g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT2), .B(G113), .ZN(new_n210));
  XNOR2_X1  g024(.A(new_n209), .B(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  NOR3_X1   g026(.A1(new_n200), .A2(KEYINPUT4), .A3(new_n201), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n204), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n193), .A2(new_n197), .A3(new_n201), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT77), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n200), .A2(KEYINPUT77), .A3(new_n201), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n209), .ZN(new_n221));
  OR2_X1    g035(.A1(new_n221), .A2(new_n210), .ZN(new_n222));
  XOR2_X1   g036(.A(G104), .B(G107), .Z(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G101), .ZN(new_n224));
  OR2_X1    g038(.A1(new_n206), .A2(KEYINPUT5), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n225), .A2(G113), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n209), .A2(KEYINPUT5), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n220), .A2(new_n222), .A3(new_n224), .A4(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n215), .A2(new_n229), .ZN(new_n230));
  XOR2_X1   g044(.A(G110), .B(G122), .Z(new_n231));
  NOR2_X1   g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT89), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n222), .B(new_n224), .C1(new_n202), .C2(new_n203), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n227), .A2(KEYINPUT88), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT88), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n209), .A2(new_n236), .A3(KEYINPUT5), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n235), .A2(new_n226), .A3(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n233), .B1(new_n234), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n224), .B1(new_n202), .B2(new_n203), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n228), .A2(new_n222), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AOI22_X1  g056(.A1(new_n218), .A2(new_n219), .B1(G101), .B2(new_n223), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n235), .A2(new_n226), .A3(new_n237), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n243), .A2(KEYINPUT89), .A3(new_n222), .A4(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n239), .A2(new_n242), .A3(new_n245), .ZN(new_n246));
  XOR2_X1   g060(.A(new_n231), .B(KEYINPUT8), .Z(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT84), .ZN(new_n249));
  INV_X1    g063(.A(G146), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G143), .ZN(new_n251));
  AND2_X1   g065(.A1(KEYINPUT0), .A2(G128), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT64), .B(G143), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n251), .B(new_n252), .C1(new_n253), .C2(new_n250), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT65), .ZN(new_n255));
  INV_X1    g069(.A(G143), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(KEYINPUT64), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT64), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G143), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G146), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT65), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n261), .A2(new_n262), .A3(new_n251), .A4(new_n252), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n255), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n250), .A2(G143), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n265), .B1(new_n253), .B2(new_n250), .ZN(new_n266));
  NOR2_X1   g080(.A1(KEYINPUT0), .A2(G128), .ZN(new_n267));
  NOR3_X1   g081(.A1(new_n266), .A2(new_n252), .A3(new_n267), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n249), .B(G125), .C1(new_n264), .C2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n257), .A2(new_n259), .A3(new_n250), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n270), .B1(G143), .B2(new_n250), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n252), .A2(new_n267), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n255), .A2(new_n263), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G125), .ZN(new_n274));
  OAI21_X1  g088(.A(KEYINPUT84), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT66), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n276), .B(KEYINPUT1), .C1(new_n256), .C2(G146), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G128), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n276), .B1(new_n251), .B2(KEYINPUT1), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(KEYINPUT67), .B1(new_n280), .B2(new_n266), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n256), .A2(G146), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT1), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT66), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n284), .A2(G128), .A3(new_n277), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT67), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(new_n271), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n282), .B1(new_n260), .B2(G146), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(new_n283), .A3(G128), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n281), .A2(new_n287), .A3(new_n274), .A4(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n269), .A2(new_n275), .A3(new_n290), .ZN(new_n291));
  XOR2_X1   g105(.A(KEYINPUT86), .B(G224), .Z(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT7), .B1(new_n293), .B2(G953), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n294), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n269), .A2(new_n275), .A3(new_n290), .A4(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n248), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT90), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n232), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n248), .A2(new_n295), .A3(KEYINPUT90), .A4(new_n297), .ZN(new_n301));
  AOI21_X1  g115(.A(G902), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(G210), .B1(G237), .B2(G902), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT91), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n293), .A2(G953), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT85), .B(KEYINPUT87), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n306), .B(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n291), .B(new_n308), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n215), .A2(KEYINPUT82), .A3(new_n229), .ZN(new_n310));
  AOI21_X1  g124(.A(KEYINPUT82), .B1(new_n215), .B2(new_n229), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n231), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n312), .B(KEYINPUT6), .C1(new_n231), .C2(new_n230), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT83), .ZN(new_n314));
  INV_X1    g128(.A(new_n231), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT82), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n230), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n215), .A2(KEYINPUT82), .A3(new_n229), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n315), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT6), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n314), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n320), .B(new_n231), .C1(new_n310), .C2(new_n311), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n322), .A2(KEYINPUT83), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n309), .B(new_n313), .C1(new_n321), .C2(new_n323), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n302), .A2(new_n305), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n305), .B1(new_n302), .B2(new_n324), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G902), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT96), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n329), .B1(new_n256), .B2(G128), .ZN(new_n330));
  INV_X1    g144(.A(G128), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(KEYINPUT96), .A3(G143), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n333), .B1(new_n331), .B2(new_n253), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n334), .B(G134), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n207), .A2(G122), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT14), .ZN(new_n337));
  INV_X1    g151(.A(G122), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G116), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n336), .A2(KEYINPUT14), .ZN(new_n341));
  OAI21_X1  g155(.A(G107), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n336), .A2(new_n339), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT95), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT95), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n336), .A2(new_n339), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n188), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n335), .A2(KEYINPUT97), .A3(new_n342), .A4(new_n348), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n334), .A2(G134), .ZN(new_n350));
  INV_X1    g164(.A(G134), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n260), .A2(G128), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n351), .B1(new_n352), .B2(new_n333), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n342), .B(new_n348), .C1(new_n350), .C2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT97), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n349), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n347), .B(new_n188), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT13), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n333), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n353), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n359), .A2(new_n351), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n358), .B(new_n361), .C1(new_n334), .C2(new_n362), .ZN(new_n363));
  XOR2_X1   g177(.A(KEYINPUT9), .B(G234), .Z(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G217), .ZN(new_n366));
  NOR3_X1   g180(.A1(new_n365), .A2(new_n366), .A3(G953), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n357), .A2(new_n363), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n367), .B1(new_n357), .B2(new_n363), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n328), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G478), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n371), .A2(KEYINPUT15), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  OAI221_X1 g187(.A(new_n328), .B1(KEYINPUT15), .B2(new_n371), .C1(new_n368), .C2(new_n369), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT98), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n373), .A2(new_n374), .A3(KEYINPUT98), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(G234), .A2(G237), .ZN(new_n380));
  INV_X1    g194(.A(G953), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n380), .A2(G952), .A3(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(KEYINPUT69), .B(G953), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n384), .A2(G902), .A3(new_n380), .ZN(new_n385));
  XOR2_X1   g199(.A(KEYINPUT21), .B(G898), .Z(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n382), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(G214), .B1(G237), .B2(G902), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n274), .A2(G140), .ZN(new_n392));
  XNOR2_X1  g206(.A(G125), .B(G140), .ZN(new_n393));
  MUX2_X1   g207(.A(new_n392), .B(new_n393), .S(KEYINPUT16), .Z(new_n394));
  AND2_X1   g208(.A1(new_n394), .A2(new_n250), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n394), .A2(new_n250), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G237), .ZN(new_n398));
  AND2_X1   g212(.A1(KEYINPUT69), .A2(G953), .ZN(new_n399));
  NOR2_X1   g213(.A1(KEYINPUT69), .A2(G953), .ZN(new_n400));
  OAI211_X1 g214(.A(G214), .B(new_n398), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n253), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n383), .A2(new_n256), .A3(G214), .A4(new_n398), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n403), .A3(G131), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT93), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n402), .A2(new_n403), .ZN(new_n406));
  INV_X1    g220(.A(G131), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT17), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT93), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n402), .A2(new_n403), .A3(new_n410), .A4(G131), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n405), .A2(new_n408), .A3(new_n409), .A4(new_n411), .ZN(new_n412));
  AND2_X1   g226(.A1(new_n405), .A2(new_n411), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n397), .B(new_n412), .C1(new_n413), .C2(new_n409), .ZN(new_n414));
  XNOR2_X1  g228(.A(G113), .B(G122), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n415), .B(new_n191), .ZN(new_n416));
  NAND2_X1  g230(.A1(KEYINPUT18), .A2(G131), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n406), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n393), .B(G146), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n402), .A2(new_n403), .A3(KEYINPUT18), .A4(G131), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n418), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT92), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n419), .B1(new_n406), .B2(new_n417), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(KEYINPUT92), .A3(new_n421), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  AND3_X1   g241(.A1(new_n414), .A2(new_n416), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n416), .B1(new_n414), .B2(new_n427), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n328), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G475), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT20), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n393), .B(KEYINPUT19), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n396), .B1(new_n250), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n405), .A2(new_n411), .A3(new_n408), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n422), .A2(new_n423), .ZN(new_n437));
  AOI21_X1  g251(.A(KEYINPUT92), .B1(new_n425), .B2(new_n421), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n416), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n414), .A2(new_n416), .A3(new_n427), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(G475), .A2(G902), .ZN(new_n444));
  XOR2_X1   g258(.A(new_n444), .B(KEYINPUT94), .Z(new_n445));
  AOI21_X1  g259(.A(new_n432), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n445), .ZN(new_n447));
  AOI211_X1 g261(.A(KEYINPUT20), .B(new_n447), .C1(new_n441), .C2(new_n442), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n431), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n379), .A2(new_n391), .A3(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n327), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(G221), .B1(new_n365), .B2(G902), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT79), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n331), .B1(new_n270), .B2(KEYINPUT1), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n454), .B1(new_n455), .B2(new_n288), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n251), .B1(new_n253), .B2(new_n250), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n283), .B1(new_n253), .B2(new_n250), .ZN(new_n458));
  OAI211_X1 g272(.A(KEYINPUT79), .B(new_n457), .C1(new_n458), .C2(new_n331), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n456), .A2(new_n459), .A3(new_n289), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n243), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT10), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n281), .A2(new_n289), .A3(new_n287), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n464), .A2(new_n243), .A3(KEYINPUT10), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT78), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n213), .B1(new_n220), .B2(new_n199), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n466), .B1(new_n467), .B2(new_n273), .ZN(new_n468));
  AND4_X1   g282(.A1(new_n466), .A2(new_n204), .A3(new_n273), .A4(new_n214), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n463), .B(new_n465), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n351), .A2(G137), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT11), .ZN(new_n472));
  INV_X1    g286(.A(G137), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n473), .A2(G134), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT11), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n476), .B1(new_n351), .B2(G137), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n472), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n478), .B(G131), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n470), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n383), .A2(G227), .ZN(new_n481));
  XNOR2_X1  g295(.A(G110), .B(G140), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n481), .B(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n460), .A2(new_n243), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n464), .A2(new_n243), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n479), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT12), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n240), .A2(new_n289), .A3(new_n281), .A4(new_n287), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n461), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(KEYINPUT12), .A3(new_n479), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n490), .A2(KEYINPUT80), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT80), .ZN(new_n495));
  AOI21_X1  g309(.A(KEYINPUT12), .B1(new_n492), .B2(new_n479), .ZN(new_n496));
  INV_X1    g310(.A(new_n479), .ZN(new_n497));
  AOI211_X1 g311(.A(new_n489), .B(new_n497), .C1(new_n491), .C2(new_n461), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n495), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n485), .A2(new_n494), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n470), .A2(new_n479), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n464), .A2(new_n243), .A3(KEYINPUT10), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n204), .A2(new_n273), .A3(new_n214), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(KEYINPUT78), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n467), .A2(new_n466), .A3(new_n273), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n502), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(new_n497), .A3(new_n463), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n501), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(KEYINPUT81), .B1(new_n508), .B2(new_n484), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT81), .ZN(new_n510));
  AOI211_X1 g324(.A(new_n510), .B(new_n483), .C1(new_n501), .C2(new_n507), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n500), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(G469), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(new_n513), .A3(new_n328), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n513), .A2(new_n328), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n485), .A2(new_n501), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n496), .A2(new_n498), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n484), .B1(new_n480), .B2(new_n518), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G469), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n514), .A2(new_n516), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n452), .A2(new_n453), .A3(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(G472), .A2(G902), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n474), .A2(new_n471), .ZN(new_n525));
  MUX2_X1   g339(.A(new_n525), .B(new_n478), .S(new_n407), .Z(new_n526));
  NAND2_X1  g340(.A1(new_n464), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n273), .A2(new_n479), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT30), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n527), .A2(KEYINPUT30), .A3(new_n528), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n212), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT68), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n383), .A2(G210), .A3(new_n398), .ZN(new_n535));
  XNOR2_X1  g349(.A(KEYINPUT26), .B(G101), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n535), .B(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n537), .B(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n527), .A2(new_n211), .A3(new_n528), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT68), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n531), .A2(new_n541), .A3(new_n212), .A4(new_n532), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n534), .A2(new_n539), .A3(new_n540), .A4(new_n542), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n543), .A2(KEYINPUT31), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n527), .A2(new_n211), .A3(new_n528), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n211), .B1(new_n527), .B2(new_n528), .ZN(new_n546));
  OAI21_X1  g360(.A(KEYINPUT28), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT28), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n540), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n539), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n552), .B1(new_n543), .B2(KEYINPUT31), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n524), .B1(new_n544), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT32), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n534), .A2(new_n540), .A3(new_n542), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n551), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT71), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n547), .A2(new_n559), .A3(new_n539), .A4(new_n549), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT29), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(KEYINPUT71), .B1(new_n550), .B2(new_n551), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n558), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT72), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n565), .B1(new_n547), .B2(new_n549), .ZN(new_n566));
  INV_X1    g380(.A(new_n546), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n540), .ZN(new_n568));
  AOI21_X1  g382(.A(KEYINPUT72), .B1(new_n568), .B2(KEYINPUT28), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n551), .A2(new_n561), .ZN(new_n571));
  AOI21_X1  g385(.A(G902), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n564), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(G472), .ZN(new_n574));
  OAI211_X1 g388(.A(KEYINPUT32), .B(new_n524), .C1(new_n544), .C2(new_n553), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n556), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(KEYINPUT75), .A2(KEYINPUT25), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n383), .A2(G221), .A3(G234), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(KEYINPUT22), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n579), .B(G137), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(KEYINPUT74), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n396), .B1(new_n250), .B2(new_n393), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n205), .A2(G128), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT23), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n331), .A2(G119), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT73), .ZN(new_n586));
  XOR2_X1   g400(.A(new_n584), .B(new_n586), .Z(new_n587));
  NAND2_X1  g401(.A1(new_n583), .A2(new_n585), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  XOR2_X1   g403(.A(KEYINPUT24), .B(G110), .Z(new_n590));
  OAI22_X1  g404(.A1(new_n587), .A2(G110), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n582), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n587), .A2(G110), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n589), .A2(new_n590), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n593), .B(new_n594), .C1(new_n395), .C2(new_n396), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n581), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n580), .A2(new_n592), .A3(new_n595), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n577), .B1(new_n599), .B2(G902), .ZN(new_n600));
  INV_X1    g414(.A(new_n577), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n597), .A2(new_n328), .A3(new_n598), .A4(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n366), .B1(G234), .B2(new_n328), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n599), .A2(G902), .A3(new_n604), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n576), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n523), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(new_n201), .ZN(G3));
  NAND2_X1  g424(.A1(new_n522), .A2(new_n453), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  OR2_X1    g426(.A1(new_n544), .A2(new_n553), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n328), .B1(new_n544), .B2(new_n553), .ZN(new_n614));
  AOI22_X1  g428(.A1(new_n524), .A2(new_n613), .B1(new_n614), .B2(G472), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n612), .A2(new_n607), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n302), .A2(new_n324), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT99), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n617), .A2(new_n618), .A3(new_n303), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n304), .A2(KEYINPUT99), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n303), .A2(new_n618), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n302), .A2(new_n324), .A3(new_n620), .A4(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n391), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n370), .A2(new_n371), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n626), .B1(new_n368), .B2(new_n369), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n357), .A2(new_n363), .ZN(new_n628));
  INV_X1    g442(.A(new_n367), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n357), .A2(new_n363), .A3(new_n367), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n630), .A2(KEYINPUT33), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n627), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n328), .A2(G478), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n625), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n449), .A2(new_n635), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n623), .A2(new_n624), .A3(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n616), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT100), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT34), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(new_n191), .ZN(G6));
  NOR2_X1   g456(.A1(new_n446), .A2(new_n448), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT101), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n431), .ZN(new_n646));
  INV_X1    g460(.A(new_n379), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n619), .A2(new_n647), .A3(new_n391), .A4(new_n622), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n616), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT35), .B(G107), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G9));
  NAND2_X1  g465(.A1(new_n603), .A2(new_n604), .ZN(new_n652));
  OR3_X1    g466(.A1(new_n581), .A2(KEYINPUT36), .A3(new_n596), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n596), .B1(new_n581), .B2(KEYINPUT36), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n604), .A2(G902), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(KEYINPUT102), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT102), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n653), .A2(new_n654), .A3(new_n658), .A4(new_n655), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n652), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n615), .A2(new_n522), .A3(new_n660), .A4(new_n453), .ZN(new_n661));
  INV_X1    g475(.A(new_n452), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT37), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G110), .ZN(G12));
  NAND3_X1  g479(.A1(new_n522), .A2(new_n660), .A3(new_n453), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n556), .A2(new_n575), .A3(new_n574), .ZN(new_n667));
  INV_X1    g481(.A(G900), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n382), .B1(new_n385), .B2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n645), .A2(new_n647), .A3(new_n431), .A4(new_n670), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n666), .A2(new_n667), .A3(new_n671), .ZN(new_n672));
  AND3_X1   g486(.A1(new_n619), .A2(new_n389), .A3(new_n622), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G128), .ZN(G30));
  XNOR2_X1  g489(.A(new_n669), .B(KEYINPUT39), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n611), .A2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT40), .ZN(new_n678));
  AOI211_X1 g492(.A(new_n390), .B(new_n660), .C1(new_n677), .C2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n327), .B(KEYINPUT38), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n568), .A2(new_n551), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n543), .A2(G472), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(G472), .A2(G902), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n682), .A2(KEYINPUT103), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(KEYINPUT103), .B1(new_n682), .B2(new_n683), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n556), .A3(new_n575), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n680), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n379), .A2(new_n450), .ZN(new_n690));
  OAI21_X1  g504(.A(KEYINPUT40), .B1(new_n611), .B2(new_n676), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n679), .A2(new_n689), .A3(new_n690), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(new_n253), .ZN(G45));
  AND3_X1   g507(.A1(new_n449), .A2(new_n635), .A3(new_n670), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n619), .A2(new_n389), .A3(new_n694), .A4(new_n622), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT104), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n666), .A2(new_n667), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G146), .ZN(G48));
  AND4_X1   g514(.A1(new_n507), .A2(new_n499), .A3(new_n494), .A4(new_n483), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n497), .B1(new_n506), .B2(new_n463), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n484), .B1(new_n480), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n510), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n508), .A2(KEYINPUT81), .A3(new_n484), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n701), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g520(.A(G469), .B1(new_n706), .B2(G902), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(new_n453), .A3(new_n514), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n608), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n637), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT41), .B(G113), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G15));
  NOR2_X1   g526(.A1(new_n648), .A2(new_n646), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G116), .ZN(G18));
  AND3_X1   g529(.A1(new_n652), .A2(new_n657), .A3(new_n659), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n619), .A2(new_n389), .A3(new_n622), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n708), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n647), .A2(new_n388), .A3(new_n449), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n718), .A2(new_n576), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G119), .ZN(G21));
  NAND4_X1  g535(.A1(new_n690), .A2(new_n619), .A3(new_n389), .A4(new_n622), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n708), .A2(new_n388), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n570), .A2(new_n539), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n543), .A2(KEYINPUT31), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n543), .A2(KEYINPUT31), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n524), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT105), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n614), .A2(new_n731), .A3(G472), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n731), .B1(new_n614), .B2(G472), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n607), .B(new_n730), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n734), .A2(KEYINPUT106), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n734), .A2(KEYINPUT106), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n723), .B(new_n724), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(KEYINPUT107), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n338), .ZN(G24));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n740));
  INV_X1    g554(.A(new_n514), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n513), .B1(new_n512), .B2(new_n328), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n743), .A2(new_n673), .A3(new_n453), .A4(new_n660), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n449), .A2(new_n635), .A3(new_n670), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(KEYINPUT108), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT108), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n449), .A2(new_n635), .A3(new_n747), .A4(new_n670), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n730), .B(new_n749), .C1(new_n732), .C2(new_n733), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n740), .B1(new_n744), .B2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n524), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n752), .B1(new_n727), .B2(new_n728), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n614), .A2(G472), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT105), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n614), .A2(new_n731), .A3(G472), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n753), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n718), .A2(KEYINPUT109), .A3(new_n757), .A4(new_n749), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n751), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G125), .ZN(G27));
  AND2_X1   g574(.A1(new_n576), .A2(new_n607), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n325), .A2(new_n326), .A3(new_n390), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n522), .A2(new_n762), .A3(new_n453), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n761), .A2(new_n749), .A3(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT42), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n761), .A2(new_n763), .A3(KEYINPUT42), .A4(new_n749), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(KEYINPUT110), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(new_n407), .ZN(G33));
  INV_X1    g584(.A(new_n671), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n763), .A2(new_n576), .A3(new_n607), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(KEYINPUT111), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n761), .A2(new_n763), .A3(new_n774), .A4(new_n771), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G134), .ZN(G36));
  INV_X1    g591(.A(KEYINPUT43), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n450), .A2(new_n778), .A3(new_n635), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT112), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n449), .B(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n635), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n779), .B1(new_n782), .B2(KEYINPUT43), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n660), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n615), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(KEYINPUT44), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT44), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n788), .B1(new_n784), .B2(new_n615), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n787), .A2(new_n762), .A3(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n453), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n520), .A2(KEYINPUT45), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n517), .A2(new_n519), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT45), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n792), .A2(G469), .A3(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT46), .B1(new_n796), .B2(new_n516), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(new_n741), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n796), .A2(KEYINPUT46), .A3(new_n516), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n791), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n801), .A2(new_n676), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n790), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(KEYINPUT113), .B(G137), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n803), .B(new_n804), .ZN(G39));
  INV_X1    g619(.A(KEYINPUT114), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT47), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n801), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n808), .ZN(new_n810));
  NOR2_X1   g624(.A1(KEYINPUT114), .A2(KEYINPUT47), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n810), .B1(new_n800), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n576), .A2(new_n607), .ZN(new_n813));
  INV_X1    g627(.A(new_n762), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n814), .A2(new_n745), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n809), .A2(new_n812), .A3(new_n813), .A4(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G140), .ZN(G42));
  AOI22_X1  g631(.A1(new_n809), .A2(new_n812), .B1(new_n791), .B2(new_n743), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n735), .A2(new_n736), .ZN(new_n819));
  INV_X1    g633(.A(new_n382), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n821), .A2(new_n762), .A3(new_n783), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n818), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n708), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n821), .A2(new_n824), .A3(new_n783), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n825), .A2(KEYINPUT50), .A3(new_n390), .A4(new_n680), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT50), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n821), .A2(new_n390), .A3(new_n824), .A4(new_n783), .ZN(new_n828));
  INV_X1    g642(.A(new_n680), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n823), .B1(new_n826), .B2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT51), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n832), .B1(new_n823), .B2(KEYINPUT117), .ZN(new_n833));
  INV_X1    g647(.A(new_n757), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n688), .A2(new_n607), .ZN(new_n835));
  OR2_X1    g649(.A1(new_n449), .A2(new_n635), .ZN(new_n836));
  OAI22_X1  g650(.A1(new_n784), .A2(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n814), .A2(new_n708), .A3(new_n820), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n831), .A2(new_n833), .A3(new_n839), .ZN(new_n840));
  AND4_X1   g654(.A1(new_n673), .A2(new_n821), .A3(new_n824), .A4(new_n783), .ZN(new_n841));
  INV_X1    g655(.A(G952), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n838), .A2(new_n761), .A3(new_n783), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT48), .ZN(new_n844));
  AOI211_X1 g658(.A(new_n842), .B(G953), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n845), .B1(new_n844), .B2(new_n843), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n841), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n840), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n833), .B1(new_n831), .B2(new_n839), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n636), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n838), .A2(new_n607), .A3(new_n851), .A4(new_n688), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT52), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n672), .A2(new_n673), .B1(new_n697), .B2(new_n698), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n759), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n687), .A2(new_n716), .A3(new_n670), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT115), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n611), .A2(new_n722), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n673), .A2(new_n453), .A3(new_n522), .A4(new_n690), .ZN(new_n861));
  OAI21_X1  g675(.A(KEYINPUT115), .B1(new_n856), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n853), .B1(new_n855), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n863), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n865), .A2(KEYINPUT52), .A3(new_n759), .A4(new_n854), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  OAI22_X1  g681(.A1(new_n523), .A2(new_n608), .B1(new_n661), .B2(new_n662), .ZN(new_n868));
  INV_X1    g682(.A(new_n327), .ZN(new_n869));
  INV_X1    g683(.A(new_n375), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n636), .B1(new_n449), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n869), .A2(new_n391), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n615), .A2(new_n607), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n872), .A2(new_n873), .A3(new_n611), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n868), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n646), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n576), .A2(new_n876), .A3(new_n870), .A4(new_n670), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n814), .B1(new_n877), .B2(new_n750), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n878), .A2(new_n612), .A3(new_n660), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n768), .A2(new_n776), .A3(new_n875), .A4(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n737), .A2(new_n710), .A3(new_n714), .A4(new_n720), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n867), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(KEYINPUT53), .ZN(new_n884));
  XNOR2_X1  g698(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n884), .B(KEYINPUT54), .C1(new_n883), .C2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n883), .A2(new_n885), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT53), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n867), .A2(new_n882), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT54), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n850), .A2(new_n852), .A3(new_n886), .A4(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n842), .A2(new_n381), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n835), .A2(new_n791), .A3(new_n390), .ZN(new_n895));
  INV_X1    g709(.A(new_n743), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n896), .A2(KEYINPUT49), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n782), .B1(new_n896), .B2(KEYINPUT49), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n895), .A2(new_n680), .A3(new_n897), .A4(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n894), .A2(new_n899), .ZN(G75));
  OAI21_X1  g714(.A(new_n313), .B1(new_n321), .B2(new_n323), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(new_n309), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(KEYINPUT55), .Z(new_n903));
  AND3_X1   g717(.A1(new_n867), .A2(new_n882), .A3(new_n888), .ZN(new_n904));
  INV_X1    g718(.A(new_n885), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n905), .B1(new_n867), .B2(new_n882), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT118), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n907), .A2(new_n908), .A3(G902), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n887), .A2(G902), .A3(new_n889), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(KEYINPUT118), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  AOI211_X1 g726(.A(KEYINPUT56), .B(new_n903), .C1(new_n912), .C2(new_n304), .ZN(new_n913));
  INV_X1    g727(.A(G210), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n903), .B1(new_n915), .B2(KEYINPUT56), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n383), .A2(G952), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n913), .A2(new_n919), .ZN(G51));
  XNOR2_X1  g734(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(new_n515), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n887), .A2(KEYINPUT54), .A3(new_n889), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n922), .B1(new_n923), .B2(new_n890), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT120), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI211_X1 g740(.A(KEYINPUT120), .B(new_n922), .C1(new_n923), .C2(new_n890), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n926), .A2(new_n512), .A3(new_n927), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n796), .B(KEYINPUT121), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n912), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n917), .B1(new_n928), .B2(new_n930), .ZN(G54));
  AOI21_X1  g745(.A(new_n908), .B1(new_n907), .B2(G902), .ZN(new_n932));
  NOR4_X1   g746(.A1(new_n904), .A2(new_n906), .A3(KEYINPUT118), .A4(new_n328), .ZN(new_n933));
  OAI211_X1 g747(.A(KEYINPUT58), .B(G475), .C1(new_n932), .C2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n443), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n912), .A2(KEYINPUT58), .A3(G475), .A4(new_n443), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n936), .A2(new_n937), .A3(new_n918), .ZN(G60));
  NAND2_X1  g752(.A1(G478), .A2(G902), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT59), .Z(new_n940));
  AOI21_X1  g754(.A(new_n940), .B1(new_n891), .B2(new_n886), .ZN(new_n941));
  INV_X1    g755(.A(new_n633), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n918), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n923), .A2(new_n890), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n944), .A2(new_n633), .A3(new_n940), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n943), .A2(new_n945), .ZN(G63));
  AND2_X1   g760(.A1(new_n653), .A2(new_n654), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT122), .ZN(new_n948));
  NAND2_X1  g762(.A1(G217), .A2(G902), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT60), .Z(new_n950));
  AOI21_X1  g764(.A(new_n948), .B1(new_n907), .B2(new_n950), .ZN(new_n951));
  AND4_X1   g765(.A1(new_n948), .A2(new_n887), .A3(new_n889), .A4(new_n950), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n947), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n907), .A2(new_n948), .A3(new_n950), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n887), .A2(new_n889), .A3(new_n950), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(KEYINPUT122), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n599), .B(KEYINPUT123), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n954), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n953), .A2(new_n918), .A3(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT61), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n953), .A2(KEYINPUT61), .A3(new_n918), .A4(new_n958), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(G66));
  OAI21_X1  g777(.A(G953), .B1(new_n293), .B2(new_n387), .ZN(new_n964));
  INV_X1    g778(.A(new_n875), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n881), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n964), .B1(new_n966), .B2(new_n384), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n901), .B1(G898), .B2(new_n383), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(G69));
  NAND2_X1  g783(.A1(new_n531), .A2(new_n532), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(new_n433), .Z(new_n971));
  NAND2_X1  g785(.A1(new_n384), .A2(G900), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n608), .A2(new_n722), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n802), .B1(new_n790), .B2(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n855), .B1(new_n775), .B2(new_n773), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n974), .A2(new_n975), .A3(new_n768), .A4(new_n816), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n971), .B(new_n972), .C1(new_n976), .C2(new_n384), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n692), .A2(new_n759), .A3(new_n854), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT62), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n692), .A2(KEYINPUT62), .A3(new_n759), .A4(new_n854), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n982), .A2(new_n816), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n677), .A2(new_n761), .A3(new_n762), .A4(new_n871), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT124), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n985), .B1(new_n790), .B2(new_n802), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n384), .B1(new_n983), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n977), .B1(new_n987), .B2(new_n971), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n383), .B1(G227), .B2(G900), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT125), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n989), .B1(new_n977), .B2(new_n990), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n988), .B(new_n991), .Z(G72));
  XNOR2_X1  g806(.A(new_n557), .B(KEYINPUT126), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n982), .A2(new_n816), .A3(new_n966), .A4(new_n986), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n683), .B(KEYINPUT63), .ZN(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  AOI211_X1 g810(.A(new_n551), .B(new_n993), .C1(new_n994), .C2(new_n996), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(KEYINPUT127), .ZN(new_n998));
  NOR3_X1   g812(.A1(new_n976), .A2(new_n881), .A3(new_n965), .ZN(new_n999));
  OAI211_X1 g813(.A(new_n551), .B(new_n993), .C1(new_n999), .C2(new_n995), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n884), .B1(new_n883), .B2(new_n885), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n1001), .A2(new_n995), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n558), .A2(new_n543), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n917), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AND3_X1   g818(.A1(new_n998), .A2(new_n1000), .A3(new_n1004), .ZN(G57));
endmodule


