

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754;

  INV_X1 U373 ( .A(n573), .ZN(n600) );
  NOR2_X2 U374 ( .A1(n695), .A2(n715), .ZN(n697) );
  XNOR2_X2 U375 ( .A(n382), .B(n381), .ZN(n547) );
  NAND2_X2 U376 ( .A1(n690), .A2(n433), .ZN(n419) );
  OR2_X2 U377 ( .A1(n690), .A2(n417), .ZN(n416) );
  XNOR2_X2 U378 ( .A(n430), .B(n739), .ZN(n690) );
  NOR2_X1 U379 ( .A1(n550), .A2(n549), .ZN(n476) );
  NOR2_X2 U380 ( .A1(n600), .A2(n644), .ZN(n611) );
  XNOR2_X1 U381 ( .A(n371), .B(KEYINPUT0), .ZN(n598) );
  XNOR2_X1 U382 ( .A(n465), .B(n464), .ZN(n550) );
  XOR2_X1 U383 ( .A(KEYINPUT104), .B(KEYINPUT11), .Z(n454) );
  INV_X2 U384 ( .A(G953), .ZN(n354) );
  XNOR2_X1 U385 ( .A(n390), .B(KEYINPUT110), .ZN(n705) );
  NOR2_X1 U386 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U387 ( .A1(n598), .A2(n481), .ZN(n485) );
  XNOR2_X1 U388 ( .A(n685), .B(n684), .ZN(n686) );
  XNOR2_X1 U389 ( .A(n521), .B(n520), .ZN(n594) );
  XNOR2_X1 U390 ( .A(n370), .B(KEYINPUT76), .ZN(n421) );
  XNOR2_X1 U391 ( .A(n486), .B(n403), .ZN(n581) );
  XNOR2_X1 U392 ( .A(n454), .B(n453), .ZN(n455) );
  INV_X1 U393 ( .A(n354), .ZN(n355) );
  XNOR2_X1 U394 ( .A(n467), .B(n466), .ZN(n486) );
  NAND2_X1 U395 ( .A1(n442), .A2(G224), .ZN(n370) );
  XNOR2_X1 U396 ( .A(G146), .B(G125), .ZN(n448) );
  INV_X1 U397 ( .A(G953), .ZN(n442) );
  BUF_X1 U398 ( .A(n564), .Z(n352) );
  BUF_X1 U399 ( .A(n698), .Z(n353) );
  AND2_X2 U400 ( .A1(n367), .A2(n365), .ZN(n698) );
  INV_X1 U401 ( .A(G134), .ZN(n466) );
  NOR2_X1 U402 ( .A1(n355), .A2(G237), .ZN(n494) );
  XNOR2_X1 U403 ( .A(n472), .B(n471), .ZN(n510) );
  XNOR2_X1 U404 ( .A(n449), .B(KEYINPUT10), .ZN(n580) );
  XNOR2_X1 U405 ( .A(n448), .B(n384), .ZN(n449) );
  INV_X1 U406 ( .A(G140), .ZN(n384) );
  XNOR2_X1 U407 ( .A(n387), .B(n544), .ZN(n572) );
  NAND2_X1 U408 ( .A1(n628), .A2(n514), .ZN(n521) );
  NOR2_X1 U409 ( .A1(n415), .A2(n576), .ZN(n414) );
  XOR2_X1 U410 ( .A(G116), .B(KEYINPUT5), .Z(n496) );
  NAND2_X1 U411 ( .A1(n356), .A2(n375), .ZN(n374) );
  XNOR2_X1 U412 ( .A(n546), .B(n363), .ZN(n375) );
  XNOR2_X1 U413 ( .A(G119), .B(G113), .ZN(n428) );
  XNOR2_X1 U414 ( .A(KEYINPUT70), .B(KEYINPUT3), .ZN(n427) );
  XNOR2_X1 U415 ( .A(n487), .B(n404), .ZN(n403) );
  INV_X1 U416 ( .A(G137), .ZN(n404) );
  NOR2_X1 U417 ( .A1(n419), .A2(n437), .ZN(n412) );
  INV_X1 U418 ( .A(G122), .ZN(n450) );
  XNOR2_X1 U419 ( .A(n455), .B(n420), .ZN(n456) );
  XNOR2_X1 U420 ( .A(G143), .B(G104), .ZN(n458) );
  AND2_X1 U421 ( .A1(n405), .A2(n538), .ZN(n558) );
  INV_X1 U422 ( .A(KEYINPUT28), .ZN(n406) );
  XNOR2_X1 U423 ( .A(n377), .B(KEYINPUT41), .ZN(n675) );
  AND2_X1 U424 ( .A1(n388), .A2(n615), .ZN(n552) );
  AND2_X1 U425 ( .A1(n542), .A2(n389), .ZN(n388) );
  INV_X1 U426 ( .A(n543), .ZN(n389) );
  INV_X1 U427 ( .A(G478), .ZN(n381) );
  OR2_X1 U428 ( .A1(n707), .A2(G902), .ZN(n382) );
  XNOR2_X1 U429 ( .A(n513), .B(n385), .ZN(n628) );
  XNOR2_X1 U430 ( .A(n580), .B(n386), .ZN(n385) );
  XNOR2_X1 U431 ( .A(n507), .B(n357), .ZN(n386) );
  INV_X1 U432 ( .A(n637), .ZN(n367) );
  NOR2_X1 U433 ( .A1(n354), .A2(G952), .ZN(n715) );
  AND2_X1 U434 ( .A1(n735), .A2(n400), .ZN(n569) );
  INV_X1 U435 ( .A(KEYINPUT47), .ZN(n401) );
  AND2_X1 U436 ( .A1(n664), .A2(n641), .ZN(n481) );
  INV_X1 U437 ( .A(KEYINPUT44), .ZN(n398) );
  XNOR2_X1 U438 ( .A(KEYINPUT12), .B(KEYINPUT102), .ZN(n453) );
  XNOR2_X1 U439 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n422) );
  NAND2_X1 U440 ( .A1(n433), .A2(n623), .ZN(n418) );
  OR2_X1 U441 ( .A1(n433), .A2(n623), .ZN(n417) );
  XNOR2_X1 U442 ( .A(n498), .B(n368), .ZN(n502) );
  XNOR2_X1 U443 ( .A(n500), .B(n497), .ZN(n368) );
  AND2_X1 U444 ( .A1(n372), .A2(n361), .ZN(n630) );
  XNOR2_X1 U445 ( .A(n374), .B(n373), .ZN(n372) );
  INV_X1 U446 ( .A(KEYINPUT48), .ZN(n373) );
  XNOR2_X1 U447 ( .A(G110), .B(G104), .ZN(n737) );
  XNOR2_X1 U448 ( .A(G119), .B(G128), .ZN(n508) );
  XOR2_X1 U449 ( .A(G110), .B(G137), .Z(n509) );
  NOR2_X1 U450 ( .A1(n563), .A2(n728), .ZN(n574) );
  NAND2_X1 U451 ( .A1(n396), .A2(n411), .ZN(n395) );
  XNOR2_X1 U452 ( .A(n574), .B(n369), .ZN(n566) );
  INV_X1 U453 ( .A(KEYINPUT114), .ZN(n369) );
  NOR2_X1 U454 ( .A1(n539), .A2(n644), .ZN(n615) );
  XOR2_X1 U455 ( .A(KEYINPUT62), .B(n699), .Z(n700) );
  XNOR2_X1 U456 ( .A(n383), .B(n473), .ZN(n707) );
  XNOR2_X1 U457 ( .A(n474), .B(n358), .ZN(n383) );
  XNOR2_X1 U458 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U459 ( .A(n690), .B(n692), .ZN(n693) );
  XNOR2_X1 U460 ( .A(n376), .B(KEYINPUT42), .ZN(n753) );
  XNOR2_X1 U461 ( .A(n545), .B(KEYINPUT40), .ZN(n754) );
  AND2_X1 U462 ( .A1(n353), .A2(G217), .ZN(n627) );
  AND2_X1 U463 ( .A1(n570), .A2(n569), .ZN(n356) );
  INV_X1 U464 ( .A(KEYINPUT85), .ZN(n437) );
  XOR2_X1 U465 ( .A(KEYINPUT94), .B(KEYINPUT24), .Z(n357) );
  XOR2_X1 U466 ( .A(n470), .B(n469), .Z(n358) );
  AND2_X1 U467 ( .A1(n630), .A2(KEYINPUT2), .ZN(n359) );
  AND2_X1 U468 ( .A1(n717), .A2(n619), .ZN(n360) );
  AND2_X1 U469 ( .A1(n736), .A2(n683), .ZN(n361) );
  AND2_X1 U470 ( .A1(n416), .A2(n418), .ZN(n362) );
  XNOR2_X1 U471 ( .A(n504), .B(n503), .ZN(n540) );
  XOR2_X1 U472 ( .A(KEYINPUT82), .B(KEYINPUT46), .Z(n363) );
  AND2_X1 U473 ( .A1(n626), .A2(n625), .ZN(n364) );
  INV_X1 U474 ( .A(n742), .ZN(n634) );
  NAND2_X1 U475 ( .A1(n366), .A2(n364), .ZN(n365) );
  NAND2_X1 U476 ( .A1(n742), .A2(n620), .ZN(n366) );
  AND2_X2 U477 ( .A1(n742), .A2(n359), .ZN(n637) );
  XNOR2_X2 U478 ( .A(n409), .B(KEYINPUT45), .ZN(n742) );
  XNOR2_X1 U479 ( .A(n457), .B(n456), .ZN(n461) );
  NAND2_X1 U480 ( .A1(n378), .A2(n360), .ZN(n409) );
  NOR2_X2 U481 ( .A1(n556), .A2(n447), .ZN(n371) );
  NAND2_X1 U482 ( .A1(n675), .A2(n558), .ZN(n376) );
  NAND2_X1 U483 ( .A1(n529), .A2(n657), .ZN(n377) );
  NAND2_X1 U484 ( .A1(n362), .A2(n419), .ZN(n578) );
  XNOR2_X1 U485 ( .A(n379), .B(n398), .ZN(n378) );
  NAND2_X1 U486 ( .A1(n380), .A2(n392), .ZN(n379) );
  XNOR2_X1 U487 ( .A(n597), .B(n399), .ZN(n380) );
  NAND2_X1 U488 ( .A1(n552), .A2(n659), .ZN(n387) );
  NAND2_X1 U489 ( .A1(n391), .A2(n595), .ZN(n390) );
  XNOR2_X1 U490 ( .A(n607), .B(n593), .ZN(n391) );
  AND2_X2 U491 ( .A1(n592), .A2(n600), .ZN(n607) );
  INV_X1 U492 ( .A(n751), .ZN(n392) );
  XNOR2_X2 U493 ( .A(n485), .B(n484), .ZN(n592) );
  XNOR2_X2 U494 ( .A(n564), .B(KEYINPUT19), .ZN(n556) );
  NAND2_X2 U495 ( .A1(n393), .A2(n395), .ZN(n564) );
  AND2_X2 U496 ( .A1(n394), .A2(n397), .ZN(n393) );
  INV_X1 U497 ( .A(n412), .ZN(n394) );
  NOR2_X1 U498 ( .A1(n410), .A2(KEYINPUT85), .ZN(n396) );
  NAND2_X1 U499 ( .A1(n413), .A2(KEYINPUT85), .ZN(n397) );
  INV_X1 U500 ( .A(KEYINPUT84), .ZN(n399) );
  XNOR2_X2 U501 ( .A(G122), .B(G116), .ZN(n426) );
  XNOR2_X2 U502 ( .A(n426), .B(G107), .ZN(n468) );
  NAND2_X1 U503 ( .A1(n402), .A2(n401), .ZN(n400) );
  OR2_X1 U504 ( .A1(n723), .A2(n726), .ZN(n402) );
  XNOR2_X1 U505 ( .A(n407), .B(n406), .ZN(n405) );
  NAND2_X1 U506 ( .A1(n614), .A2(n562), .ZN(n407) );
  INV_X1 U507 ( .A(n540), .ZN(n614) );
  XNOR2_X2 U508 ( .A(n499), .B(n737), .ZN(n491) );
  XNOR2_X2 U509 ( .A(n583), .B(n408), .ZN(n499) );
  XNOR2_X2 U510 ( .A(KEYINPUT68), .B(G101), .ZN(n408) );
  XNOR2_X2 U511 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n583) );
  INV_X1 U512 ( .A(n419), .ZN(n410) );
  INV_X1 U513 ( .A(n413), .ZN(n411) );
  NAND2_X1 U514 ( .A1(n416), .A2(n414), .ZN(n413) );
  INV_X1 U515 ( .A(n418), .ZN(n415) );
  XNOR2_X1 U516 ( .A(KEYINPUT101), .B(KEYINPUT103), .ZN(n420) );
  XNOR2_X1 U517 ( .A(G131), .B(KEYINPUT69), .ZN(n487) );
  INV_X1 U518 ( .A(KEYINPUT80), .ZN(n631) );
  XNOR2_X1 U519 ( .A(n421), .B(n448), .ZN(n424) );
  XNOR2_X2 U520 ( .A(G143), .B(G128), .ZN(n467) );
  XNOR2_X1 U521 ( .A(n467), .B(n422), .ZN(n423) );
  XNOR2_X1 U522 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U523 ( .A(n425), .B(n491), .ZN(n430) );
  XNOR2_X1 U524 ( .A(n468), .B(KEYINPUT16), .ZN(n429) );
  XNOR2_X1 U525 ( .A(n428), .B(n427), .ZN(n497) );
  XNOR2_X1 U526 ( .A(n429), .B(n497), .ZN(n739) );
  XNOR2_X1 U527 ( .A(G902), .B(KEYINPUT15), .ZN(n477) );
  INV_X1 U528 ( .A(n477), .ZN(n623) );
  INV_X1 U529 ( .A(G902), .ZN(n514) );
  INV_X1 U530 ( .A(G237), .ZN(n431) );
  NAND2_X1 U531 ( .A1(n514), .A2(n431), .ZN(n434) );
  NAND2_X1 U532 ( .A1(n434), .A2(G210), .ZN(n432) );
  XNOR2_X1 U533 ( .A(n432), .B(KEYINPUT88), .ZN(n433) );
  NAND2_X1 U534 ( .A1(n434), .A2(G214), .ZN(n436) );
  INV_X1 U535 ( .A(KEYINPUT89), .ZN(n435) );
  XNOR2_X1 U536 ( .A(n436), .B(n435), .ZN(n657) );
  INV_X1 U537 ( .A(n657), .ZN(n576) );
  XOR2_X1 U538 ( .A(KEYINPUT73), .B(KEYINPUT14), .Z(n439) );
  NAND2_X1 U539 ( .A1(G234), .A2(G237), .ZN(n438) );
  XNOR2_X1 U540 ( .A(n439), .B(n438), .ZN(n445) );
  NAND2_X1 U541 ( .A1(n445), .A2(G952), .ZN(n441) );
  INV_X1 U542 ( .A(KEYINPUT90), .ZN(n440) );
  XNOR2_X1 U543 ( .A(n441), .B(n440), .ZN(n672) );
  NAND2_X1 U544 ( .A1(n672), .A2(n354), .ZN(n443) );
  XNOR2_X1 U545 ( .A(n443), .B(KEYINPUT91), .ZN(n534) );
  AND2_X1 U546 ( .A1(n355), .A2(G902), .ZN(n444) );
  NAND2_X1 U547 ( .A1(n445), .A2(n444), .ZN(n530) );
  NOR2_X1 U548 ( .A1(n530), .A2(G898), .ZN(n446) );
  NOR2_X1 U549 ( .A1(n534), .A2(n446), .ZN(n447) );
  XNOR2_X1 U550 ( .A(G113), .B(G131), .ZN(n451) );
  XNOR2_X1 U551 ( .A(n580), .B(n452), .ZN(n463) );
  NAND2_X1 U552 ( .A1(G214), .A2(n494), .ZN(n457) );
  XOR2_X1 U553 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n459) );
  XNOR2_X1 U554 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U555 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U556 ( .A(n463), .B(n462), .ZN(n685) );
  NOR2_X1 U557 ( .A1(G902), .A2(n685), .ZN(n465) );
  XNOR2_X1 U558 ( .A(KEYINPUT13), .B(G475), .ZN(n464) );
  XNOR2_X1 U559 ( .A(n486), .B(n468), .ZN(n474) );
  XOR2_X1 U560 ( .A(KEYINPUT105), .B(KEYINPUT7), .Z(n470) );
  XNOR2_X1 U561 ( .A(KEYINPUT106), .B(KEYINPUT9), .ZN(n469) );
  NAND2_X1 U562 ( .A1(n354), .A2(G234), .ZN(n472) );
  INV_X1 U563 ( .A(KEYINPUT8), .ZN(n471) );
  NAND2_X1 U564 ( .A1(n510), .A2(G217), .ZN(n473) );
  INV_X1 U565 ( .A(n547), .ZN(n549) );
  INV_X1 U566 ( .A(KEYINPUT107), .ZN(n475) );
  XNOR2_X2 U567 ( .A(n476), .B(n475), .ZN(n664) );
  NAND2_X1 U568 ( .A1(n477), .A2(G234), .ZN(n478) );
  XNOR2_X1 U569 ( .A(n478), .B(KEYINPUT20), .ZN(n515) );
  AND2_X1 U570 ( .A1(n515), .A2(G221), .ZN(n480) );
  XNOR2_X1 U571 ( .A(KEYINPUT98), .B(KEYINPUT21), .ZN(n479) );
  XNOR2_X1 U572 ( .A(n480), .B(n479), .ZN(n641) );
  XNOR2_X1 U573 ( .A(KEYINPUT72), .B(KEYINPUT22), .ZN(n483) );
  INV_X1 U574 ( .A(KEYINPUT66), .ZN(n482) );
  XNOR2_X1 U575 ( .A(n483), .B(n482), .ZN(n484) );
  INV_X1 U576 ( .A(n592), .ZN(n525) );
  XNOR2_X1 U577 ( .A(G146), .B(n581), .ZN(n501) );
  NAND2_X1 U578 ( .A1(n354), .A2(G227), .ZN(n489) );
  XOR2_X1 U579 ( .A(G107), .B(G140), .Z(n488) );
  XNOR2_X1 U580 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U581 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U582 ( .A(n501), .B(n492), .ZN(n712) );
  NAND2_X1 U583 ( .A1(n712), .A2(n514), .ZN(n493) );
  XNOR2_X1 U584 ( .A(n493), .B(G469), .ZN(n538) );
  XNOR2_X1 U585 ( .A(n538), .B(KEYINPUT1), .ZN(n573) );
  NAND2_X1 U586 ( .A1(n494), .A2(G210), .ZN(n495) );
  XNOR2_X1 U587 ( .A(n496), .B(n495), .ZN(n498) );
  INV_X1 U588 ( .A(n499), .ZN(n500) );
  XNOR2_X1 U589 ( .A(n502), .B(n501), .ZN(n699) );
  NAND2_X1 U590 ( .A1(n699), .A2(n514), .ZN(n504) );
  INV_X1 U591 ( .A(G472), .ZN(n503) );
  XNOR2_X1 U592 ( .A(n540), .B(KEYINPUT6), .ZN(n609) );
  XOR2_X1 U593 ( .A(KEYINPUT95), .B(KEYINPUT92), .Z(n506) );
  XNOR2_X1 U594 ( .A(KEYINPUT93), .B(KEYINPUT23), .ZN(n505) );
  XNOR2_X1 U595 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U596 ( .A(n509), .B(n508), .ZN(n512) );
  AND2_X1 U597 ( .A1(n510), .A2(G221), .ZN(n511) );
  XNOR2_X1 U598 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U599 ( .A(KEYINPUT75), .B(KEYINPUT25), .ZN(n517) );
  NAND2_X1 U600 ( .A1(G217), .A2(n515), .ZN(n516) );
  XNOR2_X1 U601 ( .A(n517), .B(n516), .ZN(n519) );
  XOR2_X1 U602 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n518) );
  XNOR2_X1 U603 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U604 ( .A(n594), .B(KEYINPUT108), .ZN(n640) );
  NOR2_X1 U605 ( .A1(n609), .A2(n640), .ZN(n522) );
  NAND2_X1 U606 ( .A1(n573), .A2(n522), .ZN(n523) );
  XOR2_X1 U607 ( .A(KEYINPUT77), .B(n523), .Z(n524) );
  NOR2_X1 U608 ( .A1(n525), .A2(n524), .ZN(n527) );
  XNOR2_X1 U609 ( .A(KEYINPUT65), .B(KEYINPUT32), .ZN(n526) );
  XNOR2_X1 U610 ( .A(n527), .B(n526), .ZN(n596) );
  XNOR2_X1 U611 ( .A(n596), .B(G119), .ZN(G21) );
  XNOR2_X1 U612 ( .A(KEYINPUT74), .B(KEYINPUT38), .ZN(n528) );
  XNOR2_X1 U613 ( .A(n578), .B(n528), .ZN(n659) );
  AND2_X1 U614 ( .A1(n659), .A2(n664), .ZN(n529) );
  INV_X1 U615 ( .A(n641), .ZN(n536) );
  XOR2_X1 U616 ( .A(KEYINPUT111), .B(n530), .Z(n531) );
  NOR2_X1 U617 ( .A1(G900), .A2(n531), .ZN(n532) );
  XNOR2_X1 U618 ( .A(n532), .B(KEYINPUT112), .ZN(n533) );
  NOR2_X1 U619 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U620 ( .A(KEYINPUT78), .B(n535), .ZN(n543) );
  OR2_X1 U621 ( .A1(n536), .A2(n543), .ZN(n537) );
  NOR2_X1 U622 ( .A1(n594), .A2(n537), .ZN(n562) );
  INV_X1 U623 ( .A(n538), .ZN(n539) );
  XOR2_X1 U624 ( .A(KEYINPUT83), .B(KEYINPUT39), .Z(n544) );
  NAND2_X1 U625 ( .A1(n641), .A2(n594), .ZN(n644) );
  NOR2_X1 U626 ( .A1(n576), .A2(n540), .ZN(n541) );
  XNOR2_X1 U627 ( .A(n541), .B(KEYINPUT30), .ZN(n542) );
  NAND2_X1 U628 ( .A1(n550), .A2(n547), .ZN(n728) );
  INV_X1 U629 ( .A(n728), .ZN(n548) );
  NAND2_X1 U630 ( .A1(n572), .A2(n548), .ZN(n545) );
  NAND2_X1 U631 ( .A1(n753), .A2(n754), .ZN(n546) );
  NOR2_X1 U632 ( .A1(n550), .A2(n547), .ZN(n571) );
  NOR2_X1 U633 ( .A1(n548), .A2(n571), .ZN(n617) );
  NAND2_X1 U634 ( .A1(n617), .A2(KEYINPUT47), .ZN(n554) );
  NAND2_X1 U635 ( .A1(n550), .A2(n549), .ZN(n604) );
  NOR2_X1 U636 ( .A1(n578), .A2(n604), .ZN(n551) );
  AND2_X1 U637 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U638 ( .A(n553), .B(KEYINPUT113), .ZN(n752) );
  NAND2_X1 U639 ( .A1(n554), .A2(n752), .ZN(n555) );
  XNOR2_X1 U640 ( .A(n555), .B(KEYINPUT79), .ZN(n560) );
  INV_X1 U641 ( .A(n556), .ZN(n557) );
  NAND2_X1 U642 ( .A1(n558), .A2(n557), .ZN(n561) );
  NAND2_X1 U643 ( .A1(n561), .A2(KEYINPUT47), .ZN(n559) );
  AND2_X1 U644 ( .A1(n560), .A2(n559), .ZN(n570) );
  INV_X1 U645 ( .A(n571), .ZN(n731) );
  NOR2_X1 U646 ( .A1(n561), .A2(n731), .ZN(n723) );
  NOR2_X1 U647 ( .A1(n561), .A2(n728), .ZN(n726) );
  NAND2_X1 U648 ( .A1(n562), .A2(n609), .ZN(n563) );
  INV_X1 U649 ( .A(n352), .ZN(n565) );
  NOR2_X1 U650 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U651 ( .A(n567), .B(KEYINPUT36), .ZN(n568) );
  NAND2_X1 U652 ( .A1(n568), .A2(n573), .ZN(n735) );
  NAND2_X1 U653 ( .A1(n572), .A2(n571), .ZN(n736) );
  NAND2_X1 U654 ( .A1(n600), .A2(n574), .ZN(n575) );
  NOR2_X1 U655 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U656 ( .A(n577), .B(KEYINPUT43), .Z(n579) );
  NAND2_X1 U657 ( .A1(n579), .A2(n578), .ZN(n683) );
  XNOR2_X1 U658 ( .A(n580), .B(KEYINPUT126), .ZN(n582) );
  XNOR2_X1 U659 ( .A(n582), .B(n581), .ZN(n584) );
  XNOR2_X1 U660 ( .A(n584), .B(n583), .ZN(n586) );
  XNOR2_X1 U661 ( .A(n630), .B(n586), .ZN(n585) );
  NAND2_X1 U662 ( .A1(n585), .A2(n354), .ZN(n591) );
  XNOR2_X1 U663 ( .A(n586), .B(G227), .ZN(n587) );
  XNOR2_X1 U664 ( .A(n587), .B(KEYINPUT127), .ZN(n588) );
  NAND2_X1 U665 ( .A1(n588), .A2(G900), .ZN(n589) );
  NAND2_X1 U666 ( .A1(n355), .A2(n589), .ZN(n590) );
  NAND2_X1 U667 ( .A1(n591), .A2(n590), .ZN(G72) );
  AND2_X1 U668 ( .A1(n630), .A2(n623), .ZN(n620) );
  INV_X1 U669 ( .A(KEYINPUT109), .ZN(n593) );
  NOR2_X1 U670 ( .A1(n614), .A2(n594), .ZN(n595) );
  NAND2_X1 U671 ( .A1(n705), .A2(n596), .ZN(n597) );
  BUF_X1 U672 ( .A(n598), .Z(n599) );
  XOR2_X1 U673 ( .A(KEYINPUT33), .B(KEYINPUT71), .Z(n602) );
  NAND2_X1 U674 ( .A1(n611), .A2(n609), .ZN(n601) );
  XNOR2_X2 U675 ( .A(n602), .B(n601), .ZN(n674) );
  NAND2_X1 U676 ( .A1(n599), .A2(n674), .ZN(n603) );
  XNOR2_X1 U677 ( .A(n603), .B(KEYINPUT34), .ZN(n605) );
  XOR2_X1 U678 ( .A(KEYINPUT35), .B(n606), .Z(n751) );
  INV_X1 U679 ( .A(n640), .ZN(n608) );
  NOR2_X1 U680 ( .A1(n609), .A2(n608), .ZN(n610) );
  NAND2_X1 U681 ( .A1(n607), .A2(n610), .ZN(n717) );
  INV_X1 U682 ( .A(n599), .ZN(n612) );
  NAND2_X1 U683 ( .A1(n614), .A2(n611), .ZN(n649) );
  NOR2_X1 U684 ( .A1(n612), .A2(n649), .ZN(n613) );
  XNOR2_X1 U685 ( .A(n613), .B(KEYINPUT31), .ZN(n730) );
  AND2_X1 U686 ( .A1(n615), .A2(n540), .ZN(n616) );
  NAND2_X1 U687 ( .A1(n616), .A2(n599), .ZN(n719) );
  NAND2_X1 U688 ( .A1(n730), .A2(n719), .ZN(n618) );
  INV_X1 U689 ( .A(n617), .ZN(n653) );
  NAND2_X1 U690 ( .A1(n618), .A2(n653), .ZN(n619) );
  INV_X1 U691 ( .A(KEYINPUT67), .ZN(n621) );
  NAND2_X1 U692 ( .A1(n621), .A2(KEYINPUT2), .ZN(n622) );
  OR2_X1 U693 ( .A1(n477), .A2(n622), .ZN(n626) );
  NAND2_X1 U694 ( .A1(n623), .A2(KEYINPUT2), .ZN(n624) );
  NAND2_X1 U695 ( .A1(n624), .A2(KEYINPUT67), .ZN(n625) );
  XNOR2_X1 U696 ( .A(n628), .B(n627), .ZN(n629) );
  NOR2_X1 U697 ( .A1(n629), .A2(n715), .ZN(G66) );
  NOR2_X1 U698 ( .A1(n630), .A2(KEYINPUT2), .ZN(n632) );
  XNOR2_X1 U699 ( .A(n632), .B(n631), .ZN(n636) );
  INV_X1 U700 ( .A(KEYINPUT2), .ZN(n633) );
  NAND2_X1 U701 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U702 ( .A1(n636), .A2(n635), .ZN(n638) );
  NOR2_X1 U703 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U704 ( .A(n639), .B(KEYINPUT81), .ZN(n680) );
  NOR2_X1 U705 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U706 ( .A(n642), .B(KEYINPUT49), .ZN(n643) );
  NAND2_X1 U707 ( .A1(n540), .A2(n643), .ZN(n647) );
  NAND2_X1 U708 ( .A1(n600), .A2(n644), .ZN(n645) );
  XOR2_X1 U709 ( .A(KEYINPUT50), .B(n645), .Z(n646) );
  NOR2_X1 U710 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U711 ( .A(n648), .B(KEYINPUT119), .ZN(n650) );
  NAND2_X1 U712 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U713 ( .A(KEYINPUT51), .B(n651), .Z(n652) );
  NAND2_X1 U714 ( .A1(n652), .A2(n675), .ZN(n669) );
  NAND2_X1 U715 ( .A1(n664), .A2(KEYINPUT120), .ZN(n655) );
  NAND2_X1 U716 ( .A1(n659), .A2(n653), .ZN(n654) );
  NAND2_X1 U717 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U718 ( .A1(n656), .A2(n657), .ZN(n666) );
  NOR2_X1 U719 ( .A1(KEYINPUT120), .A2(n657), .ZN(n658) );
  NOR2_X1 U720 ( .A1(n659), .A2(n658), .ZN(n662) );
  INV_X1 U721 ( .A(n659), .ZN(n660) );
  NOR2_X1 U722 ( .A1(KEYINPUT120), .A2(n660), .ZN(n661) );
  NOR2_X1 U723 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U724 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U725 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U726 ( .A1(n667), .A2(n674), .ZN(n668) );
  NAND2_X1 U727 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U728 ( .A(n670), .B(KEYINPUT121), .ZN(n671) );
  XOR2_X1 U729 ( .A(n671), .B(KEYINPUT52), .Z(n673) );
  AND2_X1 U730 ( .A1(n673), .A2(n672), .ZN(n678) );
  NAND2_X1 U731 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U732 ( .A1(n676), .A2(n354), .ZN(n677) );
  NOR2_X1 U733 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U734 ( .A1(n680), .A2(n679), .ZN(n682) );
  XOR2_X1 U735 ( .A(KEYINPUT122), .B(KEYINPUT53), .Z(n681) );
  XNOR2_X1 U736 ( .A(n682), .B(n681), .ZN(G75) );
  XNOR2_X1 U737 ( .A(n683), .B(G140), .ZN(G42) );
  NAND2_X1 U738 ( .A1(n698), .A2(G475), .ZN(n687) );
  XNOR2_X1 U739 ( .A(KEYINPUT87), .B(KEYINPUT59), .ZN(n684) );
  XNOR2_X1 U740 ( .A(n687), .B(n686), .ZN(n688) );
  NOR2_X2 U741 ( .A1(n688), .A2(n715), .ZN(n689) );
  XNOR2_X1 U742 ( .A(n689), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U743 ( .A1(n698), .A2(G210), .ZN(n694) );
  XOR2_X1 U744 ( .A(KEYINPUT86), .B(KEYINPUT54), .Z(n691) );
  XNOR2_X1 U745 ( .A(n691), .B(KEYINPUT55), .ZN(n692) );
  XNOR2_X1 U746 ( .A(n694), .B(n693), .ZN(n695) );
  XOR2_X1 U747 ( .A(KEYINPUT123), .B(KEYINPUT56), .Z(n696) );
  XNOR2_X1 U748 ( .A(n697), .B(n696), .ZN(G51) );
  NAND2_X1 U749 ( .A1(n698), .A2(G472), .ZN(n701) );
  XNOR2_X1 U750 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X2 U751 ( .A1(n702), .A2(n715), .ZN(n704) );
  XNOR2_X1 U752 ( .A(KEYINPUT115), .B(KEYINPUT63), .ZN(n703) );
  XNOR2_X1 U753 ( .A(n704), .B(n703), .ZN(G57) );
  BUF_X1 U754 ( .A(n705), .Z(n706) );
  XNOR2_X1 U755 ( .A(n706), .B(G110), .ZN(G12) );
  NAND2_X1 U756 ( .A1(n353), .A2(G478), .ZN(n709) );
  XNOR2_X1 U757 ( .A(n707), .B(KEYINPUT124), .ZN(n708) );
  XNOR2_X1 U758 ( .A(n709), .B(n708), .ZN(n710) );
  NOR2_X1 U759 ( .A1(n710), .A2(n715), .ZN(G63) );
  NAND2_X1 U760 ( .A1(n353), .A2(G469), .ZN(n714) );
  XNOR2_X1 U761 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n711) );
  XNOR2_X1 U762 ( .A(n712), .B(n711), .ZN(n713) );
  XNOR2_X1 U763 ( .A(n714), .B(n713), .ZN(n716) );
  NOR2_X1 U764 ( .A1(n716), .A2(n715), .ZN(G54) );
  XNOR2_X1 U765 ( .A(G101), .B(n717), .ZN(G3) );
  NOR2_X1 U766 ( .A1(n728), .A2(n719), .ZN(n718) );
  XOR2_X1 U767 ( .A(G104), .B(n718), .Z(G6) );
  NOR2_X1 U768 ( .A1(n731), .A2(n719), .ZN(n721) );
  XNOR2_X1 U769 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n720) );
  XNOR2_X1 U770 ( .A(n721), .B(n720), .ZN(n722) );
  XNOR2_X1 U771 ( .A(G107), .B(n722), .ZN(G9) );
  XNOR2_X1 U772 ( .A(n723), .B(KEYINPUT116), .ZN(n724) );
  XNOR2_X1 U773 ( .A(n724), .B(KEYINPUT29), .ZN(n725) );
  XNOR2_X1 U774 ( .A(G128), .B(n725), .ZN(G30) );
  XNOR2_X1 U775 ( .A(G146), .B(n726), .ZN(n727) );
  XNOR2_X1 U776 ( .A(n727), .B(KEYINPUT117), .ZN(G48) );
  NOR2_X1 U777 ( .A1(n728), .A2(n730), .ZN(n729) );
  XOR2_X1 U778 ( .A(G113), .B(n729), .Z(G15) );
  NOR2_X1 U779 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U780 ( .A(KEYINPUT118), .B(n732), .Z(n733) );
  XNOR2_X1 U781 ( .A(G116), .B(n733), .ZN(G18) );
  XOR2_X1 U782 ( .A(G125), .B(KEYINPUT37), .Z(n734) );
  XNOR2_X1 U783 ( .A(n735), .B(n734), .ZN(G27) );
  XNOR2_X1 U784 ( .A(G134), .B(n736), .ZN(G36) );
  XNOR2_X1 U785 ( .A(n737), .B(G101), .ZN(n738) );
  XNOR2_X1 U786 ( .A(n739), .B(n738), .ZN(n741) );
  NOR2_X1 U787 ( .A1(n354), .A2(G898), .ZN(n740) );
  NOR2_X1 U788 ( .A1(n741), .A2(n740), .ZN(n750) );
  BUF_X1 U789 ( .A(n742), .Z(n743) );
  NAND2_X1 U790 ( .A1(n743), .A2(n354), .ZN(n744) );
  XOR2_X1 U791 ( .A(KEYINPUT125), .B(n744), .Z(n748) );
  NAND2_X1 U792 ( .A1(n355), .A2(G224), .ZN(n745) );
  XNOR2_X1 U793 ( .A(KEYINPUT61), .B(n745), .ZN(n746) );
  NAND2_X1 U794 ( .A1(n746), .A2(G898), .ZN(n747) );
  NAND2_X1 U795 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U796 ( .A(n750), .B(n749), .ZN(G69) );
  XOR2_X1 U797 ( .A(G122), .B(n751), .Z(G24) );
  XNOR2_X1 U798 ( .A(G143), .B(n752), .ZN(G45) );
  XNOR2_X1 U799 ( .A(G137), .B(n753), .ZN(G39) );
  XNOR2_X1 U800 ( .A(G131), .B(n754), .ZN(G33) );
endmodule

