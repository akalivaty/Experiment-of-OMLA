

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U554 ( .A1(n683), .A2(n682), .ZN(n726) );
  INV_X1 U555 ( .A(n726), .ZN(n709) );
  BUF_X1 U556 ( .A(n570), .Z(n571) );
  XNOR2_X1 U557 ( .A(n521), .B(KEYINPUT17), .ZN(n570) );
  INV_X1 U558 ( .A(G2105), .ZN(n522) );
  NOR2_X1 U559 ( .A1(n721), .A2(n720), .ZN(n723) );
  XNOR2_X1 U560 ( .A(n708), .B(n707), .ZN(n714) );
  INV_X1 U561 ( .A(KEYINPUT95), .ZN(n750) );
  NOR2_X1 U562 ( .A1(n735), .A2(n716), .ZN(n517) );
  XNOR2_X1 U563 ( .A(n587), .B(KEYINPUT13), .ZN(n518) );
  INV_X1 U564 ( .A(G8), .ZN(n716) );
  AND2_X1 U565 ( .A1(n736), .A2(n517), .ZN(n717) );
  INV_X1 U566 ( .A(KEYINPUT29), .ZN(n706) );
  XNOR2_X1 U567 ( .A(n706), .B(KEYINPUT94), .ZN(n707) );
  INV_X1 U568 ( .A(KEYINPUT31), .ZN(n722) );
  NAND2_X1 U569 ( .A1(n733), .A2(G8), .ZN(n734) );
  NAND2_X1 U570 ( .A1(G8), .A2(n726), .ZN(n727) );
  NOR2_X1 U571 ( .A1(G1384), .A2(G164), .ZN(n680) );
  NOR2_X1 U572 ( .A1(n795), .A2(n794), .ZN(n796) );
  NOR2_X1 U573 ( .A1(G543), .A2(G651), .ZN(n646) );
  NOR2_X1 U574 ( .A1(G651), .A2(n624), .ZN(n649) );
  NOR2_X1 U575 ( .A1(n591), .A2(n590), .ZN(n986) );
  AND2_X1 U576 ( .A1(n528), .A2(n527), .ZN(G164) );
  NOR2_X2 U577 ( .A1(G2104), .A2(n522), .ZN(n860) );
  NAND2_X1 U578 ( .A1(G126), .A2(n860), .ZN(n520) );
  AND2_X1 U579 ( .A1(G2105), .A2(G2104), .ZN(n861) );
  NAND2_X1 U580 ( .A1(G114), .A2(n861), .ZN(n519) );
  AND2_X1 U581 ( .A1(n520), .A2(n519), .ZN(n528) );
  OR2_X1 U582 ( .A1(G2105), .A2(G2104), .ZN(n521) );
  NAND2_X1 U583 ( .A1(G138), .A2(n570), .ZN(n525) );
  NAND2_X1 U584 ( .A1(n522), .A2(G2104), .ZN(n523) );
  XNOR2_X1 U585 ( .A(n523), .B(KEYINPUT65), .ZN(n572) );
  NAND2_X1 U586 ( .A1(G102), .A2(n572), .ZN(n524) );
  NAND2_X1 U587 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U588 ( .A(KEYINPUT79), .B(n526), .ZN(n527) );
  NAND2_X1 U589 ( .A1(n646), .A2(G89), .ZN(n529) );
  XNOR2_X1 U590 ( .A(n529), .B(KEYINPUT4), .ZN(n532) );
  XOR2_X1 U591 ( .A(G543), .B(KEYINPUT0), .Z(n624) );
  XOR2_X1 U592 ( .A(KEYINPUT66), .B(G651), .Z(n534) );
  OR2_X1 U593 ( .A1(n624), .A2(n534), .ZN(n530) );
  XNOR2_X2 U594 ( .A(n530), .B(KEYINPUT67), .ZN(n645) );
  NAND2_X1 U595 ( .A1(G76), .A2(n645), .ZN(n531) );
  NAND2_X1 U596 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U597 ( .A(n533), .B(KEYINPUT5), .ZN(n540) );
  NAND2_X1 U598 ( .A1(G51), .A2(n649), .ZN(n537) );
  NOR2_X1 U599 ( .A1(G543), .A2(n534), .ZN(n535) );
  XOR2_X2 U600 ( .A(KEYINPUT1), .B(n535), .Z(n650) );
  NAND2_X1 U601 ( .A1(G63), .A2(n650), .ZN(n536) );
  NAND2_X1 U602 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U603 ( .A(KEYINPUT6), .B(n538), .Z(n539) );
  NAND2_X1 U604 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U605 ( .A(n541), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U606 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U607 ( .A1(G125), .A2(n860), .ZN(n543) );
  NAND2_X1 U608 ( .A1(G113), .A2(n861), .ZN(n542) );
  NAND2_X1 U609 ( .A1(n543), .A2(n542), .ZN(n548) );
  NAND2_X1 U610 ( .A1(G101), .A2(n572), .ZN(n544) );
  XOR2_X1 U611 ( .A(KEYINPUT23), .B(n544), .Z(n546) );
  NAND2_X1 U612 ( .A1(n570), .A2(G137), .ZN(n545) );
  NAND2_X1 U613 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X2 U614 ( .A1(n548), .A2(n547), .ZN(G160) );
  NAND2_X1 U615 ( .A1(G52), .A2(n649), .ZN(n550) );
  NAND2_X1 U616 ( .A1(G64), .A2(n650), .ZN(n549) );
  NAND2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n555) );
  NAND2_X1 U618 ( .A1(G77), .A2(n645), .ZN(n552) );
  NAND2_X1 U619 ( .A1(G90), .A2(n646), .ZN(n551) );
  NAND2_X1 U620 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U621 ( .A(KEYINPUT9), .B(n553), .Z(n554) );
  NOR2_X1 U622 ( .A1(n555), .A2(n554), .ZN(G171) );
  XOR2_X1 U623 ( .A(G2438), .B(G2435), .Z(n557) );
  XNOR2_X1 U624 ( .A(G2430), .B(G2454), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n557), .B(n556), .ZN(n561) );
  XOR2_X1 U626 ( .A(G2427), .B(G2443), .Z(n559) );
  XNOR2_X1 U627 ( .A(KEYINPUT101), .B(G2446), .ZN(n558) );
  XNOR2_X1 U628 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U629 ( .A(n561), .B(n560), .Z(n563) );
  XNOR2_X1 U630 ( .A(KEYINPUT100), .B(G2451), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n563), .B(n562), .ZN(n566) );
  XOR2_X1 U632 ( .A(G1348), .B(G1341), .Z(n564) );
  XNOR2_X1 U633 ( .A(KEYINPUT102), .B(n564), .ZN(n565) );
  XOR2_X1 U634 ( .A(n566), .B(n565), .Z(n567) );
  AND2_X1 U635 ( .A1(G14), .A2(n567), .ZN(G401) );
  AND2_X1 U636 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U637 ( .A1(n860), .A2(G123), .ZN(n569) );
  XNOR2_X1 U638 ( .A(KEYINPUT18), .B(KEYINPUT74), .ZN(n568) );
  XNOR2_X1 U639 ( .A(n569), .B(n568), .ZN(n579) );
  NAND2_X1 U640 ( .A1(G135), .A2(n571), .ZN(n574) );
  BUF_X1 U641 ( .A(n572), .Z(n866) );
  NAND2_X1 U642 ( .A1(G99), .A2(n866), .ZN(n573) );
  NAND2_X1 U643 ( .A1(n574), .A2(n573), .ZN(n577) );
  NAND2_X1 U644 ( .A1(G111), .A2(n861), .ZN(n575) );
  XNOR2_X1 U645 ( .A(KEYINPUT75), .B(n575), .ZN(n576) );
  NOR2_X1 U646 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U647 ( .A1(n579), .A2(n578), .ZN(n938) );
  XNOR2_X1 U648 ( .A(G2096), .B(n938), .ZN(n580) );
  OR2_X1 U649 ( .A1(G2100), .A2(n580), .ZN(G156) );
  INV_X1 U650 ( .A(G57), .ZN(G237) );
  INV_X1 U651 ( .A(G132), .ZN(G219) );
  INV_X1 U652 ( .A(G82), .ZN(G220) );
  XOR2_X1 U653 ( .A(KEYINPUT10), .B(KEYINPUT69), .Z(n582) );
  NAND2_X1 U654 ( .A1(G7), .A2(G661), .ZN(n581) );
  XNOR2_X1 U655 ( .A(n582), .B(n581), .ZN(G223) );
  INV_X1 U656 ( .A(G223), .ZN(n817) );
  NAND2_X1 U657 ( .A1(n817), .A2(G567), .ZN(n583) );
  XOR2_X1 U658 ( .A(KEYINPUT11), .B(n583), .Z(G234) );
  NAND2_X1 U659 ( .A1(n646), .A2(G81), .ZN(n584) );
  XNOR2_X1 U660 ( .A(n584), .B(KEYINPUT12), .ZN(n586) );
  NAND2_X1 U661 ( .A1(G68), .A2(n645), .ZN(n585) );
  NAND2_X1 U662 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U663 ( .A1(G43), .A2(n649), .ZN(n588) );
  NAND2_X1 U664 ( .A1(n518), .A2(n588), .ZN(n591) );
  NAND2_X1 U665 ( .A1(n650), .A2(G56), .ZN(n589) );
  XOR2_X1 U666 ( .A(KEYINPUT14), .B(n589), .Z(n590) );
  NAND2_X1 U667 ( .A1(n986), .A2(G860), .ZN(G153) );
  XOR2_X1 U668 ( .A(G171), .B(KEYINPUT70), .Z(G301) );
  NAND2_X1 U669 ( .A1(G868), .A2(G301), .ZN(n603) );
  NAND2_X1 U670 ( .A1(G92), .A2(n646), .ZN(n599) );
  NAND2_X1 U671 ( .A1(G79), .A2(n645), .ZN(n593) );
  NAND2_X1 U672 ( .A1(G54), .A2(n649), .ZN(n592) );
  NAND2_X1 U673 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U674 ( .A(KEYINPUT72), .B(n594), .ZN(n597) );
  NAND2_X1 U675 ( .A1(G66), .A2(n650), .ZN(n595) );
  XNOR2_X1 U676 ( .A(KEYINPUT71), .B(n595), .ZN(n596) );
  NOR2_X1 U677 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U678 ( .A1(n599), .A2(n598), .ZN(n601) );
  XOR2_X1 U679 ( .A(KEYINPUT73), .B(KEYINPUT15), .Z(n600) );
  XNOR2_X1 U680 ( .A(n601), .B(n600), .ZN(n882) );
  INV_X1 U681 ( .A(n882), .ZN(n983) );
  INV_X1 U682 ( .A(G868), .ZN(n662) );
  NAND2_X1 U683 ( .A1(n983), .A2(n662), .ZN(n602) );
  NAND2_X1 U684 ( .A1(n603), .A2(n602), .ZN(G284) );
  NAND2_X1 U685 ( .A1(G78), .A2(n645), .ZN(n605) );
  NAND2_X1 U686 ( .A1(G53), .A2(n649), .ZN(n604) );
  NAND2_X1 U687 ( .A1(n605), .A2(n604), .ZN(n609) );
  NAND2_X1 U688 ( .A1(G91), .A2(n646), .ZN(n607) );
  NAND2_X1 U689 ( .A1(G65), .A2(n650), .ZN(n606) );
  NAND2_X1 U690 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U691 ( .A1(n609), .A2(n608), .ZN(n985) );
  INV_X1 U692 ( .A(n985), .ZN(G299) );
  NOR2_X1 U693 ( .A1(G286), .A2(n662), .ZN(n611) );
  NOR2_X1 U694 ( .A1(G868), .A2(G299), .ZN(n610) );
  NOR2_X1 U695 ( .A1(n611), .A2(n610), .ZN(G297) );
  INV_X1 U696 ( .A(G860), .ZN(n898) );
  NAND2_X1 U697 ( .A1(n898), .A2(G559), .ZN(n612) );
  NAND2_X1 U698 ( .A1(n612), .A2(n882), .ZN(n613) );
  XNOR2_X1 U699 ( .A(n613), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U700 ( .A1(n882), .A2(G868), .ZN(n614) );
  NOR2_X1 U701 ( .A1(G559), .A2(n614), .ZN(n616) );
  AND2_X1 U702 ( .A1(n662), .A2(n986), .ZN(n615) );
  NOR2_X1 U703 ( .A1(n616), .A2(n615), .ZN(G282) );
  NAND2_X1 U704 ( .A1(G47), .A2(n649), .ZN(n618) );
  NAND2_X1 U705 ( .A1(G60), .A2(n650), .ZN(n617) );
  NAND2_X1 U706 ( .A1(n618), .A2(n617), .ZN(n621) );
  NAND2_X1 U707 ( .A1(G72), .A2(n645), .ZN(n619) );
  XOR2_X1 U708 ( .A(KEYINPUT68), .B(n619), .Z(n620) );
  NOR2_X1 U709 ( .A1(n621), .A2(n620), .ZN(n623) );
  NAND2_X1 U710 ( .A1(n646), .A2(G85), .ZN(n622) );
  NAND2_X1 U711 ( .A1(n623), .A2(n622), .ZN(G290) );
  NAND2_X1 U712 ( .A1(G87), .A2(n624), .ZN(n626) );
  NAND2_X1 U713 ( .A1(G74), .A2(G651), .ZN(n625) );
  NAND2_X1 U714 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U715 ( .A1(n650), .A2(n627), .ZN(n629) );
  NAND2_X1 U716 ( .A1(n649), .A2(G49), .ZN(n628) );
  NAND2_X1 U717 ( .A1(n629), .A2(n628), .ZN(G288) );
  NAND2_X1 U718 ( .A1(G88), .A2(n646), .ZN(n631) );
  NAND2_X1 U719 ( .A1(G50), .A2(n649), .ZN(n630) );
  NAND2_X1 U720 ( .A1(n631), .A2(n630), .ZN(n635) );
  NAND2_X1 U721 ( .A1(G75), .A2(n645), .ZN(n633) );
  NAND2_X1 U722 ( .A1(G62), .A2(n650), .ZN(n632) );
  NAND2_X1 U723 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U724 ( .A1(n635), .A2(n634), .ZN(G166) );
  NAND2_X1 U725 ( .A1(G86), .A2(n646), .ZN(n637) );
  NAND2_X1 U726 ( .A1(G48), .A2(n649), .ZN(n636) );
  NAND2_X1 U727 ( .A1(n637), .A2(n636), .ZN(n641) );
  NAND2_X1 U728 ( .A1(G73), .A2(n645), .ZN(n638) );
  XNOR2_X1 U729 ( .A(n638), .B(KEYINPUT77), .ZN(n639) );
  XNOR2_X1 U730 ( .A(n639), .B(KEYINPUT2), .ZN(n640) );
  NOR2_X1 U731 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U732 ( .A1(n650), .A2(G61), .ZN(n642) );
  NAND2_X1 U733 ( .A1(n643), .A2(n642), .ZN(G305) );
  XNOR2_X1 U734 ( .A(KEYINPUT19), .B(G290), .ZN(n644) );
  XNOR2_X1 U735 ( .A(n644), .B(G288), .ZN(n656) );
  NAND2_X1 U736 ( .A1(G80), .A2(n645), .ZN(n648) );
  NAND2_X1 U737 ( .A1(G93), .A2(n646), .ZN(n647) );
  NAND2_X1 U738 ( .A1(n648), .A2(n647), .ZN(n654) );
  NAND2_X1 U739 ( .A1(G55), .A2(n649), .ZN(n652) );
  NAND2_X1 U740 ( .A1(G67), .A2(n650), .ZN(n651) );
  NAND2_X1 U741 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U742 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U743 ( .A(KEYINPUT76), .B(n655), .Z(n899) );
  XOR2_X1 U744 ( .A(n656), .B(n899), .Z(n658) );
  XNOR2_X1 U745 ( .A(n985), .B(G166), .ZN(n657) );
  XNOR2_X1 U746 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U747 ( .A(n659), .B(G305), .ZN(n883) );
  NAND2_X1 U748 ( .A1(G559), .A2(n882), .ZN(n660) );
  XNOR2_X1 U749 ( .A(n660), .B(n986), .ZN(n897) );
  XOR2_X1 U750 ( .A(n883), .B(n897), .Z(n661) );
  NOR2_X1 U751 ( .A1(n662), .A2(n661), .ZN(n664) );
  NOR2_X1 U752 ( .A1(n899), .A2(G868), .ZN(n663) );
  NOR2_X1 U753 ( .A1(n664), .A2(n663), .ZN(G295) );
  NAND2_X1 U754 ( .A1(G2078), .A2(G2084), .ZN(n665) );
  XOR2_X1 U755 ( .A(KEYINPUT20), .B(n665), .Z(n666) );
  NAND2_X1 U756 ( .A1(G2090), .A2(n666), .ZN(n667) );
  XNOR2_X1 U757 ( .A(KEYINPUT21), .B(n667), .ZN(n668) );
  NAND2_X1 U758 ( .A1(n668), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U759 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U760 ( .A1(G220), .A2(G219), .ZN(n669) );
  XOR2_X1 U761 ( .A(KEYINPUT22), .B(n669), .Z(n670) );
  NOR2_X1 U762 ( .A1(G218), .A2(n670), .ZN(n671) );
  NAND2_X1 U763 ( .A1(G96), .A2(n671), .ZN(n902) );
  NAND2_X1 U764 ( .A1(n902), .A2(G2106), .ZN(n676) );
  NAND2_X1 U765 ( .A1(G108), .A2(G120), .ZN(n672) );
  NOR2_X1 U766 ( .A1(G237), .A2(n672), .ZN(n673) );
  NAND2_X1 U767 ( .A1(n673), .A2(G69), .ZN(n674) );
  XNOR2_X1 U768 ( .A(n674), .B(KEYINPUT78), .ZN(n901) );
  NAND2_X1 U769 ( .A1(n901), .A2(G567), .ZN(n675) );
  NAND2_X1 U770 ( .A1(n676), .A2(n675), .ZN(n822) );
  NAND2_X1 U771 ( .A1(G483), .A2(G661), .ZN(n677) );
  NOR2_X1 U772 ( .A1(n822), .A2(n677), .ZN(n821) );
  NAND2_X1 U773 ( .A1(n821), .A2(G36), .ZN(G176) );
  INV_X1 U774 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U775 ( .A(G1986), .B(KEYINPUT80), .ZN(n678) );
  XNOR2_X1 U776 ( .A(n678), .B(G290), .ZN(n1009) );
  NAND2_X1 U777 ( .A1(G40), .A2(G160), .ZN(n679) );
  XNOR2_X1 U778 ( .A(KEYINPUT81), .B(n679), .ZN(n683) );
  INV_X1 U779 ( .A(n683), .ZN(n681) );
  XNOR2_X1 U780 ( .A(n680), .B(KEYINPUT64), .ZN(n682) );
  NOR2_X1 U781 ( .A1(n681), .A2(n682), .ZN(n810) );
  NAND2_X1 U782 ( .A1(n1009), .A2(n810), .ZN(n797) );
  NAND2_X1 U783 ( .A1(G1996), .A2(n709), .ZN(n684) );
  XNOR2_X1 U784 ( .A(KEYINPUT26), .B(n684), .ZN(n685) );
  NAND2_X1 U785 ( .A1(n685), .A2(n986), .ZN(n688) );
  NAND2_X1 U786 ( .A1(G1341), .A2(n726), .ZN(n686) );
  XNOR2_X1 U787 ( .A(KEYINPUT93), .B(n686), .ZN(n687) );
  NOR2_X1 U788 ( .A1(n688), .A2(n687), .ZN(n693) );
  NAND2_X1 U789 ( .A1(n693), .A2(n882), .ZN(n692) );
  NAND2_X1 U790 ( .A1(G1348), .A2(n726), .ZN(n690) );
  NAND2_X1 U791 ( .A1(G2067), .A2(n709), .ZN(n689) );
  NAND2_X1 U792 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U793 ( .A1(n692), .A2(n691), .ZN(n695) );
  OR2_X1 U794 ( .A1(n693), .A2(n882), .ZN(n694) );
  NAND2_X1 U795 ( .A1(n695), .A2(n694), .ZN(n701) );
  NAND2_X1 U796 ( .A1(G2072), .A2(n709), .ZN(n697) );
  XNOR2_X1 U797 ( .A(KEYINPUT27), .B(KEYINPUT92), .ZN(n696) );
  XNOR2_X1 U798 ( .A(n697), .B(n696), .ZN(n699) );
  INV_X1 U799 ( .A(G1956), .ZN(n913) );
  NOR2_X1 U800 ( .A1(n709), .A2(n913), .ZN(n698) );
  NOR2_X1 U801 ( .A1(n699), .A2(n698), .ZN(n702) );
  NAND2_X1 U802 ( .A1(n702), .A2(n985), .ZN(n700) );
  NAND2_X1 U803 ( .A1(n701), .A2(n700), .ZN(n705) );
  NOR2_X1 U804 ( .A1(n702), .A2(n985), .ZN(n703) );
  XOR2_X1 U805 ( .A(n703), .B(KEYINPUT28), .Z(n704) );
  NAND2_X1 U806 ( .A1(n705), .A2(n704), .ZN(n708) );
  XOR2_X1 U807 ( .A(G1961), .B(KEYINPUT90), .Z(n911) );
  NAND2_X1 U808 ( .A1(n911), .A2(n726), .ZN(n711) );
  XNOR2_X1 U809 ( .A(KEYINPUT25), .B(G2078), .ZN(n965) );
  NAND2_X1 U810 ( .A1(n709), .A2(n965), .ZN(n710) );
  NAND2_X1 U811 ( .A1(n711), .A2(n710), .ZN(n719) );
  NAND2_X1 U812 ( .A1(G171), .A2(n719), .ZN(n712) );
  XOR2_X1 U813 ( .A(KEYINPUT91), .B(n712), .Z(n713) );
  NAND2_X1 U814 ( .A1(n714), .A2(n713), .ZN(n725) );
  NOR2_X1 U815 ( .A1(n727), .A2(G1966), .ZN(n715) );
  XNOR2_X1 U816 ( .A(n715), .B(KEYINPUT89), .ZN(n736) );
  NOR2_X1 U817 ( .A1(G2084), .A2(n726), .ZN(n735) );
  XOR2_X1 U818 ( .A(KEYINPUT30), .B(n717), .Z(n718) );
  NOR2_X1 U819 ( .A1(G168), .A2(n718), .ZN(n721) );
  NOR2_X1 U820 ( .A1(G171), .A2(n719), .ZN(n720) );
  XNOR2_X1 U821 ( .A(n723), .B(n722), .ZN(n724) );
  NAND2_X1 U822 ( .A1(n725), .A2(n724), .ZN(n737) );
  NAND2_X1 U823 ( .A1(n737), .A2(G286), .ZN(n732) );
  NOR2_X1 U824 ( .A1(G2090), .A2(n726), .ZN(n729) );
  NOR2_X1 U825 ( .A1(G1971), .A2(n727), .ZN(n728) );
  NOR2_X1 U826 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U827 ( .A1(n730), .A2(G303), .ZN(n731) );
  NAND2_X1 U828 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U829 ( .A(n734), .B(KEYINPUT32), .ZN(n741) );
  NAND2_X1 U830 ( .A1(G8), .A2(n735), .ZN(n739) );
  AND2_X1 U831 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U832 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U833 ( .A1(n741), .A2(n740), .ZN(n755) );
  NOR2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n989) );
  NOR2_X1 U835 ( .A1(G1971), .A2(G303), .ZN(n995) );
  NOR2_X1 U836 ( .A1(n989), .A2(n995), .ZN(n742) );
  NAND2_X1 U837 ( .A1(n755), .A2(n742), .ZN(n743) );
  NAND2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n990) );
  NAND2_X1 U839 ( .A1(n743), .A2(n990), .ZN(n744) );
  NOR2_X1 U840 ( .A1(KEYINPUT33), .A2(n744), .ZN(n745) );
  INV_X1 U841 ( .A(n727), .ZN(n746) );
  NAND2_X1 U842 ( .A1(n745), .A2(n746), .ZN(n749) );
  NAND2_X1 U843 ( .A1(n989), .A2(n746), .ZN(n747) );
  NAND2_X1 U844 ( .A1(n747), .A2(KEYINPUT33), .ZN(n748) );
  NAND2_X1 U845 ( .A1(n749), .A2(n748), .ZN(n751) );
  XNOR2_X1 U846 ( .A(n751), .B(n750), .ZN(n752) );
  XOR2_X1 U847 ( .A(G1981), .B(G305), .Z(n1004) );
  NAND2_X1 U848 ( .A1(n752), .A2(n1004), .ZN(n758) );
  NOR2_X1 U849 ( .A1(G2090), .A2(G303), .ZN(n753) );
  NAND2_X1 U850 ( .A1(G8), .A2(n753), .ZN(n754) );
  NAND2_X1 U851 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U852 ( .A1(n756), .A2(n727), .ZN(n757) );
  NAND2_X1 U853 ( .A1(n758), .A2(n757), .ZN(n762) );
  NOR2_X1 U854 ( .A1(G1981), .A2(G305), .ZN(n759) );
  XOR2_X1 U855 ( .A(n759), .B(KEYINPUT24), .Z(n760) );
  NOR2_X1 U856 ( .A1(n727), .A2(n760), .ZN(n761) );
  NOR2_X1 U857 ( .A1(n762), .A2(n761), .ZN(n795) );
  XNOR2_X1 U858 ( .A(G2067), .B(KEYINPUT37), .ZN(n763) );
  XOR2_X1 U859 ( .A(n763), .B(KEYINPUT82), .Z(n807) );
  NAND2_X1 U860 ( .A1(G140), .A2(n571), .ZN(n765) );
  NAND2_X1 U861 ( .A1(G104), .A2(n866), .ZN(n764) );
  NAND2_X1 U862 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U863 ( .A(KEYINPUT34), .B(n766), .ZN(n771) );
  NAND2_X1 U864 ( .A1(G128), .A2(n860), .ZN(n768) );
  NAND2_X1 U865 ( .A1(G116), .A2(n861), .ZN(n767) );
  NAND2_X1 U866 ( .A1(n768), .A2(n767), .ZN(n769) );
  XOR2_X1 U867 ( .A(KEYINPUT35), .B(n769), .Z(n770) );
  NOR2_X1 U868 ( .A1(n771), .A2(n770), .ZN(n772) );
  XOR2_X1 U869 ( .A(KEYINPUT36), .B(n772), .Z(n857) );
  AND2_X1 U870 ( .A1(n807), .A2(n857), .ZN(n945) );
  NAND2_X1 U871 ( .A1(n810), .A2(n945), .ZN(n805) );
  NAND2_X1 U872 ( .A1(G129), .A2(n860), .ZN(n774) );
  NAND2_X1 U873 ( .A1(G117), .A2(n861), .ZN(n773) );
  NAND2_X1 U874 ( .A1(n774), .A2(n773), .ZN(n777) );
  NAND2_X1 U875 ( .A1(n866), .A2(G105), .ZN(n775) );
  XOR2_X1 U876 ( .A(KEYINPUT38), .B(n775), .Z(n776) );
  NOR2_X1 U877 ( .A1(n777), .A2(n776), .ZN(n779) );
  NAND2_X1 U878 ( .A1(n571), .A2(G141), .ZN(n778) );
  NAND2_X1 U879 ( .A1(n779), .A2(n778), .ZN(n876) );
  NAND2_X1 U880 ( .A1(n876), .A2(G1996), .ZN(n791) );
  NAND2_X1 U881 ( .A1(G131), .A2(n571), .ZN(n781) );
  NAND2_X1 U882 ( .A1(G95), .A2(n866), .ZN(n780) );
  NAND2_X1 U883 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U884 ( .A(n782), .B(KEYINPUT85), .ZN(n788) );
  NAND2_X1 U885 ( .A1(n860), .A2(G119), .ZN(n783) );
  XOR2_X1 U886 ( .A(KEYINPUT83), .B(n783), .Z(n785) );
  NAND2_X1 U887 ( .A1(n861), .A2(G107), .ZN(n784) );
  NAND2_X1 U888 ( .A1(n785), .A2(n784), .ZN(n786) );
  XOR2_X1 U889 ( .A(KEYINPUT84), .B(n786), .Z(n787) );
  NAND2_X1 U890 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U891 ( .A(n789), .B(KEYINPUT86), .ZN(n856) );
  NAND2_X1 U892 ( .A1(G1991), .A2(n856), .ZN(n790) );
  NAND2_X1 U893 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U894 ( .A(n792), .B(KEYINPUT87), .Z(n948) );
  NAND2_X1 U895 ( .A1(n948), .A2(n810), .ZN(n798) );
  NAND2_X1 U896 ( .A1(n805), .A2(n798), .ZN(n793) );
  XNOR2_X1 U897 ( .A(n793), .B(KEYINPUT88), .ZN(n794) );
  NAND2_X1 U898 ( .A1(n797), .A2(n796), .ZN(n813) );
  NOR2_X1 U899 ( .A1(G1996), .A2(n876), .ZN(n936) );
  INV_X1 U900 ( .A(n798), .ZN(n801) );
  NOR2_X1 U901 ( .A1(G1986), .A2(G290), .ZN(n799) );
  NOR2_X1 U902 ( .A1(G1991), .A2(n856), .ZN(n941) );
  NOR2_X1 U903 ( .A1(n799), .A2(n941), .ZN(n800) );
  NOR2_X1 U904 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U905 ( .A(n802), .B(KEYINPUT96), .ZN(n803) );
  NOR2_X1 U906 ( .A1(n936), .A2(n803), .ZN(n804) );
  XNOR2_X1 U907 ( .A(n804), .B(KEYINPUT39), .ZN(n806) );
  NAND2_X1 U908 ( .A1(n806), .A2(n805), .ZN(n809) );
  NOR2_X1 U909 ( .A1(n807), .A2(n857), .ZN(n808) );
  XNOR2_X1 U910 ( .A(n808), .B(KEYINPUT97), .ZN(n949) );
  NAND2_X1 U911 ( .A1(n809), .A2(n949), .ZN(n811) );
  NAND2_X1 U912 ( .A1(n811), .A2(n810), .ZN(n812) );
  NAND2_X1 U913 ( .A1(n813), .A2(n812), .ZN(n816) );
  XOR2_X1 U914 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n814) );
  XNOR2_X1 U915 ( .A(KEYINPUT40), .B(n814), .ZN(n815) );
  XNOR2_X1 U916 ( .A(n816), .B(n815), .ZN(G329) );
  NAND2_X1 U917 ( .A1(G2106), .A2(n817), .ZN(G217) );
  AND2_X1 U918 ( .A1(G15), .A2(G2), .ZN(n818) );
  NAND2_X1 U919 ( .A1(G661), .A2(n818), .ZN(G259) );
  NAND2_X1 U920 ( .A1(G3), .A2(G1), .ZN(n819) );
  XOR2_X1 U921 ( .A(KEYINPUT103), .B(n819), .Z(n820) );
  NAND2_X1 U922 ( .A1(n821), .A2(n820), .ZN(G188) );
  XOR2_X1 U923 ( .A(G120), .B(KEYINPUT104), .Z(G236) );
  INV_X1 U924 ( .A(n822), .ZN(G319) );
  XNOR2_X1 U925 ( .A(G1996), .B(G2474), .ZN(n832) );
  XOR2_X1 U926 ( .A(G1981), .B(G1956), .Z(n824) );
  XNOR2_X1 U927 ( .A(G1991), .B(G1966), .ZN(n823) );
  XNOR2_X1 U928 ( .A(n824), .B(n823), .ZN(n828) );
  XOR2_X1 U929 ( .A(G1976), .B(G1971), .Z(n826) );
  XNOR2_X1 U930 ( .A(G1986), .B(G1961), .ZN(n825) );
  XNOR2_X1 U931 ( .A(n826), .B(n825), .ZN(n827) );
  XOR2_X1 U932 ( .A(n828), .B(n827), .Z(n830) );
  XNOR2_X1 U933 ( .A(KEYINPUT106), .B(KEYINPUT41), .ZN(n829) );
  XNOR2_X1 U934 ( .A(n830), .B(n829), .ZN(n831) );
  XNOR2_X1 U935 ( .A(n832), .B(n831), .ZN(G229) );
  XOR2_X1 U936 ( .A(G2100), .B(G2096), .Z(n834) );
  XNOR2_X1 U937 ( .A(KEYINPUT42), .B(G2678), .ZN(n833) );
  XNOR2_X1 U938 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U939 ( .A(KEYINPUT43), .B(G2090), .Z(n836) );
  XNOR2_X1 U940 ( .A(G2067), .B(G2072), .ZN(n835) );
  XNOR2_X1 U941 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U942 ( .A(n838), .B(n837), .Z(n840) );
  XNOR2_X1 U943 ( .A(G2078), .B(G2084), .ZN(n839) );
  XNOR2_X1 U944 ( .A(n840), .B(n839), .ZN(G227) );
  NAND2_X1 U945 ( .A1(n860), .A2(G124), .ZN(n841) );
  XNOR2_X1 U946 ( .A(n841), .B(KEYINPUT44), .ZN(n843) );
  NAND2_X1 U947 ( .A1(G100), .A2(n866), .ZN(n842) );
  NAND2_X1 U948 ( .A1(n843), .A2(n842), .ZN(n847) );
  NAND2_X1 U949 ( .A1(G112), .A2(n861), .ZN(n845) );
  NAND2_X1 U950 ( .A1(G136), .A2(n571), .ZN(n844) );
  NAND2_X1 U951 ( .A1(n845), .A2(n844), .ZN(n846) );
  NOR2_X1 U952 ( .A1(n847), .A2(n846), .ZN(G162) );
  NAND2_X1 U953 ( .A1(G139), .A2(n571), .ZN(n849) );
  NAND2_X1 U954 ( .A1(G103), .A2(n866), .ZN(n848) );
  NAND2_X1 U955 ( .A1(n849), .A2(n848), .ZN(n855) );
  NAND2_X1 U956 ( .A1(n861), .A2(G115), .ZN(n850) );
  XOR2_X1 U957 ( .A(KEYINPUT109), .B(n850), .Z(n852) );
  NAND2_X1 U958 ( .A1(n860), .A2(G127), .ZN(n851) );
  NAND2_X1 U959 ( .A1(n852), .A2(n851), .ZN(n853) );
  XOR2_X1 U960 ( .A(KEYINPUT47), .B(n853), .Z(n854) );
  NOR2_X1 U961 ( .A1(n855), .A2(n854), .ZN(n931) );
  XOR2_X1 U962 ( .A(n931), .B(n856), .Z(n859) );
  XNOR2_X1 U963 ( .A(G164), .B(n857), .ZN(n858) );
  XNOR2_X1 U964 ( .A(n859), .B(n858), .ZN(n873) );
  NAND2_X1 U965 ( .A1(G130), .A2(n860), .ZN(n863) );
  NAND2_X1 U966 ( .A1(G118), .A2(n861), .ZN(n862) );
  NAND2_X1 U967 ( .A1(n863), .A2(n862), .ZN(n864) );
  XOR2_X1 U968 ( .A(KEYINPUT107), .B(n864), .Z(n871) );
  NAND2_X1 U969 ( .A1(n571), .A2(G142), .ZN(n865) );
  XNOR2_X1 U970 ( .A(n865), .B(KEYINPUT108), .ZN(n868) );
  NAND2_X1 U971 ( .A1(G106), .A2(n866), .ZN(n867) );
  NAND2_X1 U972 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U973 ( .A(n869), .B(KEYINPUT45), .Z(n870) );
  NOR2_X1 U974 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U975 ( .A(n873), .B(n872), .Z(n880) );
  XOR2_X1 U976 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n875) );
  XNOR2_X1 U977 ( .A(G160), .B(G162), .ZN(n874) );
  XNOR2_X1 U978 ( .A(n875), .B(n874), .ZN(n877) );
  XOR2_X1 U979 ( .A(n877), .B(n876), .Z(n878) );
  XNOR2_X1 U980 ( .A(n938), .B(n878), .ZN(n879) );
  XNOR2_X1 U981 ( .A(n880), .B(n879), .ZN(n881) );
  NOR2_X1 U982 ( .A1(G37), .A2(n881), .ZN(G395) );
  XNOR2_X1 U983 ( .A(n882), .B(G171), .ZN(n887) );
  XOR2_X1 U984 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n885) );
  XNOR2_X1 U985 ( .A(n986), .B(n883), .ZN(n884) );
  XNOR2_X1 U986 ( .A(n885), .B(n884), .ZN(n886) );
  XNOR2_X1 U987 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U988 ( .A(n888), .B(G286), .ZN(n889) );
  NOR2_X1 U989 ( .A1(G37), .A2(n889), .ZN(G397) );
  XNOR2_X1 U990 ( .A(KEYINPUT112), .B(KEYINPUT49), .ZN(n891) );
  NOR2_X1 U991 ( .A1(G229), .A2(G227), .ZN(n890) );
  XNOR2_X1 U992 ( .A(n891), .B(n890), .ZN(n892) );
  NOR2_X1 U993 ( .A1(G401), .A2(n892), .ZN(n893) );
  NAND2_X1 U994 ( .A1(G319), .A2(n893), .ZN(n894) );
  XNOR2_X1 U995 ( .A(KEYINPUT113), .B(n894), .ZN(n896) );
  NOR2_X1 U996 ( .A1(G395), .A2(G397), .ZN(n895) );
  NAND2_X1 U997 ( .A1(n896), .A2(n895), .ZN(G225) );
  XOR2_X1 U998 ( .A(KEYINPUT114), .B(G225), .Z(G308) );
  NAND2_X1 U1000 ( .A1(n898), .A2(n897), .ZN(n900) );
  XNOR2_X1 U1001 ( .A(n900), .B(n899), .ZN(G145) );
  INV_X1 U1002 ( .A(G108), .ZN(G238) );
  INV_X1 U1003 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1004 ( .A1(n902), .A2(n901), .ZN(n903) );
  XNOR2_X1 U1005 ( .A(n903), .B(KEYINPUT105), .ZN(G261) );
  INV_X1 U1006 ( .A(G261), .ZN(G325) );
  INV_X1 U1007 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1008 ( .A(G1971), .B(G22), .ZN(n905) );
  XNOR2_X1 U1009 ( .A(G23), .B(G1976), .ZN(n904) );
  NOR2_X1 U1010 ( .A1(n905), .A2(n904), .ZN(n907) );
  XOR2_X1 U1011 ( .A(G1986), .B(G24), .Z(n906) );
  NAND2_X1 U1012 ( .A1(n907), .A2(n906), .ZN(n910) );
  XNOR2_X1 U1013 ( .A(KEYINPUT126), .B(KEYINPUT127), .ZN(n908) );
  XNOR2_X1 U1014 ( .A(n908), .B(KEYINPUT58), .ZN(n909) );
  XNOR2_X1 U1015 ( .A(n910), .B(n909), .ZN(n924) );
  XOR2_X1 U1016 ( .A(n911), .B(G5), .Z(n922) );
  XNOR2_X1 U1017 ( .A(KEYINPUT59), .B(G1348), .ZN(n912) );
  XNOR2_X1 U1018 ( .A(n912), .B(G4), .ZN(n919) );
  XOR2_X1 U1019 ( .A(G1341), .B(G19), .Z(n915) );
  XNOR2_X1 U1020 ( .A(n913), .B(G20), .ZN(n914) );
  NAND2_X1 U1021 ( .A1(n915), .A2(n914), .ZN(n917) );
  XNOR2_X1 U1022 ( .A(G6), .B(G1981), .ZN(n916) );
  NOR2_X1 U1023 ( .A1(n917), .A2(n916), .ZN(n918) );
  NAND2_X1 U1024 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1025 ( .A(n920), .B(KEYINPUT60), .ZN(n921) );
  NOR2_X1 U1026 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1027 ( .A1(n924), .A2(n923), .ZN(n926) );
  XNOR2_X1 U1028 ( .A(G21), .B(G1966), .ZN(n925) );
  NOR2_X1 U1029 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1030 ( .A(KEYINPUT61), .B(n927), .ZN(n929) );
  INV_X1 U1031 ( .A(G16), .ZN(n928) );
  NAND2_X1 U1032 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1033 ( .A1(n930), .A2(G11), .ZN(n958) );
  XOR2_X1 U1034 ( .A(G2072), .B(n931), .Z(n933) );
  XOR2_X1 U1035 ( .A(G164), .B(G2078), .Z(n932) );
  NOR2_X1 U1036 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1037 ( .A(KEYINPUT50), .B(n934), .ZN(n947) );
  XOR2_X1 U1038 ( .A(G2090), .B(G162), .Z(n935) );
  NOR2_X1 U1039 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1040 ( .A(KEYINPUT51), .B(n937), .Z(n943) );
  XNOR2_X1 U1041 ( .A(G160), .B(G2084), .ZN(n939) );
  NAND2_X1 U1042 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1043 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1044 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1045 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1046 ( .A1(n947), .A2(n946), .ZN(n952) );
  INV_X1 U1047 ( .A(n948), .ZN(n950) );
  NAND2_X1 U1048 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1049 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1050 ( .A(KEYINPUT52), .B(n953), .Z(n954) );
  NOR2_X1 U1051 ( .A1(KEYINPUT55), .A2(n954), .ZN(n956) );
  INV_X1 U1052 ( .A(G29), .ZN(n955) );
  NOR2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n982) );
  XOR2_X1 U1055 ( .A(KEYINPUT118), .B(G29), .Z(n980) );
  XOR2_X1 U1056 ( .A(G2090), .B(G35), .Z(n974) );
  XNOR2_X1 U1057 ( .A(G1991), .B(G25), .ZN(n963) );
  XNOR2_X1 U1058 ( .A(G2067), .B(G26), .ZN(n960) );
  XNOR2_X1 U1059 ( .A(G2072), .B(G33), .ZN(n959) );
  NOR2_X1 U1060 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1061 ( .A(KEYINPUT115), .B(n961), .ZN(n962) );
  NOR2_X1 U1062 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1063 ( .A1(G28), .A2(n964), .ZN(n970) );
  XOR2_X1 U1064 ( .A(G1996), .B(G32), .Z(n967) );
  XNOR2_X1 U1065 ( .A(n965), .B(G27), .ZN(n966) );
  NAND2_X1 U1066 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1067 ( .A(KEYINPUT116), .B(n968), .ZN(n969) );
  NOR2_X1 U1068 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1069 ( .A(n971), .B(KEYINPUT117), .ZN(n972) );
  XNOR2_X1 U1070 ( .A(n972), .B(KEYINPUT53), .ZN(n973) );
  NAND2_X1 U1071 ( .A1(n974), .A2(n973), .ZN(n977) );
  XNOR2_X1 U1072 ( .A(G34), .B(G2084), .ZN(n975) );
  XNOR2_X1 U1073 ( .A(KEYINPUT54), .B(n975), .ZN(n976) );
  NOR2_X1 U1074 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1075 ( .A(KEYINPUT55), .B(n978), .ZN(n979) );
  NAND2_X1 U1076 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n1018) );
  XOR2_X1 U1078 ( .A(KEYINPUT56), .B(G16), .Z(n1016) );
  XNOR2_X1 U1079 ( .A(n983), .B(G1348), .ZN(n984) );
  XNOR2_X1 U1080 ( .A(n984), .B(KEYINPUT121), .ZN(n1001) );
  XNOR2_X1 U1081 ( .A(n985), .B(G1956), .ZN(n988) );
  XNOR2_X1 U1082 ( .A(n986), .B(G1341), .ZN(n987) );
  NAND2_X1 U1083 ( .A1(n988), .A2(n987), .ZN(n999) );
  INV_X1 U1084 ( .A(n989), .ZN(n991) );
  NAND2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1086 ( .A(n992), .B(KEYINPUT123), .ZN(n994) );
  NAND2_X1 U1087 ( .A1(G1971), .A2(G303), .ZN(n993) );
  NAND2_X1 U1088 ( .A1(n994), .A2(n993), .ZN(n996) );
  NOR2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1090 ( .A(KEYINPUT124), .B(n997), .Z(n998) );
  NOR2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1013) );
  XOR2_X1 U1093 ( .A(G1966), .B(G168), .Z(n1002) );
  XNOR2_X1 U1094 ( .A(KEYINPUT119), .B(n1002), .ZN(n1003) );
  NAND2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1006) );
  XNOR2_X1 U1096 ( .A(KEYINPUT57), .B(KEYINPUT120), .ZN(n1005) );
  XNOR2_X1 U1097 ( .A(n1006), .B(n1005), .ZN(n1011) );
  XOR2_X1 U1098 ( .A(G171), .B(G1961), .Z(n1007) );
  XNOR2_X1 U1099 ( .A(KEYINPUT122), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1100 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1103 ( .A(KEYINPUT125), .B(n1014), .Z(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1106 ( .A(n1019), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

