//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 1 0 1 1 1 1 1 1 1 0 1 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 1 0 1 0 0 1 0 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n767, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068;
  INV_X1    g000(.A(KEYINPUT29), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT64), .ZN(new_n188));
  XNOR2_X1  g002(.A(G143), .B(G146), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT0), .B(G128), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n188), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(KEYINPUT0), .A2(G128), .ZN(new_n197));
  OR2_X1    g011(.A1(KEYINPUT0), .A2(G128), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n196), .A2(KEYINPUT64), .A3(new_n197), .A4(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n189), .A2(KEYINPUT0), .A3(G128), .ZN(new_n200));
  AND3_X1   g014(.A1(new_n191), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G137), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(KEYINPUT11), .A3(G134), .ZN(new_n203));
  INV_X1    g017(.A(G134), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G137), .ZN(new_n205));
  AND2_X1   g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT11), .ZN(new_n207));
  OAI211_X1 g021(.A(KEYINPUT65), .B(new_n207), .C1(new_n204), .C2(G137), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n202), .A2(G134), .ZN(new_n210));
  AOI21_X1  g024(.A(KEYINPUT65), .B1(new_n210), .B2(new_n207), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n206), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G131), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(KEYINPUT66), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n203), .A2(new_n205), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n207), .B1(new_n204), .B2(G137), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT65), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n216), .B1(new_n219), .B2(new_n208), .ZN(new_n220));
  INV_X1    g034(.A(new_n214), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n201), .B1(new_n215), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G116), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(G119), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n226));
  INV_X1    g040(.A(G119), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n226), .B1(new_n227), .B2(G116), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n224), .A2(KEYINPUT68), .A3(G119), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n225), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT2), .B(G113), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n235));
  AOI211_X1 g049(.A(new_n235), .B(new_n225), .C1(new_n228), .C2(new_n229), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n228), .A2(new_n229), .ZN(new_n237));
  INV_X1    g051(.A(new_n225), .ZN(new_n238));
  AOI21_X1  g052(.A(KEYINPUT69), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n234), .B1(new_n240), .B2(new_n231), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n213), .B1(new_n210), .B2(new_n205), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n242), .B1(new_n220), .B2(new_n213), .ZN(new_n243));
  INV_X1    g057(.A(G128), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n192), .A2(G143), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n196), .A2(new_n244), .B1(KEYINPUT1), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT1), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n193), .A2(new_n195), .A3(new_n247), .A4(G128), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n243), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n223), .A2(new_n241), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n249), .B1(new_n243), .B2(KEYINPUT67), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n206), .B(new_n213), .C1(new_n209), .C2(new_n211), .ZN(new_n254));
  INV_X1    g068(.A(new_n242), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(KEYINPUT67), .A3(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n223), .B1(new_n253), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT30), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n212), .A2(new_n214), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n220), .A2(new_n221), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n263), .A2(new_n201), .B1(new_n249), .B2(new_n243), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n241), .B1(new_n264), .B2(KEYINPUT30), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n252), .B1(new_n260), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(G237), .A2(G953), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G210), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n268), .B(KEYINPUT27), .ZN(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT26), .B(G101), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n269), .B(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n187), .B1(new_n266), .B2(new_n271), .ZN(new_n272));
  XOR2_X1   g086(.A(KEYINPUT72), .B(KEYINPUT28), .Z(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT73), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n240), .A2(new_n231), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n233), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n258), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(new_n251), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n254), .A2(new_n255), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT67), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(new_n249), .A3(new_n256), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n241), .B1(new_n283), .B2(new_n223), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n284), .A2(new_n275), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n274), .B1(new_n279), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n191), .A2(new_n199), .A3(new_n200), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n287), .B1(new_n261), .B2(new_n262), .ZN(new_n288));
  OAI22_X1  g102(.A1(new_n189), .A2(G128), .B1(new_n247), .B2(new_n195), .ZN(new_n289));
  INV_X1    g103(.A(new_n248), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n280), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(KEYINPUT74), .B1(new_n288), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT74), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n223), .A2(new_n294), .A3(new_n250), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n293), .A2(new_n241), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT28), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n271), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n272), .B1(new_n286), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G902), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n277), .B1(new_n288), .B2(new_n292), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n251), .ZN(new_n304));
  AOI21_X1  g118(.A(KEYINPUT75), .B1(new_n304), .B2(KEYINPUT28), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT75), .ZN(new_n306));
  AOI211_X1 g120(.A(new_n306), .B(new_n297), .C1(new_n303), .C2(new_n251), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n296), .A2(new_n297), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(KEYINPUT29), .A3(new_n271), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n302), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(G472), .B1(new_n301), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g126(.A1(G472), .A2(G902), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT32), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n299), .B1(new_n264), .B2(new_n241), .ZN(new_n317));
  XOR2_X1   g131(.A(KEYINPUT71), .B(KEYINPUT31), .Z(new_n318));
  AOI21_X1  g132(.A(KEYINPUT30), .B1(new_n283), .B2(new_n223), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n223), .A2(KEYINPUT30), .A3(new_n250), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n277), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n317), .B(new_n318), .C1(new_n319), .C2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT70), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT31), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n291), .B1(new_n280), .B2(new_n281), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n288), .B1(new_n325), .B2(new_n256), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n277), .B(new_n320), .C1(new_n326), .C2(KEYINPUT30), .ZN(new_n327));
  AOI211_X1 g141(.A(new_n323), .B(new_n324), .C1(new_n327), .C2(new_n317), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n317), .B1(new_n319), .B2(new_n321), .ZN(new_n329));
  AOI21_X1  g143(.A(KEYINPUT70), .B1(new_n329), .B2(KEYINPUT31), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n322), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n271), .B1(new_n286), .B2(new_n309), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n316), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n322), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n251), .A2(new_n271), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n335), .B1(new_n260), .B2(new_n265), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n323), .B1(new_n336), .B2(new_n324), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n329), .A2(KEYINPUT70), .A3(KEYINPUT31), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n334), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n252), .B1(new_n284), .B2(new_n275), .ZN(new_n340));
  OAI21_X1  g154(.A(KEYINPUT73), .B1(new_n326), .B2(new_n241), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n273), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n299), .B1(new_n342), .B2(new_n298), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n314), .B1(new_n339), .B2(new_n343), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n312), .B(new_n333), .C1(new_n344), .C2(KEYINPUT32), .ZN(new_n345));
  INV_X1    g159(.A(G217), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n346), .B1(G234), .B2(new_n302), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT16), .ZN(new_n348));
  INV_X1    g162(.A(G140), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(new_n349), .A3(G125), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT78), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n352), .A2(new_n348), .A3(new_n349), .A4(G125), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G125), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n349), .B1(new_n355), .B2(KEYINPUT77), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT77), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n357), .A2(G125), .A3(G140), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n348), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n192), .B1(new_n354), .B2(new_n359), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n357), .A2(G125), .A3(G140), .ZN(new_n361));
  AOI21_X1  g175(.A(G140), .B1(new_n357), .B2(G125), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT16), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n363), .A2(G146), .A3(new_n351), .A4(new_n353), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT23), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n366), .B1(new_n227), .B2(G128), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n244), .A2(KEYINPUT23), .A3(G119), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n227), .A2(G128), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G110), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT76), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n370), .A2(KEYINPUT76), .A3(G110), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  XOR2_X1   g189(.A(KEYINPUT24), .B(G110), .Z(new_n376));
  XNOR2_X1  g190(.A(G119), .B(G128), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n365), .A2(new_n375), .A3(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(G125), .B(G140), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n192), .ZN(new_n381));
  OAI22_X1  g195(.A1(new_n370), .A2(G110), .B1(new_n376), .B2(new_n377), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n364), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT22), .B(G137), .ZN(new_n385));
  INV_X1    g199(.A(G953), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(G221), .A3(G234), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n385), .B(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n384), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n379), .A2(new_n383), .A3(new_n388), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n302), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT79), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT25), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT79), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n390), .A2(new_n395), .A3(new_n302), .A4(new_n391), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n393), .A2(KEYINPUT80), .A3(new_n394), .A4(new_n396), .ZN(new_n397));
  OR2_X1    g211(.A1(new_n392), .A2(new_n394), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(KEYINPUT25), .B1(new_n392), .B2(KEYINPUT79), .ZN(new_n400));
  AOI21_X1  g214(.A(KEYINPUT80), .B1(new_n400), .B2(new_n396), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n347), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(KEYINPUT9), .B(G234), .ZN(new_n403));
  OAI21_X1  g217(.A(G221), .B1(new_n403), .B2(G902), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G469), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n406), .A2(new_n302), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT10), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT83), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n248), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n189), .A2(KEYINPUT83), .A3(new_n247), .A4(G128), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n246), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT3), .ZN(new_n413));
  INV_X1    g227(.A(G104), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n413), .B1(new_n414), .B2(G107), .ZN(new_n415));
  INV_X1    g229(.A(G107), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(KEYINPUT3), .A3(G104), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n415), .A2(new_n417), .B1(new_n414), .B2(G107), .ZN(new_n418));
  INV_X1    g232(.A(G101), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT82), .B1(new_n416), .B2(G104), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n416), .A2(G104), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n414), .A2(G107), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n424), .A2(KEYINPUT82), .ZN(new_n425));
  OAI21_X1  g239(.A(G101), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n420), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n408), .B1(new_n412), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT4), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n429), .B1(new_n418), .B2(new_n419), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n415), .A2(new_n417), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n424), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G101), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n432), .A2(new_n429), .A3(G101), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n201), .A3(new_n435), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n215), .A2(new_n222), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n420), .A2(new_n426), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n408), .B1(new_n246), .B2(new_n248), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n428), .A2(new_n436), .A3(new_n437), .A4(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n246), .A2(new_n410), .A3(new_n411), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n442), .A2(new_n420), .A3(new_n426), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n427), .A2(new_n291), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AND3_X1   g259(.A1(new_n445), .A2(KEYINPUT12), .A3(new_n263), .ZN(new_n446));
  AOI21_X1  g260(.A(KEYINPUT12), .B1(new_n445), .B2(new_n263), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n441), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  XOR2_X1   g262(.A(G110), .B(G140), .Z(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(KEYINPUT81), .ZN(new_n450));
  AND2_X1   g264(.A1(new_n386), .A2(G227), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n450), .B(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n441), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n428), .A2(new_n436), .A3(new_n440), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n263), .ZN(new_n456));
  AOI22_X1  g270(.A1(new_n448), .A2(new_n452), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n407), .B1(new_n457), .B2(G469), .ZN(new_n458));
  AOI22_X1  g272(.A1(new_n443), .A2(new_n408), .B1(new_n438), .B2(new_n439), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n437), .B1(new_n459), .B2(new_n436), .ZN(new_n460));
  INV_X1    g274(.A(new_n441), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n452), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n441), .B(new_n453), .C1(new_n446), .C2(new_n447), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n464), .A2(new_n406), .A3(new_n302), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n405), .B1(new_n458), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n390), .A2(new_n391), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n347), .A2(G902), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n402), .A2(new_n466), .A3(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(G214), .B1(G237), .B2(G902), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(G210), .B1(G237), .B2(G902), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n249), .A2(new_n355), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n476), .B1(new_n355), .B2(new_n287), .ZN(new_n477));
  INV_X1    g291(.A(G224), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n478), .A2(G953), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n479), .B(KEYINPUT87), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n477), .B(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(G110), .B(G122), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT86), .B(KEYINPUT6), .ZN(new_n484));
  NOR3_X1   g298(.A1(new_n236), .A2(new_n239), .A3(new_n232), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n435), .B(new_n434), .C1(new_n485), .C2(new_n234), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n420), .A2(new_n426), .A3(new_n233), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT84), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT5), .ZN(new_n489));
  AND3_X1   g303(.A1(new_n224), .A2(KEYINPUT68), .A3(G119), .ZN(new_n490));
  AOI21_X1  g304(.A(KEYINPUT68), .B1(new_n224), .B2(G119), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n238), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n235), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n230), .A2(KEYINPUT69), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n489), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(G113), .B1(new_n238), .B2(KEYINPUT5), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n487), .B(new_n488), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n486), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n496), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n499), .B1(new_n240), .B2(new_n489), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n488), .B1(new_n500), .B2(new_n487), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n483), .B(new_n484), .C1(new_n498), .C2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n487), .B1(new_n495), .B2(new_n496), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT84), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n505), .A2(new_n482), .A3(new_n486), .A4(new_n497), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT85), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(new_n507), .A3(KEYINPUT6), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n506), .A2(KEYINPUT85), .A3(KEYINPUT6), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n483), .B1(new_n498), .B2(new_n501), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n481), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n482), .B(KEYINPUT8), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n500), .A2(new_n233), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n427), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT89), .ZN(new_n518));
  AOI21_X1  g332(.A(KEYINPUT88), .B1(new_n230), .B2(KEYINPUT5), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n519), .A2(new_n496), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n230), .A2(KEYINPUT88), .A3(KEYINPUT5), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI22_X1  g336(.A1(new_n517), .A2(new_n518), .B1(new_n487), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n516), .A2(KEYINPUT89), .A3(new_n427), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n515), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(KEYINPUT7), .B1(new_n478), .B2(G953), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n477), .B(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n506), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n302), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n475), .B1(new_n513), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n495), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n234), .B1(new_n531), .B2(new_n499), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n518), .B1(new_n532), .B2(new_n438), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n522), .A2(new_n487), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n533), .A2(new_n524), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n514), .ZN(new_n536));
  INV_X1    g350(.A(new_n528), .ZN(new_n537));
  AOI21_X1  g351(.A(G902), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AOI22_X1  g352(.A1(new_n508), .A2(new_n503), .B1(new_n510), .B2(new_n511), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n538), .B(new_n474), .C1(new_n539), .C2(new_n481), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n473), .B1(new_n530), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT20), .ZN(new_n542));
  XOR2_X1   g356(.A(G113), .B(G122), .Z(new_n543));
  XOR2_X1   g357(.A(KEYINPUT91), .B(G104), .Z(new_n544));
  XOR2_X1   g358(.A(new_n543), .B(new_n544), .Z(new_n545));
  AND3_X1   g359(.A1(new_n267), .A2(G143), .A3(G214), .ZN(new_n546));
  AOI21_X1  g360(.A(G143), .B1(new_n267), .B2(G214), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n213), .ZN(new_n549));
  OAI21_X1  g363(.A(G131), .B1(new_n546), .B2(new_n547), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n361), .A2(new_n362), .ZN(new_n552));
  MUX2_X1   g366(.A(new_n380), .B(new_n552), .S(KEYINPUT19), .Z(new_n553));
  OAI211_X1 g367(.A(new_n551), .B(new_n364), .C1(new_n553), .C2(G146), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n356), .A2(G146), .A3(new_n358), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n381), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(KEYINPUT90), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT90), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n381), .A2(new_n558), .A3(new_n555), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT18), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n548), .B1(new_n561), .B2(new_n213), .ZN(new_n562));
  OAI211_X1 g376(.A(KEYINPUT18), .B(G131), .C1(new_n546), .C2(new_n547), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n560), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n545), .B1(new_n554), .B2(new_n564), .ZN(new_n565));
  AND3_X1   g379(.A1(new_n560), .A2(new_n562), .A3(new_n563), .ZN(new_n566));
  OAI211_X1 g380(.A(KEYINPUT17), .B(G131), .C1(new_n546), .C2(new_n547), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n360), .A2(new_n364), .A3(KEYINPUT92), .A4(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT17), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n549), .A2(new_n569), .A3(new_n550), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n360), .A2(new_n364), .A3(new_n567), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT92), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n566), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n565), .B1(new_n575), .B2(new_n545), .ZN(new_n576));
  NOR2_X1   g390(.A1(G475), .A2(G902), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  OAI211_X1 g392(.A(KEYINPUT93), .B(new_n542), .C1(new_n576), .C2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n574), .A2(new_n570), .A3(new_n568), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n580), .A2(new_n564), .A3(new_n545), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n545), .B1(new_n580), .B2(new_n564), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n302), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(G475), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n580), .A2(new_n564), .A3(new_n545), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n554), .A2(new_n564), .ZN(new_n586));
  INV_X1    g400(.A(new_n545), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n578), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT93), .ZN(new_n590));
  OAI21_X1  g404(.A(KEYINPUT20), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AOI211_X1 g405(.A(KEYINPUT93), .B(new_n578), .C1(new_n585), .C2(new_n588), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n579), .B(new_n584), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(G952), .ZN(new_n594));
  AOI211_X1 g408(.A(G953), .B(new_n594), .C1(G234), .C2(G237), .ZN(new_n595));
  AOI211_X1 g409(.A(new_n302), .B(new_n386), .C1(G234), .C2(G237), .ZN(new_n596));
  XNOR2_X1  g410(.A(KEYINPUT21), .B(G898), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n224), .A2(G122), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n224), .A2(G122), .ZN(new_n601));
  OR3_X1    g415(.A1(new_n600), .A2(new_n601), .A3(G107), .ZN(new_n602));
  OAI21_X1  g416(.A(G107), .B1(new_n600), .B2(new_n601), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(G128), .B(G143), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n204), .ZN(new_n606));
  OR2_X1    g420(.A1(new_n606), .A2(KEYINPUT94), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n605), .A2(KEYINPUT13), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n194), .A2(G128), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n608), .B(G134), .C1(KEYINPUT13), .C2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n606), .A2(KEYINPUT94), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n604), .A2(new_n607), .A3(new_n610), .A4(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n599), .A2(KEYINPUT14), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n599), .B1(new_n601), .B2(KEYINPUT14), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n613), .B1(new_n614), .B2(KEYINPUT95), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n615), .B1(KEYINPUT95), .B2(new_n614), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n616), .A2(G107), .ZN(new_n617));
  INV_X1    g431(.A(new_n606), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n605), .A2(new_n204), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n602), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n612), .B1(new_n617), .B2(new_n620), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n403), .A2(new_n346), .A3(G953), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n612), .B(new_n622), .C1(new_n617), .C2(new_n620), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n302), .ZN(new_n627));
  INV_X1    g441(.A(G478), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT96), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n629), .A2(KEYINPUT15), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(KEYINPUT15), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n628), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n627), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n633), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n626), .A2(new_n302), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n593), .A2(new_n598), .A3(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n345), .A2(new_n471), .A3(new_n541), .A4(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G101), .ZN(G3));
  OAI21_X1  g454(.A(new_n302), .B1(new_n331), .B2(new_n332), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n344), .B1(new_n641), .B2(G472), .ZN(new_n642));
  AOI21_X1  g456(.A(KEYINPUT97), .B1(new_n642), .B2(new_n471), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n313), .B1(new_n331), .B2(new_n332), .ZN(new_n644));
  AOI21_X1  g458(.A(G902), .B1(new_n339), .B2(new_n343), .ZN(new_n645));
  INV_X1    g459(.A(G472), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n402), .A2(new_n466), .A3(new_n470), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT97), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n598), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT99), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n620), .B1(new_n616), .B2(G107), .ZN(new_n653));
  AND4_X1   g467(.A1(new_n604), .A2(new_n607), .A3(new_n610), .A4(new_n611), .ZN(new_n654));
  OAI211_X1 g468(.A(KEYINPUT98), .B(new_n623), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n655), .A2(new_n625), .A3(KEYINPUT33), .ZN(new_n656));
  AOI21_X1  g470(.A(KEYINPUT98), .B1(new_n621), .B2(new_n623), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n652), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT33), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n626), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT98), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n653), .A2(new_n654), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n661), .B1(new_n662), .B2(new_n622), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n659), .B1(new_n662), .B2(new_n622), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n663), .A2(new_n664), .A3(KEYINPUT99), .A4(new_n655), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n628), .A2(G902), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n658), .A2(new_n660), .A3(new_n665), .A4(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n627), .A2(new_n628), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n593), .A2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n541), .A2(new_n651), .A3(new_n671), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n643), .A2(new_n650), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(KEYINPUT34), .B(G104), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G6));
  AND2_X1   g489(.A1(new_n634), .A2(new_n636), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n593), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n541), .A2(new_n651), .A3(new_n677), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n643), .A2(new_n650), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT35), .B(G107), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G9));
  NAND2_X1  g495(.A1(new_n454), .A2(new_n456), .ZN(new_n682));
  INV_X1    g496(.A(new_n447), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n445), .A2(KEYINPUT12), .A3(new_n263), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n461), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n682), .B(G469), .C1(new_n685), .C2(new_n453), .ZN(new_n686));
  INV_X1    g500(.A(new_n407), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AOI211_X1 g502(.A(G469), .B(G902), .C1(new_n462), .C2(new_n463), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n404), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n384), .B(KEYINPUT100), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n389), .A2(KEYINPUT36), .ZN(new_n692));
  XOR2_X1   g506(.A(new_n691), .B(new_n692), .Z(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n469), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n690), .B1(new_n402), .B2(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n642), .A2(new_n695), .A3(new_n541), .A4(new_n638), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT37), .B(G110), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G12));
  INV_X1    g512(.A(G900), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n595), .B1(new_n596), .B2(new_n699), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n593), .A2(new_n676), .A3(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n345), .A2(new_n695), .A3(new_n541), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G128), .ZN(G30));
  XNOR2_X1  g517(.A(KEYINPUT102), .B(KEYINPUT39), .ZN(new_n704));
  XOR2_X1   g518(.A(new_n700), .B(new_n704), .Z(new_n705));
  NOR2_X1   g519(.A1(new_n690), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT40), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n530), .A2(new_n540), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(KEYINPUT38), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n402), .A2(new_n694), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n593), .A2(new_n637), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n710), .A2(new_n473), .A3(new_n711), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n266), .A2(new_n299), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n302), .B1(new_n304), .B2(new_n271), .ZN(new_n714));
  OAI21_X1  g528(.A(G472), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  XOR2_X1   g529(.A(new_n715), .B(KEYINPUT101), .Z(new_n716));
  NAND2_X1  g530(.A1(new_n644), .A2(new_n315), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n717), .A3(new_n333), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n707), .A2(new_n709), .A3(new_n712), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G143), .ZN(G45));
  INV_X1    g534(.A(new_n700), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n593), .A2(new_n669), .A3(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n722), .A2(new_n708), .A3(new_n472), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT103), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n541), .A2(KEYINPUT103), .A3(new_n722), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n725), .A2(new_n345), .A3(new_n695), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G146), .ZN(G48));
  AOI21_X1  g542(.A(new_n406), .B1(new_n464), .B2(new_n302), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n729), .A2(new_n689), .A3(new_n405), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n730), .A2(new_n402), .A3(new_n470), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n345), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n732), .A2(new_n672), .ZN(new_n733));
  XOR2_X1   g547(.A(KEYINPUT41), .B(G113), .Z(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(G15));
  INV_X1    g549(.A(new_n678), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT104), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n736), .A2(new_n737), .A3(new_n345), .A4(new_n731), .ZN(new_n738));
  OAI21_X1  g552(.A(KEYINPUT104), .B1(new_n732), .B2(new_n678), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G116), .ZN(G18));
  NAND2_X1  g555(.A1(new_n683), .A2(new_n684), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n456), .A2(new_n441), .ZN(new_n743));
  AOI22_X1  g557(.A1(new_n742), .A2(new_n454), .B1(new_n743), .B2(new_n452), .ZN(new_n744));
  OAI21_X1  g558(.A(G469), .B1(new_n744), .B2(G902), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(new_n404), .A3(new_n465), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n746), .B1(new_n402), .B2(new_n694), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n345), .A2(new_n541), .A3(new_n638), .A4(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G119), .ZN(G21));
  NAND2_X1  g563(.A1(new_n641), .A2(G472), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n393), .A2(new_n394), .A3(new_n396), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT80), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(new_n398), .A3(new_n397), .ZN(new_n754));
  AOI22_X1  g568(.A1(new_n754), .A2(new_n347), .B1(new_n468), .B2(new_n469), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n746), .A2(new_n598), .ZN(new_n756));
  OR2_X1    g570(.A1(new_n305), .A2(new_n307), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n271), .B1(new_n757), .B2(new_n309), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n322), .B1(new_n336), .B2(new_n324), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n313), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n750), .A2(new_n755), .A3(new_n756), .A4(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n541), .A2(new_n637), .A3(new_n593), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XOR2_X1   g577(.A(new_n763), .B(G122), .Z(G24));
  NAND3_X1  g578(.A1(new_n541), .A2(new_n722), .A3(new_n730), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n750), .A2(new_n710), .A3(new_n760), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(new_n355), .ZN(G27));
  AND3_X1   g582(.A1(new_n530), .A2(new_n472), .A3(new_n540), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n345), .A2(new_n471), .A3(new_n769), .A4(new_n722), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT42), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n333), .A2(KEYINPUT105), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT105), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n774), .B(new_n316), .C1(new_n331), .C2(new_n332), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n717), .A2(new_n773), .A3(new_n775), .A4(new_n312), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n530), .A2(new_n472), .A3(new_n540), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n593), .A2(new_n669), .A3(new_n721), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n777), .A2(new_n690), .A3(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n776), .A2(new_n779), .A3(KEYINPUT42), .A4(new_n755), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n772), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G131), .ZN(G33));
  AND2_X1   g596(.A1(new_n312), .A2(new_n333), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n648), .B1(new_n783), .B2(new_n717), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n784), .A2(KEYINPUT106), .A3(new_n701), .A4(new_n769), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n345), .A2(new_n471), .A3(new_n769), .A4(new_n701), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT106), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G134), .ZN(G36));
  OAI21_X1  g604(.A(new_n682), .B1(new_n685), .B2(new_n453), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT45), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n406), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n457), .A2(KEYINPUT45), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n687), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT46), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n689), .B1(new_n796), .B2(new_n797), .ZN(new_n800));
  AOI211_X1 g614(.A(new_n405), .B(new_n705), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n669), .ZN(new_n802));
  OAI21_X1  g616(.A(KEYINPUT43), .B1(new_n802), .B2(new_n593), .ZN(new_n803));
  INV_X1    g617(.A(new_n593), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT43), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n804), .A2(new_n805), .A3(new_n669), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n402), .A2(new_n694), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n807), .A2(new_n642), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n801), .B1(KEYINPUT44), .B2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n807), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n811), .A2(KEYINPUT44), .A3(new_n647), .A4(new_n710), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT107), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n809), .A2(KEYINPUT107), .A3(KEYINPUT44), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n814), .A2(new_n815), .A3(new_n769), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT108), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT44), .ZN(new_n818));
  NOR4_X1   g632(.A1(new_n807), .A2(new_n642), .A3(new_n808), .A4(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n777), .B1(new_n819), .B2(KEYINPUT107), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT108), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n820), .A2(new_n821), .A3(new_n814), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n810), .B1(new_n817), .B2(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(new_n202), .ZN(G39));
  INV_X1    g638(.A(new_n800), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n404), .B1(new_n825), .B2(new_n798), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT47), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g642(.A(KEYINPUT47), .B(new_n404), .C1(new_n825), .C2(new_n798), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n345), .ZN(new_n831));
  INV_X1    g645(.A(new_n755), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n831), .A2(new_n832), .A3(new_n722), .A4(new_n769), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(new_n349), .ZN(G42));
  NOR2_X1   g649(.A1(new_n729), .A2(new_n689), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n837), .A2(KEYINPUT49), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(KEYINPUT49), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n802), .A2(new_n593), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n405), .A2(new_n473), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n838), .A2(new_n839), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  OR4_X1    g656(.A1(new_n832), .A2(new_n842), .A3(new_n709), .A4(new_n718), .ZN(new_n843));
  INV_X1    g657(.A(new_n643), .ZN(new_n844));
  INV_X1    g658(.A(new_n650), .ZN(new_n845));
  OAI21_X1  g659(.A(KEYINPUT109), .B1(new_n593), .B2(new_n676), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n589), .A2(new_n590), .ZN(new_n847));
  AOI22_X1  g661(.A1(new_n847), .A2(new_n542), .B1(new_n583), .B2(G475), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT93), .B1(new_n576), .B2(new_n578), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n589), .A2(new_n590), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n849), .A2(KEYINPUT20), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT109), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n848), .A2(new_n851), .A3(new_n852), .A4(new_n637), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n846), .A2(new_n670), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n854), .A2(new_n541), .A3(new_n651), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n844), .A2(new_n845), .A3(new_n856), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n639), .A2(new_n748), .A3(new_n696), .ZN(new_n858));
  OAI22_X1  g672(.A1(new_n732), .A2(new_n672), .B1(new_n761), .B2(new_n762), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  AND4_X1   g674(.A1(new_n740), .A2(new_n857), .A3(new_n858), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n345), .A2(new_n695), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n593), .A2(new_n637), .A3(new_n700), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n769), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n769), .A2(new_n466), .A3(new_n722), .ZN(new_n865));
  OAI22_X1  g679(.A1(new_n862), .A2(new_n864), .B1(new_n865), .B2(new_n766), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n789), .A2(new_n781), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n702), .B1(new_n766), .B2(new_n765), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT52), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n690), .A2(new_n700), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n712), .A2(new_n718), .A3(new_n708), .A4(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n870), .A2(new_n871), .A3(new_n727), .A4(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n727), .A2(new_n873), .ZN(new_n875));
  OAI21_X1  g689(.A(KEYINPUT52), .B1(new_n875), .B2(new_n869), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n861), .A2(new_n868), .A3(new_n874), .A4(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT53), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(KEYINPUT112), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT54), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n740), .A2(new_n857), .A3(new_n860), .A4(new_n858), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n789), .A2(new_n781), .A3(new_n867), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT110), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n869), .A2(new_n885), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n702), .B(KEYINPUT110), .C1(new_n766), .C2(new_n765), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n886), .A2(new_n727), .A3(new_n873), .A4(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT52), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n884), .A2(new_n889), .A3(KEYINPUT53), .A4(new_n874), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT112), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n643), .A2(new_n650), .A3(new_n855), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n639), .A2(new_n748), .A3(new_n696), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n892), .A2(new_n893), .A3(new_n859), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n866), .B1(new_n772), .B2(new_n780), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n894), .A2(new_n740), .A3(new_n789), .A4(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n876), .A2(new_n874), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n891), .B(new_n878), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n880), .A2(new_n881), .A3(new_n890), .A4(new_n898), .ZN(new_n899));
  OR3_X1    g713(.A1(new_n877), .A2(KEYINPUT111), .A3(new_n878), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n884), .A2(new_n889), .A3(new_n874), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n901), .A2(new_n878), .ZN(new_n902));
  OAI21_X1  g716(.A(KEYINPUT111), .B1(new_n877), .B2(new_n878), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n900), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n899), .B1(new_n904), .B2(new_n881), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n760), .B1(new_n645), .B2(new_n646), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n906), .A2(new_n832), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n803), .A2(new_n595), .A3(new_n806), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n910), .A2(new_n541), .A3(new_n730), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT117), .Z(new_n912));
  AND2_X1   g726(.A1(new_n776), .A2(new_n755), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n777), .A2(new_n746), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n913), .A2(new_n908), .A3(new_n914), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT48), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n755), .A2(new_n595), .ZN(new_n917));
  NOR4_X1   g731(.A1(new_n718), .A2(new_n917), .A3(new_n746), .A4(new_n777), .ZN(new_n918));
  AOI211_X1 g732(.A(new_n594), .B(G953), .C1(new_n918), .C2(new_n671), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n912), .A2(new_n916), .A3(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n918), .A2(new_n804), .A3(new_n802), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n908), .A2(new_n914), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n921), .B1(new_n766), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n836), .A2(new_n405), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n830), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n909), .A2(new_n777), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(KEYINPUT113), .A2(KEYINPUT50), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n910), .A2(new_n730), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n473), .B1(KEYINPUT113), .B2(KEYINPUT50), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n709), .A2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n929), .B1(new_n930), .B2(new_n933), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n930), .A2(new_n929), .A3(new_n933), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n927), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT51), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n937), .A2(KEYINPUT114), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT114), .B1(new_n937), .B2(new_n938), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n920), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n923), .A2(new_n938), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n942), .A2(new_n936), .A3(new_n934), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT115), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n925), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n830), .A2(KEYINPUT115), .A3(new_n924), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n945), .A2(new_n926), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n943), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT116), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n905), .A2(new_n941), .A3(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(G952), .A2(G953), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n843), .B1(new_n950), .B2(new_n951), .ZN(G75));
  NAND2_X1  g766(.A1(new_n898), .A2(new_n890), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n891), .B1(new_n877), .B2(new_n878), .ZN(new_n954));
  OAI211_X1 g768(.A(G210), .B(G902), .C1(new_n953), .C2(new_n954), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n539), .B(new_n481), .ZN(new_n956));
  XNOR2_X1  g770(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n958), .A2(KEYINPUT56), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n955), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n386), .A2(G952), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(KEYINPUT56), .B1(new_n955), .B2(KEYINPUT119), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n964), .B1(KEYINPUT119), .B2(new_n955), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n963), .B1(new_n965), .B2(new_n958), .ZN(G51));
  OAI21_X1  g780(.A(KEYINPUT54), .B1(new_n953), .B2(new_n954), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n899), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n407), .B(KEYINPUT57), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n464), .ZN(new_n971));
  INV_X1    g785(.A(new_n795), .ZN(new_n972));
  OAI211_X1 g786(.A(G902), .B(new_n972), .C1(new_n953), .C2(new_n954), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT120), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n961), .B1(new_n971), .B2(new_n974), .ZN(G54));
  OAI21_X1  g789(.A(G902), .B1(new_n953), .B2(new_n954), .ZN(new_n976));
  NAND2_X1  g790(.A1(KEYINPUT58), .A2(G475), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n576), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n962), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n976), .A2(new_n576), .A3(new_n977), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n979), .A2(new_n980), .ZN(G60));
  AND3_X1   g795(.A1(new_n658), .A2(new_n660), .A3(new_n665), .ZN(new_n982));
  NAND2_X1  g796(.A1(G478), .A2(G902), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT59), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n982), .B1(new_n905), .B2(new_n984), .ZN(new_n985));
  AND3_X1   g799(.A1(new_n968), .A2(new_n982), .A3(new_n984), .ZN(new_n986));
  NOR3_X1   g800(.A1(new_n985), .A2(new_n986), .A3(new_n961), .ZN(G63));
  NAND2_X1  g801(.A1(G217), .A2(G902), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT60), .Z(new_n989));
  OAI21_X1  g803(.A(new_n989), .B1(new_n953), .B2(new_n954), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n467), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n693), .B(new_n989), .C1(new_n953), .C2(new_n954), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n991), .A2(new_n962), .A3(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT61), .ZN(new_n994));
  OR2_X1    g808(.A1(new_n994), .A2(KEYINPUT121), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(KEYINPUT121), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n993), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n961), .B1(new_n990), .B2(new_n467), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n998), .A2(KEYINPUT121), .A3(new_n994), .A4(new_n992), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n997), .A2(new_n999), .ZN(G66));
  INV_X1    g814(.A(new_n597), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n386), .B1(new_n1001), .B2(G224), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1002), .B1(new_n882), .B2(new_n386), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n539), .B1(G898), .B2(new_n386), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1004), .B(KEYINPUT122), .Z(new_n1005));
  XNOR2_X1  g819(.A(new_n1003), .B(new_n1005), .ZN(G69));
  AOI21_X1  g820(.A(new_n386), .B1(G227), .B2(G900), .ZN(new_n1007));
  INV_X1    g821(.A(new_n705), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n784), .A2(new_n1008), .A3(new_n769), .A4(new_n854), .ZN(new_n1009));
  INV_X1    g823(.A(new_n1009), .ZN(new_n1010));
  NOR3_X1   g824(.A1(new_n823), .A2(new_n834), .A3(new_n1010), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n886), .A2(new_n719), .A3(new_n727), .A4(new_n887), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1012), .B(KEYINPUT62), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(KEYINPUT124), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g829(.A(new_n810), .ZN(new_n1016));
  AND4_X1   g830(.A1(new_n821), .A2(new_n814), .A3(new_n769), .A4(new_n815), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n821), .B1(new_n820), .B2(new_n814), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1016), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(new_n834), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n1019), .A2(new_n1020), .A3(new_n1009), .ZN(new_n1021));
  INV_X1    g835(.A(KEYINPUT124), .ZN(new_n1022));
  NOR3_X1   g836(.A1(new_n1021), .A2(new_n1022), .A3(new_n1013), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n386), .B1(new_n1015), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n260), .A2(new_n320), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n1025), .B(new_n553), .ZN(new_n1026));
  XNOR2_X1  g840(.A(new_n1026), .B(KEYINPUT123), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n823), .A2(new_n834), .ZN(new_n1029));
  INV_X1    g843(.A(new_n762), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n801), .A2(new_n1030), .A3(new_n913), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1031), .A2(new_n781), .A3(new_n789), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n886), .A2(new_n727), .A3(new_n887), .ZN(new_n1033));
  NOR2_X1   g847(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g848(.A(G953), .B1(new_n1029), .B2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g849(.A1(new_n386), .A2(G900), .ZN(new_n1036));
  XNOR2_X1  g850(.A(new_n1036), .B(KEYINPUT125), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n1026), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n1007), .B1(new_n1028), .B2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g853(.A1(new_n1011), .A2(KEYINPUT124), .A3(new_n1014), .ZN(new_n1040));
  OAI21_X1  g854(.A(new_n1022), .B1(new_n1021), .B2(new_n1013), .ZN(new_n1041));
  AOI21_X1  g855(.A(G953), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g856(.A(new_n1027), .ZN(new_n1043));
  OAI211_X1 g857(.A(new_n1038), .B(new_n1007), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1044));
  INV_X1    g858(.A(new_n1044), .ZN(new_n1045));
  NOR2_X1   g859(.A1(new_n1039), .A2(new_n1045), .ZN(G72));
  NAND2_X1  g860(.A1(G472), .A2(G902), .ZN(new_n1047));
  XOR2_X1   g861(.A(new_n1047), .B(KEYINPUT63), .Z(new_n1048));
  INV_X1    g862(.A(new_n1048), .ZN(new_n1049));
  NOR2_X1   g863(.A1(new_n266), .A2(new_n271), .ZN(new_n1050));
  INV_X1    g864(.A(new_n1050), .ZN(new_n1051));
  OR2_X1    g865(.A1(new_n1051), .A2(KEYINPUT126), .ZN(new_n1052));
  AOI21_X1  g866(.A(new_n336), .B1(new_n1051), .B2(KEYINPUT126), .ZN(new_n1053));
  AOI21_X1  g867(.A(new_n1049), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OAI211_X1 g868(.A(new_n900), .B(new_n1054), .C1(new_n902), .C2(new_n903), .ZN(new_n1055));
  NAND4_X1  g869(.A1(new_n1019), .A2(new_n1020), .A3(new_n861), .A4(new_n1034), .ZN(new_n1056));
  NAND2_X1  g870(.A1(new_n1056), .A2(new_n1048), .ZN(new_n1057));
  AND2_X1   g871(.A1(new_n266), .A2(new_n299), .ZN(new_n1058));
  AOI21_X1  g872(.A(new_n961), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g873(.A1(new_n1055), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g874(.A(new_n1060), .ZN(new_n1061));
  NAND3_X1  g875(.A1(new_n1040), .A2(new_n1041), .A3(new_n861), .ZN(new_n1062));
  AND2_X1   g876(.A1(new_n1062), .A2(new_n1048), .ZN(new_n1063));
  INV_X1    g877(.A(new_n713), .ZN(new_n1064));
  OAI211_X1 g878(.A(new_n1061), .B(KEYINPUT127), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1065));
  INV_X1    g879(.A(KEYINPUT127), .ZN(new_n1066));
  AOI21_X1  g880(.A(new_n1064), .B1(new_n1062), .B2(new_n1048), .ZN(new_n1067));
  OAI21_X1  g881(.A(new_n1066), .B1(new_n1067), .B2(new_n1060), .ZN(new_n1068));
  NAND2_X1  g882(.A1(new_n1065), .A2(new_n1068), .ZN(G57));
endmodule


