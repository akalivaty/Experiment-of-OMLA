//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 0 1 0 1 0 0 0 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 1 1 0 1 1 1 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n594, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n653, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n840, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G137), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT11), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT64), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT64), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT11), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n189), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G137), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G134), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n188), .A2(G137), .ZN(new_n197));
  AOI22_X1  g011(.A1(new_n196), .A2(new_n197), .B1(KEYINPUT64), .B2(new_n190), .ZN(new_n198));
  OAI21_X1  g012(.A(G131), .B1(new_n194), .B2(new_n198), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n192), .A2(KEYINPUT11), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n190), .A2(KEYINPUT64), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n196), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n195), .A2(G134), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n191), .B1(new_n189), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G131), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n202), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n199), .A2(new_n206), .A3(KEYINPUT65), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT65), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n208), .B(G131), .C1(new_n194), .C2(new_n198), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT70), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G143), .ZN(new_n214));
  INV_X1    g028(.A(G143), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G146), .ZN(new_n216));
  AND2_X1   g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT0), .ZN(new_n218));
  INV_X1    g032(.A(G128), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  XOR2_X1   g034(.A(KEYINPUT0), .B(G128), .Z(new_n221));
  OAI21_X1  g035(.A(new_n220), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n207), .A2(KEYINPUT70), .A3(new_n209), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n212), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT71), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT1), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n217), .A2(new_n227), .A3(G128), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n214), .A2(new_n216), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT66), .B(G128), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n227), .B1(G143), .B2(new_n213), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n228), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(G131), .B1(new_n189), .B2(new_n203), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n233), .A2(new_n206), .A3(new_n234), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n212), .A2(KEYINPUT71), .A3(new_n222), .A4(new_n223), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n226), .A2(KEYINPUT30), .A3(new_n235), .A4(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G116), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G119), .ZN(new_n239));
  XNOR2_X1  g053(.A(new_n239), .B(KEYINPUT69), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT68), .B(G119), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G116), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(KEYINPUT2), .B(G113), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n246), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n241), .A2(new_n248), .A3(new_n244), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  OR2_X1    g064(.A1(new_n235), .A2(KEYINPUT67), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n235), .A2(KEYINPUT67), .ZN(new_n252));
  INV_X1    g066(.A(new_n222), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n251), .B(new_n252), .C1(new_n253), .C2(new_n210), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT30), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n237), .A2(new_n250), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT72), .ZN(new_n258));
  INV_X1    g072(.A(new_n250), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n226), .A2(new_n259), .A3(new_n235), .A4(new_n236), .ZN(new_n260));
  NOR2_X1   g074(.A1(G237), .A2(G953), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G210), .ZN(new_n262));
  INV_X1    g076(.A(G101), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n262), .B(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n265));
  XOR2_X1   g079(.A(new_n264), .B(new_n265), .Z(new_n266));
  INV_X1    g080(.A(KEYINPUT72), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n237), .A2(new_n267), .A3(new_n250), .A4(new_n256), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n258), .A2(new_n260), .A3(new_n266), .A4(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT73), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n268), .A2(new_n260), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT73), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n271), .A2(new_n272), .A3(new_n266), .A4(new_n258), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n270), .A2(new_n273), .A3(KEYINPUT31), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT31), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n269), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT28), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT74), .ZN(new_n279));
  AND3_X1   g093(.A1(new_n254), .A2(new_n279), .A3(new_n250), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n279), .B1(new_n254), .B2(new_n250), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n278), .B1(new_n282), .B2(new_n260), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n259), .A2(new_n235), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT28), .B1(new_n284), .B2(new_n224), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT75), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n285), .B(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n288), .A2(new_n266), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n277), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(G472), .A2(G902), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT76), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n289), .B1(new_n274), .B2(new_n276), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT76), .ZN(new_n295));
  INV_X1    g109(.A(new_n292), .ZN(new_n296));
  NOR3_X1   g110(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n187), .B1(new_n293), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n291), .A2(KEYINPUT32), .A3(new_n292), .ZN(new_n299));
  INV_X1    g113(.A(new_n287), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n266), .A2(KEYINPUT29), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n226), .A2(new_n235), .A3(new_n236), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n250), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n260), .ZN(new_n304));
  AOI21_X1  g118(.A(KEYINPUT77), .B1(new_n304), .B2(KEYINPUT28), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT77), .ZN(new_n306));
  AOI211_X1 g120(.A(new_n306), .B(new_n278), .C1(new_n303), .C2(new_n260), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n300), .B(new_n301), .C1(new_n305), .C2(new_n307), .ZN(new_n308));
  OR2_X1    g122(.A1(new_n308), .A2(KEYINPUT78), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT29), .B1(new_n288), .B2(new_n266), .ZN(new_n310));
  INV_X1    g124(.A(new_n266), .ZN(new_n311));
  INV_X1    g125(.A(new_n258), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n268), .A2(new_n260), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(G902), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n308), .A2(KEYINPUT78), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n309), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G472), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n298), .A2(new_n299), .A3(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G125), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n320), .A2(G140), .ZN(new_n321));
  XNOR2_X1  g135(.A(G125), .B(G140), .ZN(new_n322));
  MUX2_X1   g136(.A(new_n321), .B(new_n322), .S(KEYINPUT16), .Z(new_n323));
  XNOR2_X1  g137(.A(new_n323), .B(G146), .ZN(new_n324));
  AOI22_X1  g138(.A1(new_n243), .A2(G128), .B1(new_n230), .B2(G119), .ZN(new_n325));
  XOR2_X1   g139(.A(KEYINPUT24), .B(G110), .Z(new_n326));
  AOI21_X1  g140(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G110), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT23), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n242), .A2(new_n329), .A3(new_n219), .ZN(new_n330));
  INV_X1    g144(.A(new_n325), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n330), .B1(new_n331), .B2(new_n329), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n327), .B1(new_n328), .B2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n322), .B(KEYINPUT79), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n334), .A2(new_n213), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n323), .A2(new_n213), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n332), .A2(new_n328), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n325), .A2(new_n326), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n333), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT22), .B(G137), .ZN(new_n342));
  INV_X1    g156(.A(G953), .ZN(new_n343));
  AND3_X1   g157(.A1(new_n343), .A2(G221), .A3(G234), .ZN(new_n344));
  XOR2_X1   g158(.A(new_n342), .B(new_n344), .Z(new_n345));
  XNOR2_X1  g159(.A(new_n341), .B(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G902), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  XOR2_X1   g162(.A(new_n348), .B(KEYINPUT25), .Z(new_n349));
  INV_X1    g163(.A(G217), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n350), .B1(G234), .B2(new_n347), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n351), .A2(G902), .ZN(new_n353));
  XOR2_X1   g167(.A(new_n353), .B(KEYINPUT80), .Z(new_n354));
  NAND2_X1  g168(.A1(new_n346), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(G214), .B1(G237), .B2(G902), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(G210), .B1(G237), .B2(G902), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n233), .A2(new_n320), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n361), .B1(new_n253), .B2(new_n320), .ZN(new_n362));
  INV_X1    g176(.A(G224), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n363), .A2(G953), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n362), .B(new_n365), .ZN(new_n366));
  AND3_X1   g180(.A1(new_n241), .A2(KEYINPUT5), .A3(new_n244), .ZN(new_n367));
  OAI21_X1  g181(.A(G113), .B1(new_n244), .B2(KEYINPUT5), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n249), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G104), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G107), .ZN(new_n371));
  INV_X1    g185(.A(G107), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G104), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT3), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(KEYINPUT3), .B1(new_n372), .B2(G104), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n371), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n377), .A2(G101), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n263), .B1(new_n371), .B2(new_n373), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  OR2_X1    g195(.A1(new_n369), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT4), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n378), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n377), .A2(G101), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n377), .A2(new_n383), .A3(G101), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n250), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n382), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT86), .ZN(new_n390));
  XOR2_X1   g204(.A(G110), .B(G122), .Z(new_n391));
  NAND3_X1  g205(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT6), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n391), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n382), .A2(new_n388), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n392), .A2(new_n393), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n366), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  XOR2_X1   g213(.A(new_n391), .B(KEYINPUT8), .Z(new_n400));
  INV_X1    g214(.A(new_n382), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n369), .A2(new_n381), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n366), .B1(KEYINPUT7), .B2(new_n364), .ZN(new_n404));
  OR3_X1    g218(.A1(new_n362), .A2(KEYINPUT7), .A3(new_n364), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n403), .A2(new_n404), .A3(new_n396), .A4(new_n405), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n406), .A2(new_n347), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n360), .B1(new_n399), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n399), .A2(new_n407), .A3(new_n360), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n359), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G221), .ZN(new_n412));
  XOR2_X1   g226(.A(KEYINPUT9), .B(G234), .Z(new_n413));
  AOI21_X1  g227(.A(new_n412), .B1(new_n413), .B2(new_n347), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G469), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n231), .A2(new_n219), .ZN(new_n417));
  OAI21_X1  g231(.A(KEYINPUT83), .B1(new_n417), .B2(new_n217), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n228), .ZN(new_n419));
  NOR3_X1   g233(.A1(new_n417), .A2(new_n217), .A3(KEYINPUT83), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n380), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT10), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT84), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n423), .B(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n212), .A2(new_n223), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n386), .A2(new_n222), .A3(new_n387), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n380), .A2(KEYINPUT10), .A3(new_n233), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n425), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  XOR2_X1   g244(.A(G110), .B(G140), .Z(new_n431));
  INV_X1    g245(.A(G227), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n432), .A2(G953), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n431), .B(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(KEYINPUT81), .B(KEYINPUT82), .ZN(new_n435));
  XOR2_X1   g249(.A(new_n434), .B(new_n435), .Z(new_n436));
  NAND2_X1  g250(.A1(new_n430), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n426), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n421), .B1(new_n233), .B2(new_n380), .ZN(new_n439));
  AOI21_X1  g253(.A(KEYINPUT12), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n207), .A2(KEYINPUT12), .A3(new_n209), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n440), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n437), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n425), .A2(new_n429), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n438), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n436), .B1(new_n445), .B2(new_n430), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n416), .B(new_n347), .C1(new_n443), .C2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(G469), .A2(G902), .ZN(new_n448));
  INV_X1    g262(.A(new_n436), .ZN(new_n449));
  INV_X1    g263(.A(new_n430), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n449), .B1(new_n450), .B2(new_n442), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n437), .A2(KEYINPUT85), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n445), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n437), .A2(KEYINPUT85), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n451), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n447), .B(new_n448), .C1(new_n455), .C2(new_n416), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n411), .A2(new_n415), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n413), .ZN(new_n458));
  NOR3_X1   g272(.A1(new_n458), .A2(new_n350), .A3(G953), .ZN(new_n459));
  INV_X1    g273(.A(G122), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(G116), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(KEYINPUT91), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n238), .A2(G122), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n463), .B(KEYINPUT92), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n372), .B1(new_n462), .B2(KEYINPUT14), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n465), .B(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n230), .A2(G143), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n215), .A2(G128), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(KEYINPUT94), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT94), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n468), .A2(new_n472), .A3(new_n469), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n471), .A2(new_n188), .A3(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n188), .B1(new_n471), .B2(new_n473), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n467), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT95), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT95), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n467), .B(new_n479), .C1(new_n475), .C2(new_n476), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n465), .B(new_n372), .ZN(new_n482));
  AOI22_X1  g296(.A1(new_n468), .A2(KEYINPUT13), .B1(G128), .B2(new_n215), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n215), .A2(KEYINPUT13), .A3(G128), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n484), .B(KEYINPUT93), .ZN(new_n485));
  OAI21_X1  g299(.A(G134), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n482), .A2(new_n474), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n459), .B1(new_n481), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n481), .A2(new_n487), .A3(new_n459), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n347), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(G478), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n492), .A2(KEYINPUT15), .ZN(new_n493));
  OR2_X1    g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n261), .A2(G214), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT87), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n495), .A2(new_n496), .A3(G143), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(G143), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n215), .A2(KEYINPUT87), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n498), .A2(new_n499), .A3(G214), .A4(new_n261), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n501), .B(G131), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n502), .A2(new_n336), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT19), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n334), .A2(new_n504), .ZN(new_n505));
  XOR2_X1   g319(.A(new_n505), .B(KEYINPUT89), .Z(new_n506));
  NOR2_X1   g320(.A1(new_n322), .A2(new_n504), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n507), .B(KEYINPUT88), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n503), .B1(new_n509), .B2(G146), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT18), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n501), .B1(new_n511), .B2(new_n205), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n501), .A2(new_n205), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n322), .A2(new_n213), .ZN(new_n515));
  OAI221_X1 g329(.A(new_n512), .B1(new_n514), .B2(new_n511), .C1(new_n335), .C2(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(G113), .B(G122), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(new_n370), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT17), .ZN(new_n521));
  AND2_X1   g335(.A1(new_n502), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n324), .B1(new_n521), .B2(new_n514), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n516), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g338(.A1(new_n510), .A2(new_n520), .B1(new_n524), .B2(new_n518), .ZN(new_n525));
  NOR2_X1   g339(.A1(G475), .A2(G902), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT20), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT20), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n525), .A2(new_n529), .A3(new_n526), .ZN(new_n530));
  OR2_X1    g344(.A1(new_n518), .A2(KEYINPUT90), .ZN(new_n531));
  AOI21_X1  g345(.A(G902), .B1(new_n524), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n532), .B1(new_n531), .B2(new_n524), .ZN(new_n533));
  AOI22_X1  g347(.A1(new_n528), .A2(new_n530), .B1(G475), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G952), .ZN(new_n535));
  AOI211_X1 g349(.A(G953), .B(new_n535), .C1(G234), .C2(G237), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  AOI211_X1 g351(.A(new_n347), .B(new_n343), .C1(G234), .C2(G237), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  XOR2_X1   g353(.A(KEYINPUT21), .B(G898), .Z(new_n540));
  OAI21_X1  g354(.A(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(KEYINPUT96), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n491), .A2(new_n493), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n494), .A2(new_n534), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n457), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n319), .A2(new_n357), .A3(new_n545), .ZN(new_n546));
  XNOR2_X1  g360(.A(KEYINPUT97), .B(G101), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n546), .B(new_n547), .ZN(G3));
  NAND3_X1  g362(.A1(new_n291), .A2(KEYINPUT76), .A3(new_n292), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n295), .B1(new_n294), .B2(new_n296), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(G472), .B1(new_n294), .B2(G902), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n357), .A2(new_n415), .A3(new_n456), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n411), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT98), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT33), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(KEYINPUT98), .A2(KEYINPUT33), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n560), .B(new_n561), .C1(new_n490), .C2(new_n488), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n481), .A2(new_n487), .ZN(new_n563));
  INV_X1    g377(.A(new_n459), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n565), .A2(new_n558), .A3(new_n559), .A4(new_n489), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n492), .A2(G902), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n567), .A2(new_n568), .B1(new_n491), .B2(new_n492), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n534), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n542), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n557), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n556), .A2(new_n574), .ZN(new_n575));
  XOR2_X1   g389(.A(KEYINPUT34), .B(G104), .Z(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(G6));
  XNOR2_X1  g391(.A(new_n542), .B(KEYINPUT99), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n411), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n494), .A2(new_n543), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n534), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n556), .A2(new_n582), .ZN(new_n583));
  XOR2_X1   g397(.A(KEYINPUT35), .B(G107), .Z(new_n584));
  XNOR2_X1  g398(.A(new_n583), .B(new_n584), .ZN(G9));
  INV_X1    g399(.A(new_n345), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n586), .A2(KEYINPUT36), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n341), .B(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n354), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n352), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n551), .A2(new_n545), .A3(new_n552), .A4(new_n590), .ZN(new_n591));
  XOR2_X1   g405(.A(KEYINPUT37), .B(G110), .Z(new_n592));
  XNOR2_X1  g406(.A(new_n591), .B(new_n592), .ZN(G12));
  INV_X1    g407(.A(new_n581), .ZN(new_n594));
  INV_X1    g408(.A(G900), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n536), .B1(new_n538), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g412(.A(new_n598), .B(KEYINPUT100), .Z(new_n599));
  INV_X1    g413(.A(new_n457), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n319), .A2(new_n599), .A3(new_n600), .A4(new_n590), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(G128), .ZN(G30));
  NAND2_X1  g416(.A1(new_n270), .A2(new_n273), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n304), .A2(new_n311), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(G472), .B1(new_n605), .B2(G902), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n299), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(KEYINPUT101), .B1(new_n298), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(KEYINPUT32), .B1(new_n549), .B2(new_n550), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n299), .A2(new_n606), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT101), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n590), .ZN(new_n615));
  INV_X1    g429(.A(new_n410), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n616), .A2(new_n408), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(KEYINPUT38), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n580), .A2(new_n571), .ZN(new_n619));
  NOR3_X1   g433(.A1(new_n618), .A2(new_n359), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n456), .A2(new_n415), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n596), .B(KEYINPUT39), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n620), .B1(KEYINPUT40), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n626), .B1(KEYINPUT40), .B2(new_n625), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n614), .A2(new_n615), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT102), .ZN(new_n629));
  XNOR2_X1  g443(.A(KEYINPUT103), .B(G143), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G45));
  NAND2_X1  g445(.A1(new_n299), .A2(new_n318), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n600), .B(new_n590), .C1(new_n609), .C2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n570), .A2(new_n571), .A3(new_n597), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(new_n213), .ZN(G48));
  NOR2_X1   g450(.A1(new_n609), .A2(new_n632), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n637), .A2(new_n356), .ZN(new_n638));
  INV_X1    g452(.A(new_n443), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n445), .A2(new_n430), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n449), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n416), .B1(new_n642), .B2(new_n347), .ZN(new_n643));
  INV_X1    g457(.A(new_n447), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n415), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n638), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n574), .ZN(new_n650));
  XNOR2_X1  g464(.A(KEYINPUT41), .B(G113), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G15));
  NAND2_X1  g466(.A1(new_n649), .A2(new_n582), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G116), .ZN(G18));
  NOR3_X1   g468(.A1(new_n646), .A2(new_n557), .A3(new_n544), .ZN(new_n655));
  OAI211_X1 g469(.A(new_n655), .B(new_n590), .C1(new_n609), .C2(new_n632), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G119), .ZN(G21));
  NAND3_X1  g471(.A1(new_n645), .A2(new_n415), .A3(new_n578), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n411), .A2(new_n580), .A3(new_n571), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n300), .B1(new_n305), .B2(new_n307), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n311), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n277), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n292), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n660), .A2(new_n357), .A3(new_n552), .A4(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G122), .ZN(G24));
  NAND2_X1  g480(.A1(new_n664), .A2(new_n552), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n667), .A2(new_n615), .ZN(new_n668));
  INV_X1    g482(.A(new_n634), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n646), .A2(new_n557), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT104), .B(G125), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G27));
  OAI21_X1  g487(.A(new_n187), .B1(new_n294), .B2(new_n296), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n299), .A2(new_n318), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n617), .A2(new_n358), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n621), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n675), .A2(new_n357), .A3(new_n669), .A4(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(KEYINPUT42), .ZN(new_n679));
  OAI211_X1 g493(.A(new_n357), .B(new_n677), .C1(new_n609), .C2(new_n632), .ZN(new_n680));
  OR2_X1    g494(.A1(new_n634), .A2(KEYINPUT42), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n679), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(new_n205), .ZN(G33));
  XNOR2_X1  g497(.A(new_n598), .B(KEYINPUT100), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(new_n188), .ZN(G36));
  XNOR2_X1  g500(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n687), .B1(new_n569), .B2(new_n571), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT107), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n569), .A2(new_n571), .ZN(new_n690));
  AOI22_X1  g504(.A1(new_n688), .A2(new_n689), .B1(new_n690), .B2(KEYINPUT43), .ZN(new_n691));
  OR2_X1    g505(.A1(new_n688), .A2(new_n689), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n590), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n553), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n676), .B1(new_n695), .B2(KEYINPUT44), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n697));
  OR2_X1    g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n696), .A2(new_n697), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n695), .A2(KEYINPUT44), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT45), .ZN(new_n701));
  OR2_X1    g515(.A1(new_n455), .A2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n416), .B1(new_n455), .B2(new_n701), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n703), .B1(new_n702), .B2(new_n704), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n448), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT46), .ZN(new_n708));
  AND2_X1   g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n447), .B1(new_n707), .B2(new_n708), .ZN(new_n710));
  OR2_X1    g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n711), .A2(new_n415), .A3(new_n624), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n698), .A2(new_n699), .A3(new_n700), .A4(new_n713), .ZN(new_n714));
  XOR2_X1   g528(.A(KEYINPUT109), .B(G137), .Z(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G39));
  INV_X1    g530(.A(KEYINPUT47), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n711), .A2(new_n717), .A3(new_n415), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n357), .A2(new_n676), .A3(new_n634), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n637), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(KEYINPUT110), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n717), .B1(new_n711), .B2(new_n415), .ZN(new_n723));
  OR3_X1    g537(.A1(new_n719), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G140), .ZN(G42));
  NAND4_X1  g539(.A1(new_n357), .A2(new_n358), .A3(new_n415), .A4(new_n690), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(KEYINPUT111), .ZN(new_n727));
  OAI21_X1  g541(.A(KEYINPUT49), .B1(new_n643), .B2(new_n644), .ZN(new_n728));
  OR3_X1    g542(.A1(new_n643), .A2(KEYINPUT49), .A3(new_n644), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n618), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n613), .A2(new_n727), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n537), .B1(new_n691), .B2(new_n692), .ZN(new_n732));
  AND4_X1   g546(.A1(new_n358), .A2(new_n732), .A3(new_n617), .A4(new_n647), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n675), .A2(new_n357), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g549(.A(KEYINPUT48), .B1(new_n735), .B2(KEYINPUT119), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(KEYINPUT119), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n667), .A2(new_n356), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n732), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n740), .A2(new_n557), .A3(new_n646), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n741), .A2(new_n535), .A3(G953), .ZN(new_n742));
  NOR4_X1   g556(.A1(new_n646), .A2(new_n356), .A3(new_n676), .A4(new_n537), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n613), .A2(new_n743), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n738), .B(new_n742), .C1(new_n572), .C2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n645), .A2(new_n414), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n746), .B1(new_n719), .B2(new_n723), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n740), .A2(new_n676), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n618), .A2(new_n359), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n739), .A2(new_n647), .A3(new_n750), .A4(new_n732), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(KEYINPUT117), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(KEYINPUT118), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT50), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT118), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n754), .B1(new_n751), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n752), .A2(KEYINPUT118), .A3(new_n754), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n733), .A2(new_n668), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n613), .A2(new_n534), .A3(new_n569), .A4(new_n743), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n757), .A2(new_n758), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n749), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT116), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n764), .B1(new_n761), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n749), .A2(new_n762), .A3(new_n765), .A4(new_n764), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n745), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n319), .A2(new_n600), .A3(new_n590), .A4(new_n669), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n601), .A2(new_n770), .A3(new_n671), .ZN(new_n771));
  INV_X1    g585(.A(new_n659), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(new_n622), .A3(new_n597), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n611), .B1(new_n609), .B2(new_n610), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n298), .A2(new_n607), .A3(KEYINPUT101), .ZN(new_n775));
  AOI211_X1 g589(.A(new_n590), .B(new_n773), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n771), .A2(new_n776), .A3(KEYINPUT52), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n671), .B1(new_n633), .B2(new_n684), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(new_n635), .ZN(new_n780));
  INV_X1    g594(.A(new_n773), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n615), .B(new_n781), .C1(new_n608), .C2(new_n612), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n778), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(KEYINPUT115), .B1(new_n777), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(KEYINPUT52), .B1(new_n771), .B2(new_n776), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n780), .A2(new_n778), .A3(new_n782), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n682), .A2(new_n685), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n591), .A2(new_n665), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n594), .B1(new_n572), .B2(KEYINPUT112), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n572), .A2(KEYINPUT112), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n579), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n553), .A2(new_n554), .A3(new_n793), .ZN(new_n794));
  AND4_X1   g608(.A1(new_n546), .A2(new_n790), .A3(new_n656), .A4(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT114), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n494), .A2(new_n534), .A3(new_n543), .A4(new_n597), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT113), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n677), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n319), .A2(new_n796), .A3(new_n590), .A4(new_n799), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n799), .B(new_n590), .C1(new_n609), .C2(new_n632), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT114), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n667), .A2(new_n615), .A3(new_n634), .ZN(new_n803));
  AOI22_X1  g617(.A1(new_n800), .A2(new_n802), .B1(new_n803), .B2(new_n677), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n638), .B(new_n647), .C1(new_n574), .C2(new_n582), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n789), .A2(new_n795), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n784), .A2(KEYINPUT53), .A3(new_n788), .A4(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n785), .A2(new_n786), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n810), .B1(new_n811), .B2(new_n806), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n808), .A2(new_n809), .A3(new_n812), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n811), .A2(new_n806), .A3(new_n810), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n784), .A2(new_n788), .A3(new_n807), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n814), .B1(new_n815), .B2(new_n810), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n769), .B(new_n813), .C1(new_n809), .C2(new_n816), .ZN(new_n817));
  OAI22_X1  g631(.A1(new_n817), .A2(KEYINPUT120), .B1(G952), .B2(G953), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n817), .A2(KEYINPUT120), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n731), .B1(new_n818), .B2(new_n819), .ZN(G75));
  AOI21_X1  g634(.A(new_n347), .B1(new_n808), .B2(new_n812), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT56), .B1(new_n821), .B2(G210), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n397), .A2(new_n398), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(new_n366), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(KEYINPUT55), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n822), .A2(new_n825), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n343), .A2(G952), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(G51));
  XNOR2_X1  g643(.A(new_n642), .B(KEYINPUT121), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n808), .A2(new_n812), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(KEYINPUT54), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(new_n813), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n448), .B(KEYINPUT57), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n830), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n821), .ZN(new_n837));
  OR3_X1    g651(.A1(new_n837), .A2(new_n705), .A3(new_n706), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n828), .B1(new_n836), .B2(new_n838), .ZN(G54));
  AND2_X1   g653(.A1(KEYINPUT58), .A2(G475), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n821), .A2(new_n525), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n525), .B1(new_n821), .B2(new_n840), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n841), .A2(new_n842), .A3(new_n828), .ZN(G60));
  OAI21_X1  g657(.A(new_n813), .B1(new_n816), .B2(new_n809), .ZN(new_n844));
  NAND2_X1  g658(.A1(G478), .A2(G902), .ZN(new_n845));
  XOR2_X1   g659(.A(new_n845), .B(KEYINPUT59), .Z(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n567), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT122), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n849), .A2(new_n846), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n828), .B1(new_n833), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n850), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n808), .A2(new_n809), .A3(new_n812), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n809), .B1(new_n808), .B2(new_n812), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n852), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n828), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n567), .B1(new_n844), .B2(new_n847), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT122), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n854), .A2(new_n861), .ZN(G63));
  NAND2_X1  g676(.A1(G217), .A2(G902), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(KEYINPUT60), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n864), .B1(new_n808), .B2(new_n812), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n828), .B1(new_n865), .B2(new_n588), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n866), .B1(new_n346), .B2(new_n865), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT61), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n867), .B(new_n868), .ZN(G66));
  INV_X1    g683(.A(new_n540), .ZN(new_n870));
  OAI21_X1  g684(.A(G953), .B1(new_n870), .B2(new_n363), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n795), .A2(new_n805), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n871), .B1(new_n873), .B2(G953), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n823), .B1(G898), .B2(new_n343), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n874), .B(new_n875), .ZN(G69));
  NAND2_X1  g690(.A1(new_n791), .A2(new_n792), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT124), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n624), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n879), .B1(new_n878), .B2(new_n877), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n880), .A2(new_n638), .A3(new_n677), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n882), .A2(KEYINPUT125), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(KEYINPUT125), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n724), .A2(new_n714), .A3(new_n883), .A4(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT62), .ZN(new_n886));
  OR3_X1    g700(.A1(new_n629), .A2(new_n886), .A3(new_n771), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n886), .B1(new_n629), .B2(new_n771), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n885), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n509), .B(KEYINPUT123), .Z(new_n890));
  NAND2_X1  g704(.A1(new_n237), .A2(new_n256), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n890), .B(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n343), .B1(new_n892), .B2(G900), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n713), .A2(new_n772), .A3(new_n734), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n771), .A2(new_n682), .A3(new_n685), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n724), .A2(new_n714), .A3(new_n896), .A4(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n893), .A2(G953), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n895), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n894), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n343), .B1(G227), .B2(G900), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT126), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n901), .B(new_n903), .ZN(G72));
  XNOR2_X1  g718(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n905));
  NAND2_X1  g719(.A1(G472), .A2(G902), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n905), .B(new_n906), .Z(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n908), .B1(new_n898), .B2(new_n872), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n312), .A2(new_n313), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n911), .A2(new_n266), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n828), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n907), .B1(new_n889), .B2(new_n873), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n911), .A2(new_n266), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AOI211_X1 g730(.A(new_n907), .B(new_n816), .C1(new_n603), .C2(new_n314), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n916), .A2(new_n917), .ZN(G57));
endmodule


