//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 1 1 0 1 0 0 0 0 1 1 0 0 1 0 1 0 1 1 1 1 0 1 0 0 0 0 1 0 1 1 0 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955;
  XNOR2_X1  g000(.A(KEYINPUT69), .B(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(G143), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G146), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT0), .A2(G128), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  NOR2_X1   g007(.A1(KEYINPUT0), .A2(G128), .ZN(new_n194));
  OAI22_X1  g008(.A1(new_n189), .A2(new_n191), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(G143), .B(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(new_n192), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT66), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT11), .ZN(new_n200));
  INV_X1    g014(.A(G134), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(G137), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(G137), .ZN(new_n203));
  INV_X1    g017(.A(G137), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT11), .A3(G134), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n202), .A2(new_n203), .A3(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G131), .ZN(new_n207));
  INV_X1    g021(.A(G131), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n202), .A2(new_n205), .A3(new_n208), .A4(new_n203), .ZN(new_n209));
  AND2_X1   g023(.A1(new_n209), .A2(KEYINPUT64), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n209), .A2(KEYINPUT64), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n199), .B(new_n207), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(new_n209), .B(KEYINPUT64), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n199), .B1(new_n214), .B2(new_n207), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n198), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n203), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n201), .A2(G137), .ZN(new_n218));
  OAI21_X1  g032(.A(G131), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G128), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n196), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n189), .A2(new_n220), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n191), .B1(KEYINPUT1), .B2(new_n220), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n214), .A2(new_n219), .A3(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n216), .A2(KEYINPUT30), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G119), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G116), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT65), .B(G116), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n229), .B1(new_n230), .B2(new_n228), .ZN(new_n231));
  XOR2_X1   g045(.A(KEYINPUT2), .B(G113), .Z(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n232), .B(new_n229), .C1(new_n228), .C2(new_n230), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n207), .B1(new_n210), .B2(new_n211), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(new_n198), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(new_n226), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT30), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n227), .A2(new_n236), .A3(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n236), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n216), .A2(new_n243), .A3(new_n226), .ZN(new_n244));
  XOR2_X1   g058(.A(KEYINPUT67), .B(KEYINPUT27), .Z(new_n245));
  INV_X1    g059(.A(G237), .ZN(new_n246));
  INV_X1    g060(.A(G953), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n247), .A3(G210), .ZN(new_n248));
  XNOR2_X1  g062(.A(new_n245), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT26), .B(G101), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n249), .B(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n242), .A2(new_n244), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT31), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT28), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n244), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n239), .A2(new_n236), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n216), .A2(KEYINPUT28), .A3(new_n243), .A4(new_n226), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n251), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT31), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n242), .A2(new_n261), .A3(new_n244), .A4(new_n251), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n253), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT68), .ZN(new_n264));
  NOR2_X1   g078(.A1(G472), .A2(G902), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n264), .B1(new_n263), .B2(new_n265), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n187), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n242), .A2(new_n244), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n259), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT29), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n255), .A2(new_n251), .A3(new_n256), .A4(new_n257), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G902), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n270), .A2(KEYINPUT70), .A3(new_n271), .A4(new_n272), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n237), .A2(KEYINPUT66), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n278), .A2(new_n212), .B1(new_n195), .B2(new_n197), .ZN(new_n279));
  INV_X1    g093(.A(new_n226), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n236), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n254), .B1(new_n281), .B2(new_n244), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT71), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n259), .A2(new_n271), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n255), .A2(KEYINPUT71), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n283), .B(new_n284), .C1(new_n285), .C2(new_n282), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n275), .A2(new_n276), .A3(new_n277), .A4(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G472), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n263), .A2(KEYINPUT32), .A3(new_n265), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n268), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(G113), .B(G122), .ZN(new_n291));
  INV_X1    g105(.A(G104), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n291), .B(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G140), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G125), .ZN(new_n295));
  INV_X1    g109(.A(G125), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G140), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  XOR2_X1   g112(.A(new_n298), .B(KEYINPUT19), .Z(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n190), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT87), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n246), .A2(new_n247), .A3(G214), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n188), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n246), .A2(new_n247), .A3(G143), .A4(G214), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n208), .A3(new_n305), .ZN(new_n306));
  OR2_X1    g120(.A1(new_n306), .A2(KEYINPUT86), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n304), .A2(new_n305), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G131), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n306), .A2(KEYINPUT86), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n307), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT72), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n312), .B1(new_n295), .B2(KEYINPUT16), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT16), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n314), .A2(new_n294), .A3(KEYINPUT72), .A4(G125), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n313), .B(new_n315), .C1(new_n298), .C2(new_n314), .ZN(new_n316));
  OR2_X1    g130(.A1(new_n316), .A2(new_n190), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n299), .A2(KEYINPUT87), .A3(new_n190), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n302), .A2(new_n311), .A3(new_n317), .A4(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n309), .ZN(new_n320));
  INV_X1    g134(.A(new_n298), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n190), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n298), .A2(G146), .ZN(new_n323));
  AOI22_X1  g137(.A1(new_n320), .A2(KEYINPUT18), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n306), .B1(new_n308), .B2(KEYINPUT18), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT85), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n325), .A2(new_n326), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n324), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n293), .B1(new_n319), .B2(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n316), .B(G146), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n320), .A2(KEYINPUT17), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n331), .B(new_n332), .C1(new_n311), .C2(KEYINPUT17), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n293), .B(KEYINPUT88), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(new_n329), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT89), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT89), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n333), .A2(new_n329), .A3(new_n337), .A4(new_n334), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n330), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NOR3_X1   g153(.A1(new_n339), .A2(G475), .A3(G902), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n336), .A2(new_n338), .ZN(new_n341));
  INV_X1    g155(.A(new_n330), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT90), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT20), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n340), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G475), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n343), .A2(new_n348), .A3(new_n276), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n346), .B1(new_n339), .B2(KEYINPUT90), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n347), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(G128), .B(G143), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT13), .ZN(new_n354));
  NOR3_X1   g168(.A1(new_n220), .A2(KEYINPUT13), .A3(G143), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n355), .A2(new_n201), .ZN(new_n356));
  AOI22_X1  g170(.A1(new_n354), .A2(new_n356), .B1(new_n201), .B2(new_n353), .ZN(new_n357));
  INV_X1    g171(.A(G122), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G116), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n359), .B1(new_n230), .B2(new_n358), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n360), .A2(G107), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n360), .A2(G107), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n357), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n230), .A2(new_n358), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT14), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n365), .B(G107), .C1(KEYINPUT14), .C2(new_n360), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n366), .B1(G107), .B2(new_n360), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n353), .B(G134), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n363), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  XOR2_X1   g183(.A(KEYINPUT9), .B(G234), .Z(new_n370));
  XNOR2_X1  g184(.A(new_n370), .B(KEYINPUT74), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n371), .A2(G217), .A3(new_n247), .ZN(new_n372));
  OR2_X1    g186(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n369), .A2(new_n372), .ZN(new_n374));
  AOI21_X1  g188(.A(G902), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT91), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G478), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n378), .A2(KEYINPUT15), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  OAI22_X1  g194(.A1(new_n375), .A2(new_n376), .B1(KEYINPUT15), .B2(new_n378), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n380), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n293), .B1(new_n333), .B2(new_n329), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n383), .B1(new_n336), .B2(new_n338), .ZN(new_n384));
  OAI21_X1  g198(.A(G475), .B1(new_n384), .B2(G902), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n352), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(G110), .B(G140), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n247), .A2(G227), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n387), .B(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G107), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT3), .ZN(new_n391));
  OAI211_X1 g205(.A(G104), .B(new_n390), .C1(new_n391), .C2(KEYINPUT75), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n292), .A2(G107), .ZN(new_n393));
  XNOR2_X1  g207(.A(KEYINPUT75), .B(KEYINPUT3), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n390), .A2(G104), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n392), .B(new_n393), .C1(new_n394), .C2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G101), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n391), .A2(KEYINPUT75), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT75), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n400), .A2(KEYINPUT3), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n395), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G101), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n402), .A2(new_n403), .A3(new_n392), .A4(new_n393), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n398), .A2(KEYINPUT4), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT4), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n397), .A2(new_n406), .A3(G101), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n405), .A2(new_n198), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n395), .A2(new_n393), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G101), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n404), .A2(new_n225), .A3(KEYINPUT10), .A4(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n404), .A2(new_n225), .A3(new_n410), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT10), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n408), .A2(new_n411), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n278), .A2(new_n212), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n389), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT77), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n412), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n225), .B1(new_n404), .B2(new_n410), .ZN(new_n421));
  OAI211_X1 g235(.A(KEYINPUT12), .B(new_n237), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n421), .ZN(new_n423));
  AOI22_X1  g237(.A1(new_n278), .A2(new_n212), .B1(new_n423), .B2(new_n412), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n422), .B1(new_n424), .B2(KEYINPUT12), .ZN(new_n425));
  OAI211_X1 g239(.A(KEYINPUT77), .B(new_n389), .C1(new_n415), .C2(new_n416), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n419), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n389), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n415), .A2(new_n416), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n415), .A2(new_n416), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n427), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(G469), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(new_n433), .A3(new_n276), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n433), .A2(new_n276), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT76), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n429), .B1(new_n437), .B2(new_n417), .ZN(new_n438));
  OR2_X1    g252(.A1(new_n417), .A2(new_n437), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n430), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n425), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n428), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n440), .A2(G469), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n434), .A2(new_n436), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G221), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n446), .B1(new_n371), .B2(new_n276), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(KEYINPUT78), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT78), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n445), .A2(new_n451), .A3(new_n448), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n386), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(G214), .B1(G237), .B2(G902), .ZN(new_n454));
  XOR2_X1   g268(.A(new_n454), .B(KEYINPUT79), .Z(new_n455));
  NAND3_X1  g269(.A1(new_n195), .A2(new_n197), .A3(G125), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT82), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n456), .B(new_n457), .C1(new_n225), .C2(G125), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n195), .A2(new_n197), .A3(KEYINPUT82), .A4(G125), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(G224), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(G953), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n460), .B(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT6), .ZN(new_n465));
  XOR2_X1   g279(.A(G110), .B(G122), .Z(new_n466));
  AND3_X1   g280(.A1(new_n404), .A2(new_n235), .A3(new_n410), .ZN(new_n467));
  OAI211_X1 g281(.A(KEYINPUT5), .B(new_n229), .C1(new_n230), .C2(new_n228), .ZN(new_n468));
  OR2_X1    g282(.A1(new_n229), .A2(KEYINPUT5), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(G113), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT80), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n468), .A2(KEYINPUT80), .A3(G113), .A4(new_n469), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n467), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n405), .A2(new_n236), .A3(new_n407), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n474), .A2(KEYINPUT81), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(KEYINPUT81), .B1(new_n474), .B2(new_n475), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n466), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n474), .A2(new_n475), .ZN(new_n479));
  OR2_X1    g293(.A1(new_n479), .A2(new_n466), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n465), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT81), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n474), .A2(KEYINPUT81), .A3(new_n475), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(KEYINPUT6), .B1(new_n485), .B2(new_n466), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n464), .B1(new_n481), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT84), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n463), .A2(KEYINPUT7), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n458), .A2(new_n459), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n462), .B1(new_n458), .B2(new_n459), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT83), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n491), .A2(new_n492), .A3(KEYINPUT7), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n492), .B1(new_n491), .B2(KEYINPUT7), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n490), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  XOR2_X1   g309(.A(new_n466), .B(KEYINPUT8), .Z(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n472), .A2(new_n235), .A3(new_n473), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n404), .A2(new_n410), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n467), .A2(new_n470), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n497), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n488), .B1(new_n495), .B2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n494), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n491), .A2(new_n492), .A3(KEYINPUT7), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n502), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n506), .A2(new_n507), .A3(KEYINPUT84), .A4(new_n490), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n503), .A2(new_n508), .A3(new_n480), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n487), .A2(new_n509), .A3(new_n276), .ZN(new_n510));
  OAI21_X1  g324(.A(G210), .B1(G237), .B2(G902), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n487), .A2(new_n509), .A3(new_n276), .A4(new_n511), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n455), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(G234), .A2(G237), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(G952), .A3(new_n247), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  XOR2_X1   g332(.A(KEYINPUT21), .B(G898), .Z(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n516), .A2(G902), .A3(G953), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n518), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  AND2_X1   g338(.A1(new_n515), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n247), .A2(G221), .A3(G234), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n526), .B(KEYINPUT22), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(G137), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(KEYINPUT73), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n527), .B(new_n204), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT73), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n317), .A2(new_n322), .ZN(new_n534));
  OR3_X1    g348(.A1(new_n228), .A2(KEYINPUT23), .A3(G128), .ZN(new_n535));
  OAI21_X1  g349(.A(KEYINPUT23), .B1(new_n228), .B2(G128), .ZN(new_n536));
  AOI22_X1  g350(.A1(new_n535), .A2(new_n536), .B1(new_n228), .B2(G128), .ZN(new_n537));
  INV_X1    g351(.A(G110), .ZN(new_n538));
  XOR2_X1   g352(.A(G119), .B(G128), .Z(new_n539));
  XNOR2_X1  g353(.A(KEYINPUT24), .B(G110), .ZN(new_n540));
  AOI22_X1  g354(.A1(new_n537), .A2(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OR2_X1    g355(.A1(new_n534), .A2(new_n541), .ZN(new_n542));
  OAI22_X1  g356(.A1(new_n537), .A2(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n543));
  OR2_X1    g357(.A1(new_n331), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n533), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n542), .A2(new_n544), .A3(new_n530), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT25), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n548), .A2(new_n549), .A3(new_n276), .ZN(new_n550));
  INV_X1    g364(.A(new_n547), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n276), .B1(new_n551), .B2(new_n545), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT25), .ZN(new_n553));
  INV_X1    g367(.A(G234), .ZN(new_n554));
  OAI21_X1  g368(.A(G217), .B1(new_n554), .B2(G902), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n550), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n556), .A2(G902), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n548), .A2(new_n558), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n290), .A2(new_n453), .A3(new_n525), .A4(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT92), .B(G101), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n561), .B(new_n562), .ZN(G3));
  NAND2_X1  g377(.A1(new_n263), .A2(new_n265), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT68), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n263), .A2(new_n276), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n568), .A2(KEYINPUT93), .A3(G472), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(KEYINPUT93), .B1(new_n568), .B2(G472), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n567), .B(new_n560), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(G902), .B1(new_n427), .B2(new_n431), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n435), .B1(new_n573), .B2(new_n433), .ZN(new_n574));
  AOI211_X1 g388(.A(KEYINPUT78), .B(new_n447), .C1(new_n574), .C2(new_n444), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n451), .B1(new_n445), .B2(new_n448), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n515), .B(new_n524), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n352), .A2(new_n385), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n373), .A2(new_n374), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n374), .A2(KEYINPUT94), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(KEYINPUT33), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT33), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n373), .B(new_n374), .C1(KEYINPUT94), .C2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n581), .A2(G478), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n375), .A2(new_n378), .ZN(new_n585));
  NAND2_X1  g399(.A1(G478), .A2(G902), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n578), .A2(new_n588), .ZN(new_n589));
  NOR3_X1   g403(.A1(new_n572), .A2(new_n577), .A3(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT34), .B(G104), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(G6));
  NAND2_X1  g406(.A1(new_n568), .A2(G472), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT93), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI22_X1  g409(.A1(new_n595), .A2(new_n569), .B1(new_n565), .B2(new_n566), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n450), .A2(new_n452), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n596), .A2(new_n525), .A3(new_n560), .A4(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n340), .B(new_n346), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n381), .A2(new_n377), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n600), .B1(new_n379), .B2(new_n377), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n599), .A2(new_n601), .A3(new_n385), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(KEYINPUT35), .B(G107), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G9));
  NOR2_X1   g419(.A1(new_n533), .A2(KEYINPUT36), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n542), .A2(new_n544), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n558), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n557), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n596), .A2(new_n453), .A3(new_n525), .A4(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(KEYINPUT37), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(new_n538), .ZN(G12));
  AND2_X1   g428(.A1(new_n515), .A2(new_n611), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n517), .B1(new_n521), .B2(G900), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n602), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n290), .A2(new_n615), .A3(new_n597), .A4(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G128), .ZN(G30));
  INV_X1    g434(.A(new_n289), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(new_n567), .B2(new_n187), .ZN(new_n622));
  INV_X1    g436(.A(new_n269), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n623), .A2(new_n259), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n281), .A2(new_n244), .A3(new_n259), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n276), .ZN(new_n626));
  OAI21_X1  g440(.A(G472), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n622), .A2(KEYINPUT95), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n268), .A2(new_n289), .A3(new_n627), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT95), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  OR2_X1    g446(.A1(new_n632), .A2(KEYINPUT96), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(KEYINPUT96), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n455), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n578), .A2(new_n636), .A3(new_n601), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n616), .B(KEYINPUT39), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n597), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(new_n640), .B(KEYINPUT97), .Z(new_n641));
  INV_X1    g455(.A(KEYINPUT40), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n611), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n513), .A2(new_n514), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT38), .ZN(new_n645));
  OR2_X1    g459(.A1(new_n641), .A2(new_n642), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n638), .A2(new_n643), .A3(new_n645), .A4(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G143), .ZN(G45));
  NOR2_X1   g462(.A1(new_n575), .A2(new_n576), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n649), .B1(new_n622), .B2(new_n288), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n589), .A2(new_n617), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n650), .A2(KEYINPUT98), .A3(new_n615), .A4(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n290), .A2(new_n651), .A3(new_n615), .A4(new_n597), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT98), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G146), .ZN(G48));
  INV_X1    g471(.A(new_n434), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n573), .A2(new_n433), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n658), .A2(new_n659), .A3(new_n447), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n290), .A2(new_n525), .A3(new_n560), .A4(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n661), .A2(new_n589), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT41), .B(G113), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G15));
  NOR2_X1   g478(.A1(new_n661), .A2(new_n602), .ZN(new_n665));
  XOR2_X1   g479(.A(new_n665), .B(G116), .Z(G18));
  INV_X1    g480(.A(new_n386), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n290), .A2(new_n524), .A3(new_n667), .A4(new_n660), .ZN(new_n668));
  INV_X1    g482(.A(new_n615), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(new_n228), .ZN(G21));
  INV_X1    g485(.A(KEYINPUT99), .ZN(new_n672));
  AND3_X1   g486(.A1(new_n557), .A2(new_n672), .A3(new_n559), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n672), .B1(new_n557), .B2(new_n559), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OR2_X1    g489(.A1(new_n285), .A2(new_n282), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n251), .B1(new_n676), .B2(new_n283), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n253), .A2(new_n262), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n265), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  AND4_X1   g493(.A1(new_n593), .A2(new_n675), .A3(new_n679), .A4(new_n660), .ZN(new_n680));
  INV_X1    g494(.A(new_n644), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n637), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n680), .A2(new_n524), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G122), .ZN(G24));
  AND2_X1   g498(.A1(new_n515), .A2(new_n660), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n679), .A2(new_n593), .ZN(new_n686));
  INV_X1    g500(.A(new_n589), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n610), .A2(new_n617), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n685), .A2(new_n686), .A3(new_n687), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G125), .ZN(G27));
  INV_X1    g504(.A(KEYINPUT32), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n564), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n289), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT103), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n692), .A2(KEYINPUT103), .A3(new_n289), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n695), .A2(new_n288), .A3(new_n696), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n697), .A2(new_n675), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n440), .A2(KEYINPUT100), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n440), .A2(KEYINPUT100), .ZN(new_n700));
  OAI211_X1 g514(.A(G469), .B(new_n443), .C1(new_n699), .C2(new_n700), .ZN(new_n701));
  OR2_X1    g515(.A1(new_n701), .A2(KEYINPUT101), .ZN(new_n702));
  INV_X1    g516(.A(new_n574), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n703), .B1(new_n701), .B2(KEYINPUT101), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n447), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n687), .A2(new_n616), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n644), .A2(new_n455), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n698), .A2(KEYINPUT42), .A3(new_n705), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n705), .A2(new_n290), .A3(new_n560), .A4(new_n707), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n711), .B1(new_n712), .B2(new_n706), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G131), .ZN(G33));
  NOR3_X1   g529(.A1(new_n712), .A2(new_n602), .A3(new_n617), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT104), .B(G134), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G36));
  OAI211_X1 g532(.A(KEYINPUT45), .B(new_n443), .C1(new_n699), .C2(new_n700), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n440), .A2(new_n443), .ZN(new_n720));
  OR2_X1    g534(.A1(new_n720), .A2(KEYINPUT45), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n719), .A2(new_n721), .A3(G469), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n722), .A2(KEYINPUT46), .A3(new_n436), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT105), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT46), .ZN(new_n726));
  INV_X1    g540(.A(new_n722), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n726), .B1(new_n727), .B2(new_n435), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n722), .A2(KEYINPUT105), .A3(KEYINPUT46), .A4(new_n436), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n725), .A2(new_n728), .A3(new_n434), .A4(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n730), .A2(new_n448), .A3(new_n639), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n578), .A2(KEYINPUT43), .A3(new_n587), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n352), .A2(new_n385), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(KEYINPUT106), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n352), .A2(KEYINPUT106), .A3(new_n385), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n588), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n732), .B1(new_n736), .B2(KEYINPUT43), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n567), .B1(new_n570), .B2(new_n571), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n738), .A2(KEYINPUT107), .A3(new_n611), .ZN(new_n739));
  AOI21_X1  g553(.A(KEYINPUT107), .B1(new_n738), .B2(new_n611), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n737), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n731), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n737), .B(KEYINPUT44), .C1(new_n740), .C2(new_n739), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n744), .A2(KEYINPUT108), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n744), .A2(KEYINPUT108), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n707), .B(new_n743), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G137), .ZN(G39));
  NAND2_X1  g562(.A1(new_n730), .A2(new_n448), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT47), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n730), .A2(KEYINPUT47), .A3(new_n448), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n290), .A2(new_n560), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(new_n709), .A3(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G140), .ZN(G42));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n619), .A2(new_n689), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n758), .B1(new_n652), .B2(new_n655), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n611), .A2(new_n617), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n632), .A2(new_n682), .A3(new_n705), .A4(new_n760), .ZN(new_n761));
  AND3_X1   g575(.A1(new_n759), .A2(KEYINPUT52), .A3(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n763), .B1(new_n759), .B2(new_n761), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT109), .ZN(new_n766));
  AND4_X1   g580(.A1(new_n290), .A2(new_n453), .A3(new_n525), .A4(new_n560), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n766), .B1(new_n767), .B2(new_n590), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n561), .B(KEYINPUT109), .C1(new_n598), .C2(new_n589), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n662), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n716), .B1(new_n710), .B2(new_n713), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n733), .A2(new_n601), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n683), .B(new_n612), .C1(new_n598), .C2(new_n772), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n773), .A2(new_n665), .A3(new_n670), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n599), .A2(new_n385), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n650), .A2(new_n382), .A3(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n705), .A2(new_n687), .A3(new_n686), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n778), .A2(new_n688), .A3(new_n707), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n770), .A2(new_n771), .A3(new_n774), .A4(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n757), .B1(new_n765), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(KEYINPUT111), .ZN(new_n782));
  AND4_X1   g596(.A1(new_n771), .A2(new_n770), .A3(new_n774), .A4(new_n779), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n784));
  INV_X1    g598(.A(new_n758), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n653), .A2(new_n654), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n653), .A2(new_n654), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n785), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n761), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n784), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n759), .A2(KEYINPUT52), .A3(new_n761), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XOR2_X1   g606(.A(KEYINPUT112), .B(KEYINPUT53), .Z(new_n793));
  NAND3_X1  g607(.A1(new_n783), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT111), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n795), .B(new_n757), .C1(new_n765), .C2(new_n780), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n782), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT54), .ZN(new_n798));
  INV_X1    g612(.A(new_n793), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT52), .B1(new_n759), .B2(new_n761), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n762), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n799), .B1(new_n801), .B2(new_n780), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n788), .A2(new_n789), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n791), .B1(new_n803), .B2(new_n763), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n783), .A2(new_n804), .A3(KEYINPUT53), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n802), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n798), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(KEYINPUT113), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n658), .A2(new_n659), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(KEYINPUT115), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n751), .B(new_n752), .C1(new_n448), .C2(new_n811), .ZN(new_n812));
  AOI211_X1 g626(.A(new_n517), .B(new_n732), .C1(new_n736), .C2(KEYINPUT43), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n686), .A2(new_n675), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n813), .A2(new_n814), .A3(new_n707), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT114), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n737), .A2(new_n518), .A3(new_n814), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(KEYINPUT114), .A3(new_n707), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n812), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n645), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n821), .A2(new_n455), .A3(new_n660), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT116), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n821), .A2(KEYINPUT116), .A3(new_n455), .A4(new_n660), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n813), .A2(new_n824), .A3(new_n814), .A4(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT50), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n818), .A2(KEYINPUT50), .A3(new_n824), .A4(new_n825), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n707), .A2(new_n660), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n813), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n832), .A2(new_n611), .A3(new_n686), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n820), .A2(new_n830), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n831), .A2(new_n560), .ZN(new_n835));
  AOI211_X1 g649(.A(new_n517), .B(new_n835), .C1(new_n633), .C2(new_n634), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n836), .A2(new_n733), .A3(new_n587), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT117), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n836), .A2(KEYINPUT117), .A3(new_n733), .A4(new_n587), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n834), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI211_X1 g655(.A(G952), .B(new_n247), .C1(new_n841), .C2(KEYINPUT51), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT51), .ZN(new_n843));
  AOI211_X1 g657(.A(new_n843), .B(new_n834), .C1(new_n839), .C2(new_n840), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n836), .A2(new_n687), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n832), .A2(new_n698), .ZN(new_n846));
  XOR2_X1   g660(.A(new_n846), .B(KEYINPUT48), .Z(new_n847));
  NOR4_X1   g661(.A1(new_n842), .A2(new_n844), .A3(new_n845), .A4(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT113), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n798), .A2(new_n849), .A3(new_n807), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n818), .A2(new_n685), .ZN(new_n851));
  XOR2_X1   g665(.A(new_n851), .B(KEYINPUT118), .Z(new_n852));
  NAND4_X1  g666(.A1(new_n809), .A2(new_n848), .A3(new_n850), .A4(new_n852), .ZN(new_n853));
  OR2_X1    g667(.A1(G952), .A2(G953), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n635), .A2(new_n636), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n856), .A2(new_n645), .A3(new_n736), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n810), .B(KEYINPUT49), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n857), .A2(new_n448), .A3(new_n675), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n855), .A2(new_n859), .ZN(G75));
  NOR3_X1   g674(.A1(new_n765), .A2(new_n757), .A3(new_n780), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n793), .B1(new_n783), .B2(new_n792), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n863), .A2(new_n276), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT56), .B1(new_n864), .B2(G210), .ZN(new_n865));
  OR2_X1    g679(.A1(new_n481), .A2(new_n486), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(new_n464), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n867), .B(KEYINPUT55), .Z(new_n868));
  XNOR2_X1  g682(.A(new_n865), .B(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n247), .A2(G952), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(G51));
  OAI21_X1  g685(.A(KEYINPUT54), .B1(new_n861), .B2(new_n862), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT119), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n872), .A2(new_n873), .A3(new_n807), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n863), .A2(KEYINPUT119), .A3(new_n806), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n435), .B(KEYINPUT57), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT120), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n877), .A2(new_n878), .A3(new_n432), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n878), .B1(new_n877), .B2(new_n432), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n864), .A2(new_n727), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n882), .B(KEYINPUT121), .Z(new_n883));
  AOI21_X1  g697(.A(new_n870), .B1(new_n881), .B2(new_n883), .ZN(G54));
  NAND3_X1  g698(.A1(new_n864), .A2(KEYINPUT58), .A3(G475), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(new_n339), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n886), .A2(new_n870), .ZN(G60));
  NAND2_X1  g701(.A1(new_n874), .A2(new_n875), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n581), .A2(new_n583), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n586), .B(KEYINPUT59), .Z(new_n890));
  NOR3_X1   g704(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n890), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n802), .A2(new_n805), .A3(new_n806), .ZN(new_n893));
  AOI211_X1 g707(.A(KEYINPUT113), .B(new_n893), .C1(new_n797), .C2(KEYINPUT54), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n849), .B1(new_n798), .B2(new_n807), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n892), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AOI211_X1 g710(.A(new_n870), .B(new_n891), .C1(new_n896), .C2(new_n889), .ZN(G63));
  NAND2_X1  g711(.A1(G217), .A2(G902), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT60), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n802), .B2(new_n805), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(new_n608), .ZN(new_n901));
  INV_X1    g715(.A(new_n870), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n901), .B(new_n902), .C1(new_n548), .C2(new_n900), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT122), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT61), .ZN(G66));
  NAND2_X1  g720(.A1(new_n770), .A2(new_n774), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT123), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n247), .B1(new_n519), .B2(G224), .ZN(new_n909));
  AOI22_X1  g723(.A1(new_n907), .A2(new_n247), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n910), .B1(new_n908), .B2(new_n909), .ZN(new_n911));
  INV_X1    g725(.A(G898), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n866), .B1(new_n912), .B2(G953), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n911), .B(new_n913), .Z(G69));
  AOI21_X1  g728(.A(new_n247), .B1(G227), .B2(G900), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n227), .A2(new_n241), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(new_n299), .ZN(new_n917));
  NAND2_X1  g731(.A1(G900), .A2(G953), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n747), .A2(new_n755), .A3(new_n759), .A4(new_n771), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n698), .A2(new_n682), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n731), .A2(new_n920), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n917), .B(new_n918), .C1(new_n922), .C2(G953), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n915), .B1(new_n923), .B2(KEYINPUT125), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n917), .B(KEYINPUT124), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n290), .A2(new_n560), .A3(new_n707), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n772), .A2(new_n589), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n641), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n747), .A2(new_n755), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n647), .A2(new_n759), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT62), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n647), .A2(KEYINPUT62), .A3(new_n759), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n929), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n925), .B1(new_n934), .B2(G953), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n923), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n924), .B(new_n936), .Z(G72));
  NAND2_X1  g751(.A1(G472), .A2(G902), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT63), .Z(new_n939));
  OAI21_X1  g753(.A(new_n939), .B1(new_n922), .B2(new_n907), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n940), .A2(new_n623), .A3(new_n259), .ZN(new_n941));
  INV_X1    g755(.A(new_n939), .ZN(new_n942));
  INV_X1    g756(.A(new_n907), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n942), .B1(new_n934), .B2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n624), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n941), .B(new_n902), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n942), .B1(new_n270), .B2(new_n252), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT126), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n797), .A2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(KEYINPUT127), .B1(new_n946), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n944), .A2(new_n945), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n952), .A2(new_n870), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n953), .A2(new_n954), .A3(new_n941), .A4(new_n949), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n951), .A2(new_n955), .ZN(G57));
endmodule


