

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U555 ( .A1(G543), .A2(G651), .ZN(n643) );
  NOR2_X2 U556 ( .A1(n721), .A2(n720), .ZN(n722) );
  AND2_X1 U557 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U558 ( .A1(n812), .A2(n802), .ZN(n522) );
  INV_X1 U559 ( .A(KEYINPUT32), .ZN(n741) );
  NAND2_X1 U560 ( .A1(n771), .A2(n769), .ZN(n729) );
  XNOR2_X1 U561 ( .A(KEYINPUT72), .B(KEYINPUT4), .ZN(n551) );
  AND2_X1 U562 ( .A1(G160), .A2(G40), .ZN(n769) );
  XNOR2_X1 U563 ( .A(n552), .B(n551), .ZN(n554) );
  NOR2_X1 U564 ( .A1(G164), .A2(G1384), .ZN(n771) );
  INV_X1 U565 ( .A(KEYINPUT17), .ZN(n523) );
  NAND2_X1 U566 ( .A1(n803), .A2(n522), .ZN(n804) );
  NOR2_X1 U567 ( .A1(G543), .A2(n543), .ZN(n539) );
  XNOR2_X1 U568 ( .A(n524), .B(n523), .ZN(n875) );
  OR2_X1 U569 ( .A1(n805), .A2(n804), .ZN(n820) );
  XOR2_X1 U570 ( .A(KEYINPUT15), .B(n586), .Z(n977) );
  NOR2_X1 U571 ( .A1(G651), .A2(n634), .ZN(n647) );
  NAND2_X1 U572 ( .A1(n875), .A2(G138), .ZN(n526) );
  NOR2_X1 U573 ( .A1(G2105), .A2(G2104), .ZN(n524) );
  INV_X1 U574 ( .A(G2104), .ZN(n527) );
  NOR2_X4 U575 ( .A1(G2105), .A2(n527), .ZN(n876) );
  NAND2_X1 U576 ( .A1(G102), .A2(n876), .ZN(n525) );
  NAND2_X1 U577 ( .A1(n526), .A2(n525), .ZN(n531) );
  AND2_X1 U578 ( .A1(n527), .A2(G2105), .ZN(n871) );
  NAND2_X1 U579 ( .A1(G126), .A2(n871), .ZN(n529) );
  AND2_X1 U580 ( .A1(G2105), .A2(G2104), .ZN(n872) );
  NAND2_X1 U581 ( .A1(G114), .A2(n872), .ZN(n528) );
  NAND2_X1 U582 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U583 ( .A1(n531), .A2(n530), .ZN(G164) );
  NAND2_X1 U584 ( .A1(n875), .A2(G137), .ZN(n534) );
  NAND2_X1 U585 ( .A1(G101), .A2(n876), .ZN(n532) );
  XOR2_X1 U586 ( .A(KEYINPUT23), .B(n532), .Z(n533) );
  NAND2_X1 U587 ( .A1(n534), .A2(n533), .ZN(n538) );
  NAND2_X1 U588 ( .A1(G125), .A2(n871), .ZN(n536) );
  NAND2_X1 U589 ( .A1(G113), .A2(n872), .ZN(n535) );
  NAND2_X1 U590 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U591 ( .A1(n538), .A2(n537), .ZN(G160) );
  AND2_X1 U592 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U593 ( .A(G57), .ZN(G237) );
  XOR2_X1 U594 ( .A(G543), .B(KEYINPUT0), .Z(n634) );
  NAND2_X1 U595 ( .A1(G50), .A2(n647), .ZN(n541) );
  INV_X1 U596 ( .A(G651), .ZN(n543) );
  XOR2_X1 U597 ( .A(KEYINPUT1), .B(n539), .Z(n641) );
  NAND2_X1 U598 ( .A1(G62), .A2(n641), .ZN(n540) );
  NAND2_X1 U599 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U600 ( .A(KEYINPUT81), .B(n542), .ZN(n547) );
  NAND2_X1 U601 ( .A1(G88), .A2(n643), .ZN(n545) );
  NOR2_X1 U602 ( .A1(n634), .A2(n543), .ZN(n644) );
  NAND2_X1 U603 ( .A1(G75), .A2(n644), .ZN(n544) );
  AND2_X1 U604 ( .A1(n545), .A2(n544), .ZN(n546) );
  NAND2_X1 U605 ( .A1(n547), .A2(n546), .ZN(G303) );
  NAND2_X1 U606 ( .A1(G51), .A2(n647), .ZN(n549) );
  NAND2_X1 U607 ( .A1(G63), .A2(n641), .ZN(n548) );
  NAND2_X1 U608 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U609 ( .A(KEYINPUT6), .B(n550), .ZN(n557) );
  NAND2_X1 U610 ( .A1(G89), .A2(n643), .ZN(n552) );
  NAND2_X1 U611 ( .A1(G76), .A2(n644), .ZN(n553) );
  NAND2_X1 U612 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U613 ( .A(n555), .B(KEYINPUT5), .Z(n556) );
  NOR2_X1 U614 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U615 ( .A(KEYINPUT7), .B(n558), .Z(n559) );
  XOR2_X1 U616 ( .A(KEYINPUT73), .B(n559), .Z(G168) );
  XOR2_X1 U617 ( .A(G168), .B(KEYINPUT8), .Z(n560) );
  XNOR2_X1 U618 ( .A(KEYINPUT74), .B(n560), .ZN(G286) );
  NAND2_X1 U619 ( .A1(G7), .A2(G661), .ZN(n561) );
  XNOR2_X1 U620 ( .A(n561), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U621 ( .A(G223), .ZN(n822) );
  NAND2_X1 U622 ( .A1(n822), .A2(G567), .ZN(n562) );
  XOR2_X1 U623 ( .A(KEYINPUT11), .B(n562), .Z(G234) );
  XOR2_X1 U624 ( .A(G860), .B(KEYINPUT70), .Z(n601) );
  NAND2_X1 U625 ( .A1(G56), .A2(n641), .ZN(n563) );
  XOR2_X1 U626 ( .A(KEYINPUT14), .B(n563), .Z(n569) );
  NAND2_X1 U627 ( .A1(n643), .A2(G81), .ZN(n564) );
  XNOR2_X1 U628 ( .A(n564), .B(KEYINPUT12), .ZN(n566) );
  NAND2_X1 U629 ( .A1(G68), .A2(n644), .ZN(n565) );
  NAND2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U631 ( .A(KEYINPUT13), .B(n567), .Z(n568) );
  NOR2_X1 U632 ( .A1(n569), .A2(n568), .ZN(n571) );
  NAND2_X1 U633 ( .A1(n647), .A2(G43), .ZN(n570) );
  NAND2_X1 U634 ( .A1(n571), .A2(n570), .ZN(n985) );
  OR2_X1 U635 ( .A1(n601), .A2(n985), .ZN(G153) );
  NAND2_X1 U636 ( .A1(n643), .A2(G90), .ZN(n572) );
  XOR2_X1 U637 ( .A(KEYINPUT67), .B(n572), .Z(n574) );
  NAND2_X1 U638 ( .A1(n644), .A2(G77), .ZN(n573) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(KEYINPUT9), .B(n575), .ZN(n579) );
  NAND2_X1 U641 ( .A1(G52), .A2(n647), .ZN(n577) );
  NAND2_X1 U642 ( .A1(G64), .A2(n641), .ZN(n576) );
  AND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(G301) );
  NAND2_X1 U645 ( .A1(G92), .A2(n643), .ZN(n581) );
  NAND2_X1 U646 ( .A1(G79), .A2(n644), .ZN(n580) );
  NAND2_X1 U647 ( .A1(n581), .A2(n580), .ZN(n585) );
  NAND2_X1 U648 ( .A1(G54), .A2(n647), .ZN(n583) );
  NAND2_X1 U649 ( .A1(G66), .A2(n641), .ZN(n582) );
  NAND2_X1 U650 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U651 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U652 ( .A1(n977), .A2(G868), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n587), .B(KEYINPUT71), .ZN(n589) );
  NAND2_X1 U654 ( .A1(G868), .A2(G301), .ZN(n588) );
  NAND2_X1 U655 ( .A1(n589), .A2(n588), .ZN(G284) );
  NAND2_X1 U656 ( .A1(G91), .A2(n643), .ZN(n591) );
  NAND2_X1 U657 ( .A1(G78), .A2(n644), .ZN(n590) );
  NAND2_X1 U658 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U659 ( .A(KEYINPUT68), .B(n592), .ZN(n595) );
  NAND2_X1 U660 ( .A1(G65), .A2(n641), .ZN(n593) );
  XNOR2_X1 U661 ( .A(KEYINPUT69), .B(n593), .ZN(n594) );
  NOR2_X1 U662 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U663 ( .A1(n647), .A2(G53), .ZN(n596) );
  NAND2_X1 U664 ( .A1(n597), .A2(n596), .ZN(G299) );
  INV_X1 U665 ( .A(G868), .ZN(n662) );
  NAND2_X1 U666 ( .A1(G299), .A2(n662), .ZN(n599) );
  NAND2_X1 U667 ( .A1(G868), .A2(G286), .ZN(n598) );
  NAND2_X1 U668 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U669 ( .A(KEYINPUT75), .B(n600), .Z(G297) );
  NAND2_X1 U670 ( .A1(n601), .A2(G559), .ZN(n602) );
  NAND2_X1 U671 ( .A1(n602), .A2(n977), .ZN(n603) );
  XNOR2_X1 U672 ( .A(n603), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U673 ( .A1(G868), .A2(n985), .ZN(n604) );
  XNOR2_X1 U674 ( .A(KEYINPUT76), .B(n604), .ZN(n607) );
  NAND2_X1 U675 ( .A1(G868), .A2(n977), .ZN(n605) );
  NOR2_X1 U676 ( .A1(G559), .A2(n605), .ZN(n606) );
  NOR2_X1 U677 ( .A1(n607), .A2(n606), .ZN(G282) );
  XNOR2_X1 U678 ( .A(G2100), .B(KEYINPUT79), .ZN(n618) );
  NAND2_X1 U679 ( .A1(G123), .A2(n871), .ZN(n608) );
  XOR2_X1 U680 ( .A(KEYINPUT18), .B(n608), .Z(n609) );
  XNOR2_X1 U681 ( .A(n609), .B(KEYINPUT77), .ZN(n611) );
  NAND2_X1 U682 ( .A1(G135), .A2(n875), .ZN(n610) );
  NAND2_X1 U683 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U684 ( .A(KEYINPUT78), .B(n612), .ZN(n616) );
  NAND2_X1 U685 ( .A1(G99), .A2(n876), .ZN(n614) );
  NAND2_X1 U686 ( .A1(G111), .A2(n872), .ZN(n613) );
  NAND2_X1 U687 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U688 ( .A1(n616), .A2(n615), .ZN(n930) );
  XNOR2_X1 U689 ( .A(n930), .B(G2096), .ZN(n617) );
  NAND2_X1 U690 ( .A1(n618), .A2(n617), .ZN(G156) );
  NAND2_X1 U691 ( .A1(G559), .A2(n977), .ZN(n619) );
  XNOR2_X1 U692 ( .A(n985), .B(n619), .ZN(n659) );
  NOR2_X1 U693 ( .A1(n659), .A2(G860), .ZN(n626) );
  NAND2_X1 U694 ( .A1(G55), .A2(n647), .ZN(n621) );
  NAND2_X1 U695 ( .A1(G67), .A2(n641), .ZN(n620) );
  NAND2_X1 U696 ( .A1(n621), .A2(n620), .ZN(n625) );
  NAND2_X1 U697 ( .A1(G93), .A2(n643), .ZN(n623) );
  NAND2_X1 U698 ( .A1(G80), .A2(n644), .ZN(n622) );
  NAND2_X1 U699 ( .A1(n623), .A2(n622), .ZN(n624) );
  OR2_X1 U700 ( .A1(n625), .A2(n624), .ZN(n661) );
  XOR2_X1 U701 ( .A(n626), .B(n661), .Z(G145) );
  NAND2_X1 U702 ( .A1(G86), .A2(n643), .ZN(n628) );
  NAND2_X1 U703 ( .A1(G48), .A2(n647), .ZN(n627) );
  NAND2_X1 U704 ( .A1(n628), .A2(n627), .ZN(n631) );
  NAND2_X1 U705 ( .A1(n644), .A2(G73), .ZN(n629) );
  XOR2_X1 U706 ( .A(KEYINPUT2), .B(n629), .Z(n630) );
  NOR2_X1 U707 ( .A1(n631), .A2(n630), .ZN(n633) );
  NAND2_X1 U708 ( .A1(n641), .A2(G61), .ZN(n632) );
  NAND2_X1 U709 ( .A1(n633), .A2(n632), .ZN(G305) );
  NAND2_X1 U710 ( .A1(G74), .A2(G651), .ZN(n639) );
  NAND2_X1 U711 ( .A1(G49), .A2(n647), .ZN(n636) );
  NAND2_X1 U712 ( .A1(G87), .A2(n634), .ZN(n635) );
  NAND2_X1 U713 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U714 ( .A1(n641), .A2(n637), .ZN(n638) );
  NAND2_X1 U715 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U716 ( .A(n640), .B(KEYINPUT80), .ZN(G288) );
  NAND2_X1 U717 ( .A1(n641), .A2(G60), .ZN(n642) );
  XNOR2_X1 U718 ( .A(n642), .B(KEYINPUT64), .ZN(n652) );
  NAND2_X1 U719 ( .A1(G85), .A2(n643), .ZN(n646) );
  NAND2_X1 U720 ( .A1(G72), .A2(n644), .ZN(n645) );
  NAND2_X1 U721 ( .A1(n646), .A2(n645), .ZN(n650) );
  NAND2_X1 U722 ( .A1(G47), .A2(n647), .ZN(n648) );
  XNOR2_X1 U723 ( .A(KEYINPUT65), .B(n648), .ZN(n649) );
  NOR2_X1 U724 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U725 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U726 ( .A(KEYINPUT66), .B(n653), .ZN(G290) );
  INV_X1 U727 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U728 ( .A(G305), .B(G288), .ZN(n655) );
  XNOR2_X1 U729 ( .A(G290), .B(G166), .ZN(n654) );
  XNOR2_X1 U730 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U731 ( .A(n656), .B(n661), .ZN(n658) );
  INV_X1 U732 ( .A(G299), .ZN(n970) );
  XNOR2_X1 U733 ( .A(n970), .B(KEYINPUT19), .ZN(n657) );
  XNOR2_X1 U734 ( .A(n658), .B(n657), .ZN(n890) );
  XOR2_X1 U735 ( .A(n659), .B(n890), .Z(n660) );
  NAND2_X1 U736 ( .A1(n660), .A2(G868), .ZN(n664) );
  NAND2_X1 U737 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U738 ( .A1(n664), .A2(n663), .ZN(G295) );
  NAND2_X1 U739 ( .A1(G2084), .A2(G2078), .ZN(n665) );
  XOR2_X1 U740 ( .A(KEYINPUT20), .B(n665), .Z(n666) );
  NAND2_X1 U741 ( .A1(G2090), .A2(n666), .ZN(n667) );
  XNOR2_X1 U742 ( .A(KEYINPUT21), .B(n667), .ZN(n668) );
  NAND2_X1 U743 ( .A1(n668), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U744 ( .A(KEYINPUT82), .B(G44), .ZN(n669) );
  XNOR2_X1 U745 ( .A(n669), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U746 ( .A1(G483), .A2(G661), .ZN(n678) );
  XOR2_X1 U747 ( .A(KEYINPUT83), .B(KEYINPUT22), .Z(n671) );
  NAND2_X1 U748 ( .A1(G132), .A2(G82), .ZN(n670) );
  XNOR2_X1 U749 ( .A(n671), .B(n670), .ZN(n672) );
  NOR2_X1 U750 ( .A1(G218), .A2(n672), .ZN(n673) );
  NAND2_X1 U751 ( .A1(G96), .A2(n673), .ZN(n827) );
  NAND2_X1 U752 ( .A1(n827), .A2(G2106), .ZN(n677) );
  NAND2_X1 U753 ( .A1(G108), .A2(G120), .ZN(n674) );
  NOR2_X1 U754 ( .A1(G237), .A2(n674), .ZN(n675) );
  NAND2_X1 U755 ( .A1(G69), .A2(n675), .ZN(n828) );
  NAND2_X1 U756 ( .A1(n828), .A2(G567), .ZN(n676) );
  NAND2_X1 U757 ( .A1(n677), .A2(n676), .ZN(n829) );
  NOR2_X1 U758 ( .A1(n678), .A2(n829), .ZN(n679) );
  XNOR2_X1 U759 ( .A(n679), .B(KEYINPUT84), .ZN(n826) );
  NAND2_X1 U760 ( .A1(G36), .A2(n826), .ZN(G176) );
  INV_X1 U761 ( .A(G301), .ZN(G171) );
  NAND2_X1 U762 ( .A1(G8), .A2(n729), .ZN(n763) );
  NOR2_X1 U763 ( .A1(G1976), .A2(G288), .ZN(n751) );
  NOR2_X1 U764 ( .A1(G1971), .A2(G303), .ZN(n680) );
  NOR2_X1 U765 ( .A1(n751), .A2(n680), .ZN(n971) );
  INV_X1 U766 ( .A(n971), .ZN(n745) );
  NOR2_X1 U767 ( .A1(G1966), .A2(n763), .ZN(n724) );
  NOR2_X1 U768 ( .A1(G2084), .A2(n729), .ZN(n725) );
  NOR2_X1 U769 ( .A1(n724), .A2(n725), .ZN(n681) );
  NAND2_X1 U770 ( .A1(G8), .A2(n681), .ZN(n682) );
  XNOR2_X1 U771 ( .A(KEYINPUT30), .B(n682), .ZN(n683) );
  NOR2_X1 U772 ( .A1(G168), .A2(n683), .ZN(n688) );
  XOR2_X1 U773 ( .A(G2078), .B(KEYINPUT25), .Z(n948) );
  NOR2_X1 U774 ( .A1(n948), .A2(n729), .ZN(n684) );
  XNOR2_X1 U775 ( .A(n684), .B(KEYINPUT91), .ZN(n686) );
  INV_X1 U776 ( .A(n729), .ZN(n699) );
  OR2_X1 U777 ( .A1(G1961), .A2(n699), .ZN(n685) );
  NAND2_X1 U778 ( .A1(n686), .A2(n685), .ZN(n719) );
  NOR2_X1 U779 ( .A1(G171), .A2(n719), .ZN(n687) );
  NOR2_X1 U780 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U781 ( .A(KEYINPUT31), .B(n689), .ZN(n734) );
  INV_X1 U782 ( .A(n729), .ZN(n690) );
  NAND2_X1 U783 ( .A1(n690), .A2(G2072), .ZN(n691) );
  XNOR2_X1 U784 ( .A(n691), .B(KEYINPUT27), .ZN(n693) );
  AND2_X1 U785 ( .A1(G1956), .A2(n729), .ZN(n692) );
  NOR2_X1 U786 ( .A1(n693), .A2(n692), .ZN(n712) );
  NOR2_X1 U787 ( .A1(n970), .A2(n712), .ZN(n694) );
  XOR2_X1 U788 ( .A(n694), .B(KEYINPUT28), .Z(n716) );
  AND2_X1 U789 ( .A1(n729), .A2(G1348), .ZN(n696) );
  AND2_X1 U790 ( .A1(n699), .A2(G2067), .ZN(n695) );
  NOR2_X1 U791 ( .A1(n696), .A2(n695), .ZN(n709) );
  NAND2_X1 U792 ( .A1(n709), .A2(n977), .ZN(n708) );
  AND2_X1 U793 ( .A1(n729), .A2(G1341), .ZN(n701) );
  AND2_X1 U794 ( .A1(n701), .A2(KEYINPUT26), .ZN(n697) );
  NOR2_X1 U795 ( .A1(KEYINPUT92), .A2(n697), .ZN(n698) );
  NOR2_X1 U796 ( .A1(n698), .A2(n985), .ZN(n706) );
  NAND2_X1 U797 ( .A1(G1996), .A2(n699), .ZN(n700) );
  XNOR2_X1 U798 ( .A(KEYINPUT26), .B(n700), .ZN(n703) );
  INV_X1 U799 ( .A(n701), .ZN(n702) );
  NAND2_X1 U800 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U801 ( .A1(n704), .A2(KEYINPUT92), .ZN(n705) );
  NAND2_X1 U802 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U803 ( .A1(n708), .A2(n707), .ZN(n711) );
  OR2_X1 U804 ( .A1(n709), .A2(n977), .ZN(n710) );
  NAND2_X1 U805 ( .A1(n711), .A2(n710), .ZN(n714) );
  NAND2_X1 U806 ( .A1(n970), .A2(n712), .ZN(n713) );
  NAND2_X1 U807 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U808 ( .A1(n716), .A2(n715), .ZN(n718) );
  XOR2_X1 U809 ( .A(KEYINPUT29), .B(KEYINPUT93), .Z(n717) );
  XNOR2_X1 U810 ( .A(n718), .B(n717), .ZN(n721) );
  AND2_X1 U811 ( .A1(n719), .A2(G171), .ZN(n720) );
  XNOR2_X1 U812 ( .A(n722), .B(KEYINPUT94), .ZN(n736) );
  NOR2_X1 U813 ( .A1(n734), .A2(n736), .ZN(n723) );
  NOR2_X1 U814 ( .A1(n724), .A2(n723), .ZN(n727) );
  NAND2_X1 U815 ( .A1(G8), .A2(n725), .ZN(n726) );
  NAND2_X1 U816 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U817 ( .A(KEYINPUT95), .B(n728), .ZN(n744) );
  NOR2_X1 U818 ( .A1(G1971), .A2(n763), .ZN(n731) );
  NOR2_X1 U819 ( .A1(G2090), .A2(n729), .ZN(n730) );
  NOR2_X1 U820 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U821 ( .A(n732), .B(KEYINPUT96), .ZN(n733) );
  AND2_X1 U822 ( .A1(n733), .A2(G303), .ZN(n737) );
  OR2_X1 U823 ( .A1(n734), .A2(n737), .ZN(n735) );
  OR2_X1 U824 ( .A1(n736), .A2(n735), .ZN(n739) );
  OR2_X1 U825 ( .A1(n737), .A2(G286), .ZN(n738) );
  NAND2_X1 U826 ( .A1(n740), .A2(G8), .ZN(n742) );
  XNOR2_X1 U827 ( .A(n742), .B(n741), .ZN(n743) );
  NOR2_X1 U828 ( .A1(n744), .A2(n743), .ZN(n756) );
  OR2_X1 U829 ( .A1(n745), .A2(n756), .ZN(n747) );
  NAND2_X1 U830 ( .A1(G288), .A2(G1976), .ZN(n746) );
  XOR2_X1 U831 ( .A(KEYINPUT97), .B(n746), .Z(n973) );
  NAND2_X1 U832 ( .A1(n747), .A2(n973), .ZN(n748) );
  XNOR2_X1 U833 ( .A(KEYINPUT98), .B(n748), .ZN(n749) );
  NOR2_X1 U834 ( .A1(n763), .A2(n749), .ZN(n750) );
  NOR2_X1 U835 ( .A1(KEYINPUT33), .A2(n750), .ZN(n754) );
  NAND2_X1 U836 ( .A1(n751), .A2(KEYINPUT33), .ZN(n752) );
  NOR2_X1 U837 ( .A1(n752), .A2(n763), .ZN(n753) );
  NOR2_X1 U838 ( .A1(n754), .A2(n753), .ZN(n755) );
  XOR2_X1 U839 ( .A(G1981), .B(G305), .Z(n967) );
  AND2_X1 U840 ( .A1(n755), .A2(n967), .ZN(n767) );
  NAND2_X1 U841 ( .A1(G166), .A2(G8), .ZN(n757) );
  NOR2_X1 U842 ( .A1(G2090), .A2(n757), .ZN(n758) );
  NOR2_X1 U843 ( .A1(n756), .A2(n758), .ZN(n759) );
  XNOR2_X1 U844 ( .A(n759), .B(KEYINPUT99), .ZN(n760) );
  NAND2_X1 U845 ( .A1(n760), .A2(n763), .ZN(n765) );
  NOR2_X1 U846 ( .A1(G1981), .A2(G305), .ZN(n761) );
  XOR2_X1 U847 ( .A(n761), .B(KEYINPUT24), .Z(n762) );
  OR2_X1 U848 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U849 ( .A1(n765), .A2(n764), .ZN(n766) );
  NOR2_X1 U850 ( .A1(n767), .A2(n766), .ZN(n805) );
  XOR2_X1 U851 ( .A(G1986), .B(G290), .Z(n768) );
  XNOR2_X1 U852 ( .A(KEYINPUT85), .B(n768), .ZN(n981) );
  INV_X1 U853 ( .A(n769), .ZN(n770) );
  NOR2_X1 U854 ( .A1(n771), .A2(n770), .ZN(n817) );
  NAND2_X1 U855 ( .A1(n981), .A2(n817), .ZN(n803) );
  XNOR2_X1 U856 ( .A(KEYINPUT87), .B(KEYINPUT36), .ZN(n782) );
  NAND2_X1 U857 ( .A1(G128), .A2(n871), .ZN(n773) );
  NAND2_X1 U858 ( .A1(G116), .A2(n872), .ZN(n772) );
  NAND2_X1 U859 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U860 ( .A(KEYINPUT35), .B(n774), .ZN(n780) );
  NAND2_X1 U861 ( .A1(n875), .A2(G140), .ZN(n775) );
  XNOR2_X1 U862 ( .A(n775), .B(KEYINPUT86), .ZN(n777) );
  NAND2_X1 U863 ( .A1(G104), .A2(n876), .ZN(n776) );
  NAND2_X1 U864 ( .A1(n777), .A2(n776), .ZN(n778) );
  XOR2_X1 U865 ( .A(KEYINPUT34), .B(n778), .Z(n779) );
  NAND2_X1 U866 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U867 ( .A(n782), .B(n781), .ZN(n868) );
  XNOR2_X1 U868 ( .A(KEYINPUT37), .B(G2067), .ZN(n815) );
  NOR2_X1 U869 ( .A1(n868), .A2(n815), .ZN(n922) );
  NAND2_X1 U870 ( .A1(n817), .A2(n922), .ZN(n812) );
  NAND2_X1 U871 ( .A1(G131), .A2(n875), .ZN(n784) );
  NAND2_X1 U872 ( .A1(G119), .A2(n871), .ZN(n783) );
  NAND2_X1 U873 ( .A1(n784), .A2(n783), .ZN(n787) );
  NAND2_X1 U874 ( .A1(n876), .A2(G95), .ZN(n785) );
  XOR2_X1 U875 ( .A(KEYINPUT88), .B(n785), .Z(n786) );
  NOR2_X1 U876 ( .A1(n787), .A2(n786), .ZN(n789) );
  NAND2_X1 U877 ( .A1(n872), .A2(G107), .ZN(n788) );
  NAND2_X1 U878 ( .A1(n789), .A2(n788), .ZN(n854) );
  NAND2_X1 U879 ( .A1(G1991), .A2(n854), .ZN(n790) );
  XNOR2_X1 U880 ( .A(n790), .B(KEYINPUT89), .ZN(n800) );
  XOR2_X1 U881 ( .A(KEYINPUT38), .B(KEYINPUT90), .Z(n792) );
  NAND2_X1 U882 ( .A1(G105), .A2(n876), .ZN(n791) );
  XNOR2_X1 U883 ( .A(n792), .B(n791), .ZN(n796) );
  NAND2_X1 U884 ( .A1(G141), .A2(n875), .ZN(n794) );
  NAND2_X1 U885 ( .A1(G117), .A2(n872), .ZN(n793) );
  NAND2_X1 U886 ( .A1(n794), .A2(n793), .ZN(n795) );
  NOR2_X1 U887 ( .A1(n796), .A2(n795), .ZN(n798) );
  NAND2_X1 U888 ( .A1(n871), .A2(G129), .ZN(n797) );
  NAND2_X1 U889 ( .A1(n798), .A2(n797), .ZN(n855) );
  AND2_X1 U890 ( .A1(G1996), .A2(n855), .ZN(n799) );
  NOR2_X1 U891 ( .A1(n800), .A2(n799), .ZN(n933) );
  INV_X1 U892 ( .A(n817), .ZN(n801) );
  NOR2_X1 U893 ( .A1(n933), .A2(n801), .ZN(n808) );
  INV_X1 U894 ( .A(n808), .ZN(n802) );
  NOR2_X1 U895 ( .A1(G1996), .A2(n855), .ZN(n925) );
  NOR2_X1 U896 ( .A1(G1986), .A2(G290), .ZN(n806) );
  NOR2_X1 U897 ( .A1(G1991), .A2(n854), .ZN(n929) );
  NOR2_X1 U898 ( .A1(n806), .A2(n929), .ZN(n807) );
  NOR2_X1 U899 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U900 ( .A(n809), .B(KEYINPUT100), .ZN(n810) );
  NOR2_X1 U901 ( .A1(n925), .A2(n810), .ZN(n811) );
  XNOR2_X1 U902 ( .A(n811), .B(KEYINPUT39), .ZN(n813) );
  NAND2_X1 U903 ( .A1(n813), .A2(n812), .ZN(n814) );
  XOR2_X1 U904 ( .A(KEYINPUT101), .B(n814), .Z(n816) );
  NAND2_X1 U905 ( .A1(n868), .A2(n815), .ZN(n919) );
  NAND2_X1 U906 ( .A1(n816), .A2(n919), .ZN(n818) );
  NAND2_X1 U907 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U908 ( .A1(n820), .A2(n819), .ZN(n821) );
  XNOR2_X1 U909 ( .A(n821), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U910 ( .A1(n822), .A2(G2106), .ZN(n823) );
  XNOR2_X1 U911 ( .A(n823), .B(KEYINPUT104), .ZN(G217) );
  AND2_X1 U912 ( .A1(G15), .A2(G2), .ZN(n824) );
  NAND2_X1 U913 ( .A1(G661), .A2(n824), .ZN(G259) );
  NAND2_X1 U914 ( .A1(G3), .A2(G1), .ZN(n825) );
  NAND2_X1 U915 ( .A1(n826), .A2(n825), .ZN(G188) );
  XNOR2_X1 U916 ( .A(G120), .B(KEYINPUT105), .ZN(G236) );
  INV_X1 U918 ( .A(G132), .ZN(G219) );
  INV_X1 U919 ( .A(G108), .ZN(G238) );
  INV_X1 U920 ( .A(G96), .ZN(G221) );
  INV_X1 U921 ( .A(G82), .ZN(G220) );
  NOR2_X1 U922 ( .A1(n828), .A2(n827), .ZN(G325) );
  INV_X1 U923 ( .A(G325), .ZN(G261) );
  INV_X1 U924 ( .A(n829), .ZN(G319) );
  XOR2_X1 U925 ( .A(G2096), .B(G2100), .Z(n831) );
  XNOR2_X1 U926 ( .A(KEYINPUT42), .B(G2678), .ZN(n830) );
  XNOR2_X1 U927 ( .A(n831), .B(n830), .ZN(n835) );
  XOR2_X1 U928 ( .A(KEYINPUT43), .B(G2090), .Z(n833) );
  XNOR2_X1 U929 ( .A(G2067), .B(G2072), .ZN(n832) );
  XNOR2_X1 U930 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U931 ( .A(n835), .B(n834), .Z(n837) );
  XNOR2_X1 U932 ( .A(G2084), .B(G2078), .ZN(n836) );
  XNOR2_X1 U933 ( .A(n837), .B(n836), .ZN(G227) );
  XOR2_X1 U934 ( .A(G1976), .B(G1961), .Z(n839) );
  XNOR2_X1 U935 ( .A(G1986), .B(G1966), .ZN(n838) );
  XNOR2_X1 U936 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U937 ( .A(n840), .B(KEYINPUT41), .Z(n842) );
  XNOR2_X1 U938 ( .A(G1956), .B(G1971), .ZN(n841) );
  XNOR2_X1 U939 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U940 ( .A(G2474), .B(G1981), .Z(n844) );
  XNOR2_X1 U941 ( .A(G1996), .B(G1991), .ZN(n843) );
  XNOR2_X1 U942 ( .A(n844), .B(n843), .ZN(n845) );
  XNOR2_X1 U943 ( .A(n846), .B(n845), .ZN(G229) );
  NAND2_X1 U944 ( .A1(n871), .A2(G124), .ZN(n847) );
  XNOR2_X1 U945 ( .A(n847), .B(KEYINPUT44), .ZN(n849) );
  NAND2_X1 U946 ( .A1(G112), .A2(n872), .ZN(n848) );
  NAND2_X1 U947 ( .A1(n849), .A2(n848), .ZN(n853) );
  NAND2_X1 U948 ( .A1(G136), .A2(n875), .ZN(n851) );
  NAND2_X1 U949 ( .A1(G100), .A2(n876), .ZN(n850) );
  NAND2_X1 U950 ( .A1(n851), .A2(n850), .ZN(n852) );
  NOR2_X1 U951 ( .A1(n853), .A2(n852), .ZN(G162) );
  XNOR2_X1 U952 ( .A(n854), .B(G162), .ZN(n857) );
  XOR2_X1 U953 ( .A(G160), .B(n855), .Z(n856) );
  XNOR2_X1 U954 ( .A(n857), .B(n856), .ZN(n858) );
  XNOR2_X1 U955 ( .A(n930), .B(n858), .ZN(n870) );
  NAND2_X1 U956 ( .A1(G139), .A2(n875), .ZN(n860) );
  NAND2_X1 U957 ( .A1(G103), .A2(n876), .ZN(n859) );
  NAND2_X1 U958 ( .A1(n860), .A2(n859), .ZN(n867) );
  XNOR2_X1 U959 ( .A(KEYINPUT47), .B(KEYINPUT108), .ZN(n865) );
  NAND2_X1 U960 ( .A1(n871), .A2(G127), .ZN(n863) );
  NAND2_X1 U961 ( .A1(n872), .A2(G115), .ZN(n861) );
  XOR2_X1 U962 ( .A(KEYINPUT107), .B(n861), .Z(n862) );
  NAND2_X1 U963 ( .A1(n863), .A2(n862), .ZN(n864) );
  XOR2_X1 U964 ( .A(n865), .B(n864), .Z(n866) );
  NOR2_X1 U965 ( .A1(n867), .A2(n866), .ZN(n914) );
  XNOR2_X1 U966 ( .A(n868), .B(n914), .ZN(n869) );
  XNOR2_X1 U967 ( .A(n870), .B(n869), .ZN(n888) );
  XOR2_X1 U968 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n885) );
  NAND2_X1 U969 ( .A1(G130), .A2(n871), .ZN(n874) );
  NAND2_X1 U970 ( .A1(G118), .A2(n872), .ZN(n873) );
  NAND2_X1 U971 ( .A1(n874), .A2(n873), .ZN(n882) );
  NAND2_X1 U972 ( .A1(G142), .A2(n875), .ZN(n878) );
  NAND2_X1 U973 ( .A1(G106), .A2(n876), .ZN(n877) );
  NAND2_X1 U974 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U975 ( .A(KEYINPUT45), .B(n879), .Z(n880) );
  XNOR2_X1 U976 ( .A(KEYINPUT106), .B(n880), .ZN(n881) );
  NOR2_X1 U977 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U978 ( .A(KEYINPUT109), .B(n883), .ZN(n884) );
  XNOR2_X1 U979 ( .A(n885), .B(n884), .ZN(n886) );
  XOR2_X1 U980 ( .A(G164), .B(n886), .Z(n887) );
  XNOR2_X1 U981 ( .A(n888), .B(n887), .ZN(n889) );
  NOR2_X1 U982 ( .A1(G37), .A2(n889), .ZN(G395) );
  XNOR2_X1 U983 ( .A(n977), .B(KEYINPUT110), .ZN(n893) );
  XNOR2_X1 U984 ( .A(n890), .B(G301), .ZN(n891) );
  XNOR2_X1 U985 ( .A(n891), .B(n985), .ZN(n892) );
  XNOR2_X1 U986 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U987 ( .A(G286), .B(n894), .Z(n895) );
  NOR2_X1 U988 ( .A1(G37), .A2(n895), .ZN(n896) );
  XOR2_X1 U989 ( .A(KEYINPUT111), .B(n896), .Z(G397) );
  XNOR2_X1 U990 ( .A(G2451), .B(G2427), .ZN(n906) );
  XOR2_X1 U991 ( .A(G2430), .B(G2443), .Z(n898) );
  XNOR2_X1 U992 ( .A(G2435), .B(KEYINPUT102), .ZN(n897) );
  XNOR2_X1 U993 ( .A(n898), .B(n897), .ZN(n902) );
  XOR2_X1 U994 ( .A(G2438), .B(G2454), .Z(n900) );
  XNOR2_X1 U995 ( .A(G1341), .B(G1348), .ZN(n899) );
  XNOR2_X1 U996 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U997 ( .A(n902), .B(n901), .Z(n904) );
  XNOR2_X1 U998 ( .A(G2446), .B(KEYINPUT103), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U1000 ( .A(n906), .B(n905), .ZN(n907) );
  NAND2_X1 U1001 ( .A1(n907), .A2(G14), .ZN(n913) );
  NAND2_X1 U1002 ( .A1(G319), .A2(n913), .ZN(n910) );
  NOR2_X1 U1003 ( .A1(G227), .A2(G229), .ZN(n908) );
  XNOR2_X1 U1004 ( .A(KEYINPUT49), .B(n908), .ZN(n909) );
  NOR2_X1 U1005 ( .A1(n910), .A2(n909), .ZN(n912) );
  NOR2_X1 U1006 ( .A1(G395), .A2(G397), .ZN(n911) );
  NAND2_X1 U1007 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1008 ( .A(G225), .ZN(G308) );
  INV_X1 U1009 ( .A(G69), .ZN(G235) );
  INV_X1 U1010 ( .A(n913), .ZN(G401) );
  INV_X1 U1011 ( .A(KEYINPUT55), .ZN(n942) );
  XNOR2_X1 U1012 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n940) );
  XOR2_X1 U1013 ( .A(G2072), .B(n914), .Z(n916) );
  XOR2_X1 U1014 ( .A(G164), .B(G2078), .Z(n915) );
  NOR2_X1 U1015 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1016 ( .A(KEYINPUT114), .B(n917), .ZN(n918) );
  XNOR2_X1 U1017 ( .A(n918), .B(KEYINPUT50), .ZN(n920) );
  NAND2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(n921) );
  NOR2_X1 U1019 ( .A1(n922), .A2(n921), .ZN(n937) );
  XNOR2_X1 U1020 ( .A(G2084), .B(G160), .ZN(n923) );
  XNOR2_X1 U1021 ( .A(n923), .B(KEYINPUT112), .ZN(n928) );
  XOR2_X1 U1022 ( .A(G2090), .B(G162), .Z(n924) );
  NOR2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1024 ( .A(KEYINPUT51), .B(n926), .Z(n927) );
  NAND2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n935) );
  NOR2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1027 ( .A(KEYINPUT113), .B(n931), .Z(n932) );
  NAND2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1029 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1030 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1031 ( .A(KEYINPUT52), .B(n938), .ZN(n939) );
  XNOR2_X1 U1032 ( .A(n940), .B(n939), .ZN(n941) );
  NAND2_X1 U1033 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1034 ( .A1(n943), .A2(G29), .ZN(n1025) );
  XNOR2_X1 U1035 ( .A(G2084), .B(G34), .ZN(n944) );
  XNOR2_X1 U1036 ( .A(n944), .B(KEYINPUT54), .ZN(n960) );
  XNOR2_X1 U1037 ( .A(G2090), .B(G35), .ZN(n957) );
  XOR2_X1 U1038 ( .A(G1991), .B(G25), .Z(n945) );
  NAND2_X1 U1039 ( .A1(n945), .A2(G28), .ZN(n954) );
  XNOR2_X1 U1040 ( .A(G2067), .B(G26), .ZN(n947) );
  XNOR2_X1 U1041 ( .A(G33), .B(G2072), .ZN(n946) );
  NOR2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n952) );
  XNOR2_X1 U1043 ( .A(G1996), .B(G32), .ZN(n950) );
  XNOR2_X1 U1044 ( .A(G27), .B(n948), .ZN(n949) );
  NOR2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1048 ( .A(KEYINPUT53), .B(n955), .ZN(n956) );
  NOR2_X1 U1049 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1050 ( .A(n958), .B(KEYINPUT117), .ZN(n959) );
  NOR2_X1 U1051 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1052 ( .A(KEYINPUT55), .B(n961), .Z(n963) );
  XNOR2_X1 U1053 ( .A(G29), .B(KEYINPUT118), .ZN(n962) );
  NOR2_X1 U1054 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1055 ( .A(KEYINPUT119), .B(n964), .ZN(n965) );
  NAND2_X1 U1056 ( .A1(n965), .A2(G11), .ZN(n966) );
  XNOR2_X1 U1057 ( .A(n966), .B(KEYINPUT120), .ZN(n1023) );
  XNOR2_X1 U1058 ( .A(G16), .B(KEYINPUT56), .ZN(n991) );
  XNOR2_X1 U1059 ( .A(G1966), .B(G168), .ZN(n968) );
  NAND2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1061 ( .A(n969), .B(KEYINPUT57), .ZN(n989) );
  XNOR2_X1 U1062 ( .A(n970), .B(G1956), .ZN(n972) );
  NAND2_X1 U1063 ( .A1(n972), .A2(n971), .ZN(n976) );
  XNOR2_X1 U1064 ( .A(G171), .B(G1961), .ZN(n974) );
  NAND2_X1 U1065 ( .A1(n974), .A2(n973), .ZN(n975) );
  NOR2_X1 U1066 ( .A1(n976), .A2(n975), .ZN(n983) );
  XNOR2_X1 U1067 ( .A(n977), .B(G1348), .ZN(n979) );
  NAND2_X1 U1068 ( .A1(G1971), .A2(G303), .ZN(n978) );
  NAND2_X1 U1069 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1070 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1071 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1072 ( .A(KEYINPUT121), .B(n984), .Z(n987) );
  XNOR2_X1 U1073 ( .A(G1341), .B(n985), .ZN(n986) );
  NOR2_X1 U1074 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1075 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1076 ( .A1(n991), .A2(n990), .ZN(n1021) );
  INV_X1 U1077 ( .A(G16), .ZN(n1019) );
  XOR2_X1 U1078 ( .A(G1986), .B(G24), .Z(n995) );
  XNOR2_X1 U1079 ( .A(G1971), .B(G22), .ZN(n993) );
  XNOR2_X1 U1080 ( .A(G23), .B(G1976), .ZN(n992) );
  NOR2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1082 ( .A1(n995), .A2(n994), .ZN(n997) );
  XNOR2_X1 U1083 ( .A(KEYINPUT58), .B(KEYINPUT127), .ZN(n996) );
  XNOR2_X1 U1084 ( .A(n997), .B(n996), .ZN(n1001) );
  XNOR2_X1 U1085 ( .A(G1966), .B(G21), .ZN(n999) );
  XNOR2_X1 U1086 ( .A(G5), .B(G1961), .ZN(n998) );
  NOR2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1088 ( .A1(n1001), .A2(n1000), .ZN(n1016) );
  XOR2_X1 U1089 ( .A(KEYINPUT126), .B(G4), .Z(n1003) );
  XNOR2_X1 U1090 ( .A(G1348), .B(KEYINPUT59), .ZN(n1002) );
  XNOR2_X1 U1091 ( .A(n1003), .B(n1002), .ZN(n1013) );
  XNOR2_X1 U1092 ( .A(G1956), .B(KEYINPUT122), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(n1004), .B(G20), .ZN(n1010) );
  XOR2_X1 U1094 ( .A(G1981), .B(G6), .Z(n1005) );
  XNOR2_X1 U1095 ( .A(KEYINPUT123), .B(n1005), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(G19), .B(G1341), .ZN(n1006) );
  NOR2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1098 ( .A(KEYINPUT124), .B(n1008), .Z(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(n1011), .B(KEYINPUT125), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1102 ( .A(KEYINPUT60), .B(n1014), .Z(n1015) );
  NOR2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1104 ( .A(KEYINPUT61), .B(n1017), .ZN(n1018) );
  NAND2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1108 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1026), .Z(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

