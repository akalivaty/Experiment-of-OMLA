

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586;

  XNOR2_X1 U325 ( .A(n343), .B(n342), .ZN(n370) );
  XNOR2_X1 U326 ( .A(n341), .B(n340), .ZN(n343) );
  XNOR2_X1 U327 ( .A(KEYINPUT120), .B(n493), .ZN(n293) );
  NOR2_X1 U328 ( .A1(n383), .A2(n382), .ZN(n384) );
  INV_X1 U329 ( .A(G57GAT), .ZN(n340) );
  INV_X1 U330 ( .A(n529), .ZN(n411) );
  INV_X1 U331 ( .A(n406), .ZN(n374) );
  NAND2_X1 U332 ( .A1(n411), .A2(n293), .ZN(n412) );
  XNOR2_X1 U333 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U334 ( .A(n377), .B(n376), .ZN(n380) );
  XNOR2_X1 U335 ( .A(n431), .B(n430), .ZN(n449) );
  INV_X1 U336 ( .A(G190GAT), .ZN(n450) );
  XOR2_X1 U337 ( .A(n574), .B(KEYINPUT41), .Z(n560) );
  XNOR2_X1 U338 ( .A(n450), .B(KEYINPUT58), .ZN(n451) );
  XNOR2_X1 U339 ( .A(n452), .B(n451), .ZN(G1351GAT) );
  XOR2_X1 U340 ( .A(KEYINPUT9), .B(KEYINPUT77), .Z(n295) );
  XNOR2_X1 U341 ( .A(G92GAT), .B(KEYINPUT78), .ZN(n294) );
  XNOR2_X1 U342 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U343 ( .A(n296), .B(G106GAT), .Z(n298) );
  XOR2_X1 U344 ( .A(G43GAT), .B(G134GAT), .Z(n437) );
  XNOR2_X1 U345 ( .A(n437), .B(G218GAT), .ZN(n297) );
  XNOR2_X1 U346 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U347 ( .A(G36GAT), .B(G190GAT), .Z(n401) );
  XOR2_X1 U348 ( .A(n299), .B(n401), .Z(n302) );
  XNOR2_X1 U349 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n300) );
  XNOR2_X1 U350 ( .A(n300), .B(KEYINPUT7), .ZN(n357) );
  XOR2_X1 U351 ( .A(G50GAT), .B(G162GAT), .Z(n426) );
  XNOR2_X1 U352 ( .A(n357), .B(n426), .ZN(n301) );
  XNOR2_X1 U353 ( .A(n302), .B(n301), .ZN(n311) );
  XOR2_X1 U354 ( .A(KEYINPUT76), .B(KEYINPUT11), .Z(n304) );
  XNOR2_X1 U355 ( .A(KEYINPUT79), .B(KEYINPUT65), .ZN(n303) );
  XNOR2_X1 U356 ( .A(n304), .B(n303), .ZN(n309) );
  XNOR2_X1 U357 ( .A(G99GAT), .B(G85GAT), .ZN(n305) );
  XNOR2_X1 U358 ( .A(n305), .B(KEYINPUT73), .ZN(n378) );
  XOR2_X1 U359 ( .A(KEYINPUT10), .B(n378), .Z(n307) );
  NAND2_X1 U360 ( .A1(G232GAT), .A2(G233GAT), .ZN(n306) );
  XNOR2_X1 U361 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U362 ( .A(n309), .B(n308), .Z(n310) );
  XNOR2_X1 U363 ( .A(n311), .B(n310), .ZN(n556) );
  XOR2_X1 U364 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n313) );
  XNOR2_X1 U365 ( .A(KEYINPUT5), .B(KEYINPUT90), .ZN(n312) );
  XNOR2_X1 U366 ( .A(n313), .B(n312), .ZN(n321) );
  XNOR2_X1 U367 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n314) );
  XNOR2_X1 U368 ( .A(n314), .B(G120GAT), .ZN(n441) );
  XNOR2_X1 U369 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n315) );
  XNOR2_X1 U370 ( .A(n315), .B(KEYINPUT2), .ZN(n414) );
  XNOR2_X1 U371 ( .A(n441), .B(n414), .ZN(n319) );
  XOR2_X1 U372 ( .A(KEYINPUT1), .B(G57GAT), .Z(n317) );
  XNOR2_X1 U373 ( .A(G1GAT), .B(G127GAT), .ZN(n316) );
  XNOR2_X1 U374 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U375 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U376 ( .A(n321), .B(n320), .ZN(n329) );
  NAND2_X1 U377 ( .A1(G225GAT), .A2(G233GAT), .ZN(n327) );
  XOR2_X1 U378 ( .A(G155GAT), .B(G148GAT), .Z(n323) );
  XNOR2_X1 U379 ( .A(G29GAT), .B(G134GAT), .ZN(n322) );
  XNOR2_X1 U380 ( .A(n323), .B(n322), .ZN(n325) );
  XOR2_X1 U381 ( .A(G162GAT), .B(G85GAT), .Z(n324) );
  XNOR2_X1 U382 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U383 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U384 ( .A(n329), .B(n328), .ZN(n527) );
  XNOR2_X1 U385 ( .A(KEYINPUT111), .B(KEYINPUT48), .ZN(n392) );
  XNOR2_X1 U386 ( .A(G8GAT), .B(G183GAT), .ZN(n330) );
  XNOR2_X1 U387 ( .A(n330), .B(G211GAT), .ZN(n402) );
  XOR2_X1 U388 ( .A(KEYINPUT81), .B(KEYINPUT14), .Z(n332) );
  XNOR2_X1 U389 ( .A(G1GAT), .B(G64GAT), .ZN(n331) );
  XNOR2_X1 U390 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U391 ( .A(n402), .B(n333), .Z(n335) );
  XOR2_X1 U392 ( .A(G15GAT), .B(G127GAT), .Z(n436) );
  XOR2_X1 U393 ( .A(G22GAT), .B(G155GAT), .Z(n420) );
  XNOR2_X1 U394 ( .A(n436), .B(n420), .ZN(n334) );
  XNOR2_X1 U395 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U396 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n337) );
  NAND2_X1 U397 ( .A1(G231GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U398 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U399 ( .A(n339), .B(n338), .Z(n345) );
  XNOR2_X1 U400 ( .A(G71GAT), .B(G78GAT), .ZN(n341) );
  XOR2_X1 U401 ( .A(KEYINPUT72), .B(KEYINPUT13), .Z(n342) );
  XNOR2_X1 U402 ( .A(n370), .B(KEYINPUT80), .ZN(n344) );
  XNOR2_X1 U403 ( .A(n345), .B(n344), .ZN(n468) );
  XNOR2_X1 U404 ( .A(n468), .B(KEYINPUT109), .ZN(n565) );
  NAND2_X1 U405 ( .A1(n556), .A2(n565), .ZN(n383) );
  XOR2_X1 U406 ( .A(G15GAT), .B(G141GAT), .Z(n347) );
  XNOR2_X1 U407 ( .A(G169GAT), .B(G22GAT), .ZN(n346) );
  XNOR2_X1 U408 ( .A(n347), .B(n346), .ZN(n351) );
  XOR2_X1 U409 ( .A(KEYINPUT29), .B(KEYINPUT71), .Z(n349) );
  XNOR2_X1 U410 ( .A(G113GAT), .B(G8GAT), .ZN(n348) );
  XNOR2_X1 U411 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U412 ( .A(n351), .B(n350), .Z(n356) );
  XOR2_X1 U413 ( .A(G1GAT), .B(KEYINPUT70), .Z(n353) );
  NAND2_X1 U414 ( .A1(G229GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U415 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U416 ( .A(KEYINPUT66), .B(n354), .ZN(n355) );
  XNOR2_X1 U417 ( .A(n356), .B(n355), .ZN(n361) );
  XOR2_X1 U418 ( .A(G36GAT), .B(G50GAT), .Z(n359) );
  XNOR2_X1 U419 ( .A(n357), .B(G197GAT), .ZN(n358) );
  XNOR2_X1 U420 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U421 ( .A(n361), .B(n360), .Z(n366) );
  XOR2_X1 U422 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n363) );
  XNOR2_X1 U423 ( .A(KEYINPUT69), .B(KEYINPUT68), .ZN(n362) );
  XNOR2_X1 U424 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U425 ( .A(n364), .B(G43GAT), .ZN(n365) );
  XNOR2_X1 U426 ( .A(n366), .B(n365), .ZN(n569) );
  XOR2_X1 U427 ( .A(KEYINPUT31), .B(G204GAT), .Z(n368) );
  XNOR2_X1 U428 ( .A(G176GAT), .B(G120GAT), .ZN(n367) );
  XNOR2_X1 U429 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U430 ( .A(n370), .B(n369), .ZN(n377) );
  XOR2_X1 U431 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n372) );
  NAND2_X1 U432 ( .A1(G230GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U433 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U434 ( .A(n373), .B(KEYINPUT74), .Z(n375) );
  XOR2_X1 U435 ( .A(G92GAT), .B(G64GAT), .Z(n406) );
  XOR2_X1 U436 ( .A(G106GAT), .B(G148GAT), .Z(n421) );
  XNOR2_X1 U437 ( .A(n421), .B(n378), .ZN(n379) );
  XNOR2_X1 U438 ( .A(n380), .B(n379), .ZN(n574) );
  NOR2_X1 U439 ( .A1(n569), .A2(n560), .ZN(n381) );
  XNOR2_X1 U440 ( .A(n381), .B(KEYINPUT46), .ZN(n382) );
  XNOR2_X1 U441 ( .A(n384), .B(KEYINPUT47), .ZN(n390) );
  XNOR2_X1 U442 ( .A(KEYINPUT36), .B(n556), .ZN(n584) );
  INV_X1 U443 ( .A(n468), .ZN(n578) );
  NOR2_X1 U444 ( .A1(n584), .A2(n578), .ZN(n385) );
  XNOR2_X1 U445 ( .A(KEYINPUT45), .B(n385), .ZN(n386) );
  NAND2_X1 U446 ( .A1(n386), .A2(n574), .ZN(n387) );
  XOR2_X1 U447 ( .A(KEYINPUT110), .B(n387), .Z(n388) );
  NAND2_X1 U448 ( .A1(n388), .A2(n569), .ZN(n389) );
  NAND2_X1 U449 ( .A1(n390), .A2(n389), .ZN(n391) );
  XNOR2_X1 U450 ( .A(n392), .B(n391), .ZN(n529) );
  XOR2_X1 U451 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n394) );
  XNOR2_X1 U452 ( .A(KEYINPUT18), .B(G176GAT), .ZN(n393) );
  XNOR2_X1 U453 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U454 ( .A(G169GAT), .B(n395), .Z(n435) );
  XOR2_X1 U455 ( .A(KEYINPUT87), .B(KEYINPUT86), .Z(n397) );
  XNOR2_X1 U456 ( .A(G218GAT), .B(KEYINPUT21), .ZN(n396) );
  XNOR2_X1 U457 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U458 ( .A(n398), .B(KEYINPUT88), .Z(n400) );
  XNOR2_X1 U459 ( .A(G197GAT), .B(G204GAT), .ZN(n399) );
  XNOR2_X1 U460 ( .A(n400), .B(n399), .ZN(n427) );
  XNOR2_X1 U461 ( .A(n435), .B(n427), .ZN(n410) );
  XOR2_X1 U462 ( .A(n402), .B(n401), .Z(n404) );
  NAND2_X1 U463 ( .A1(G226GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U464 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U465 ( .A(n405), .B(KEYINPUT92), .Z(n408) );
  XNOR2_X1 U466 ( .A(n406), .B(KEYINPUT91), .ZN(n407) );
  XNOR2_X1 U467 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U468 ( .A(n410), .B(n409), .ZN(n493) );
  XNOR2_X1 U469 ( .A(n412), .B(KEYINPUT54), .ZN(n413) );
  NOR2_X1 U470 ( .A1(n527), .A2(n413), .ZN(n568) );
  XOR2_X1 U471 ( .A(KEYINPUT89), .B(n414), .Z(n419) );
  XOR2_X1 U472 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n416) );
  XNOR2_X1 U473 ( .A(G211GAT), .B(G78GAT), .ZN(n415) );
  XNOR2_X1 U474 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U475 ( .A(n417), .B(KEYINPUT22), .ZN(n418) );
  XNOR2_X1 U476 ( .A(n419), .B(n418), .ZN(n425) );
  XOR2_X1 U477 ( .A(n421), .B(n420), .Z(n423) );
  NAND2_X1 U478 ( .A1(G228GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U480 ( .A(n425), .B(n424), .Z(n429) );
  XNOR2_X1 U481 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U482 ( .A(n429), .B(n428), .ZN(n462) );
  NAND2_X1 U483 ( .A1(n568), .A2(n462), .ZN(n431) );
  XOR2_X1 U484 ( .A(KEYINPUT121), .B(KEYINPUT55), .Z(n430) );
  XOR2_X1 U485 ( .A(KEYINPUT83), .B(KEYINPUT64), .Z(n433) );
  XNOR2_X1 U486 ( .A(G183GAT), .B(KEYINPUT20), .ZN(n432) );
  XNOR2_X1 U487 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U488 ( .A(n435), .B(n434), .ZN(n448) );
  XOR2_X1 U489 ( .A(G71GAT), .B(KEYINPUT82), .Z(n439) );
  XNOR2_X1 U490 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U491 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U492 ( .A(n440), .B(G190GAT), .Z(n446) );
  XOR2_X1 U493 ( .A(n441), .B(KEYINPUT84), .Z(n443) );
  NAND2_X1 U494 ( .A1(G227GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U495 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U496 ( .A(n444), .B(G99GAT), .ZN(n445) );
  XNOR2_X1 U497 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U498 ( .A(n448), .B(n447), .ZN(n531) );
  NAND2_X1 U499 ( .A1(n449), .A2(n531), .ZN(n564) );
  NOR2_X1 U500 ( .A1(n556), .A2(n564), .ZN(n452) );
  INV_X1 U501 ( .A(n527), .ZN(n517) );
  INV_X1 U502 ( .A(n569), .ZN(n503) );
  NAND2_X1 U503 ( .A1(n503), .A2(n574), .ZN(n453) );
  XNOR2_X1 U504 ( .A(n453), .B(KEYINPUT75), .ZN(n489) );
  NAND2_X1 U505 ( .A1(n531), .A2(n493), .ZN(n454) );
  NAND2_X1 U506 ( .A1(n462), .A2(n454), .ZN(n455) );
  XOR2_X1 U507 ( .A(KEYINPUT25), .B(n455), .Z(n460) );
  XNOR2_X1 U508 ( .A(KEYINPUT26), .B(KEYINPUT94), .ZN(n457) );
  NOR2_X1 U509 ( .A1(n531), .A2(n462), .ZN(n456) );
  XNOR2_X1 U510 ( .A(n457), .B(n456), .ZN(n567) );
  XOR2_X1 U511 ( .A(n493), .B(KEYINPUT27), .Z(n458) );
  XNOR2_X1 U512 ( .A(KEYINPUT93), .B(n458), .ZN(n526) );
  NAND2_X1 U513 ( .A1(n567), .A2(n526), .ZN(n459) );
  NAND2_X1 U514 ( .A1(n460), .A2(n459), .ZN(n461) );
  NOR2_X1 U515 ( .A1(n527), .A2(n461), .ZN(n467) );
  XNOR2_X1 U516 ( .A(n462), .B(KEYINPUT28), .ZN(n533) );
  NAND2_X1 U517 ( .A1(n533), .A2(n526), .ZN(n464) );
  XOR2_X1 U518 ( .A(n531), .B(KEYINPUT85), .Z(n463) );
  NOR2_X1 U519 ( .A1(n464), .A2(n463), .ZN(n465) );
  NOR2_X1 U520 ( .A1(n517), .A2(n465), .ZN(n466) );
  NOR2_X1 U521 ( .A1(n467), .A2(n466), .ZN(n484) );
  NAND2_X1 U522 ( .A1(n468), .A2(n556), .ZN(n469) );
  XOR2_X1 U523 ( .A(KEYINPUT16), .B(n469), .Z(n470) );
  AND2_X1 U524 ( .A1(n484), .A2(n470), .ZN(n504) );
  NAND2_X1 U525 ( .A1(n489), .A2(n504), .ZN(n479) );
  NOR2_X1 U526 ( .A1(n517), .A2(n479), .ZN(n472) );
  XNOR2_X1 U527 ( .A(KEYINPUT34), .B(KEYINPUT95), .ZN(n471) );
  XNOR2_X1 U528 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U529 ( .A(G1GAT), .B(n473), .ZN(G1324GAT) );
  INV_X1 U530 ( .A(n493), .ZN(n519) );
  NOR2_X1 U531 ( .A1(n519), .A2(n479), .ZN(n474) );
  XOR2_X1 U532 ( .A(G8GAT), .B(n474), .Z(G1325GAT) );
  INV_X1 U533 ( .A(n531), .ZN(n521) );
  NOR2_X1 U534 ( .A1(n479), .A2(n521), .ZN(n478) );
  XOR2_X1 U535 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n476) );
  XNOR2_X1 U536 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n475) );
  XNOR2_X1 U537 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U538 ( .A(n478), .B(n477), .ZN(G1326GAT) );
  NOR2_X1 U539 ( .A1(n533), .A2(n479), .ZN(n480) );
  XOR2_X1 U540 ( .A(KEYINPUT98), .B(n480), .Z(n481) );
  XNOR2_X1 U541 ( .A(G22GAT), .B(n481), .ZN(G1327GAT) );
  XOR2_X1 U542 ( .A(KEYINPUT99), .B(KEYINPUT102), .Z(n483) );
  XNOR2_X1 U543 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n482) );
  XNOR2_X1 U544 ( .A(n483), .B(n482), .ZN(n492) );
  NAND2_X1 U545 ( .A1(n484), .A2(n578), .ZN(n485) );
  XNOR2_X1 U546 ( .A(KEYINPUT100), .B(n485), .ZN(n486) );
  NOR2_X1 U547 ( .A1(n584), .A2(n486), .ZN(n488) );
  XNOR2_X1 U548 ( .A(KEYINPUT101), .B(KEYINPUT37), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n488), .B(n487), .ZN(n516) );
  NAND2_X1 U550 ( .A1(n516), .A2(n489), .ZN(n490) );
  XOR2_X1 U551 ( .A(KEYINPUT38), .B(n490), .Z(n500) );
  NAND2_X1 U552 ( .A1(n527), .A2(n500), .ZN(n491) );
  XOR2_X1 U553 ( .A(n492), .B(n491), .Z(G1328GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n495) );
  NAND2_X1 U555 ( .A1(n493), .A2(n500), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U557 ( .A(G36GAT), .B(n496), .ZN(G1329GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n498) );
  NAND2_X1 U559 ( .A1(n531), .A2(n500), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U561 ( .A(G43GAT), .B(n499), .ZN(G1330GAT) );
  INV_X1 U562 ( .A(n533), .ZN(n501) );
  NAND2_X1 U563 ( .A1(n501), .A2(n500), .ZN(n502) );
  XNOR2_X1 U564 ( .A(G50GAT), .B(n502), .ZN(G1331GAT) );
  NOR2_X1 U565 ( .A1(n560), .A2(n503), .ZN(n515) );
  NAND2_X1 U566 ( .A1(n515), .A2(n504), .ZN(n511) );
  NOR2_X1 U567 ( .A1(n517), .A2(n511), .ZN(n506) );
  XNOR2_X1 U568 ( .A(KEYINPUT106), .B(KEYINPUT42), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X1 U570 ( .A(G57GAT), .B(n507), .Z(G1332GAT) );
  NOR2_X1 U571 ( .A1(n519), .A2(n511), .ZN(n509) );
  XNOR2_X1 U572 ( .A(G64GAT), .B(KEYINPUT107), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n509), .B(n508), .ZN(G1333GAT) );
  NOR2_X1 U574 ( .A1(n521), .A2(n511), .ZN(n510) );
  XOR2_X1 U575 ( .A(G71GAT), .B(n510), .Z(G1334GAT) );
  NOR2_X1 U576 ( .A1(n533), .A2(n511), .ZN(n513) );
  XNOR2_X1 U577 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U579 ( .A(G78GAT), .B(n514), .ZN(G1335GAT) );
  NAND2_X1 U580 ( .A1(n516), .A2(n515), .ZN(n523) );
  NOR2_X1 U581 ( .A1(n517), .A2(n523), .ZN(n518) );
  XOR2_X1 U582 ( .A(G85GAT), .B(n518), .Z(G1336GAT) );
  NOR2_X1 U583 ( .A1(n519), .A2(n523), .ZN(n520) );
  XOR2_X1 U584 ( .A(G92GAT), .B(n520), .Z(G1337GAT) );
  NOR2_X1 U585 ( .A1(n521), .A2(n523), .ZN(n522) );
  XOR2_X1 U586 ( .A(G99GAT), .B(n522), .Z(G1338GAT) );
  NOR2_X1 U587 ( .A1(n533), .A2(n523), .ZN(n524) );
  XOR2_X1 U588 ( .A(KEYINPUT44), .B(n524), .Z(n525) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n525), .ZN(G1339GAT) );
  NAND2_X1 U590 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U591 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U592 ( .A(KEYINPUT112), .B(n530), .ZN(n546) );
  NAND2_X1 U593 ( .A1(n531), .A2(n546), .ZN(n532) );
  XNOR2_X1 U594 ( .A(n532), .B(KEYINPUT113), .ZN(n534) );
  NAND2_X1 U595 ( .A1(n534), .A2(n533), .ZN(n543) );
  NOR2_X1 U596 ( .A1(n569), .A2(n543), .ZN(n536) );
  XNOR2_X1 U597 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n535) );
  XNOR2_X1 U598 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U599 ( .A(G113GAT), .B(n537), .ZN(G1340GAT) );
  NOR2_X1 U600 ( .A1(n560), .A2(n543), .ZN(n539) );
  XNOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n538) );
  XNOR2_X1 U602 ( .A(n539), .B(n538), .ZN(G1341GAT) );
  NOR2_X1 U603 ( .A1(n565), .A2(n543), .ZN(n541) );
  XNOR2_X1 U604 ( .A(KEYINPUT50), .B(KEYINPUT116), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U606 ( .A(G127GAT), .B(n542), .Z(G1342GAT) );
  NOR2_X1 U607 ( .A1(n556), .A2(n543), .ZN(n545) );
  XNOR2_X1 U608 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n544) );
  XNOR2_X1 U609 ( .A(n545), .B(n544), .ZN(G1343GAT) );
  NAND2_X1 U610 ( .A1(n567), .A2(n546), .ZN(n555) );
  NOR2_X1 U611 ( .A1(n569), .A2(n555), .ZN(n548) );
  XNOR2_X1 U612 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(G1344GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n550) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(n552) );
  NOR2_X1 U617 ( .A1(n560), .A2(n555), .ZN(n551) );
  XOR2_X1 U618 ( .A(n552), .B(n551), .Z(G1345GAT) );
  NOR2_X1 U619 ( .A1(n578), .A2(n555), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G155GAT), .B(KEYINPUT119), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(G1346GAT) );
  NOR2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U623 ( .A(G162GAT), .B(n557), .Z(G1347GAT) );
  NOR2_X1 U624 ( .A1(n569), .A2(n564), .ZN(n558) );
  XOR2_X1 U625 ( .A(n558), .B(G169GAT), .Z(n559) );
  XNOR2_X1 U626 ( .A(KEYINPUT122), .B(n559), .ZN(G1348GAT) );
  NOR2_X1 U627 ( .A1(n564), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(G176GAT), .B(n563), .ZN(G1349GAT) );
  NOR2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U632 ( .A(G183GAT), .B(n566), .Z(G1350GAT) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n583) );
  NOR2_X1 U634 ( .A1(n569), .A2(n583), .ZN(n571) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n573) );
  XOR2_X1 U637 ( .A(KEYINPUT60), .B(KEYINPUT123), .Z(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  NOR2_X1 U639 ( .A1(n574), .A2(n583), .ZN(n576) );
  XNOR2_X1 U640 ( .A(KEYINPUT124), .B(KEYINPUT61), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G204GAT), .B(n577), .ZN(G1353GAT) );
  NOR2_X1 U643 ( .A1(n578), .A2(n583), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G211GAT), .B(KEYINPUT125), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1354GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n582) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(n586) );
  NOR2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U650 ( .A(n586), .B(n585), .Z(G1355GAT) );
endmodule

