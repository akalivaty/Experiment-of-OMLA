//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 1 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 1 0 1 0 0 0 0 0 0 1 1 0 0 1 0 1 1 1 1 1 1 0 0 1 0 1 0 1 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1328, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1400, new_n1401,
    new_n1402, new_n1403, new_n1404, new_n1405, new_n1406, new_n1407;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G58), .B2(G232), .ZN(new_n212));
  NAND4_X1  g0012(.A1(new_n209), .A2(new_n210), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n208), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT1), .ZN(new_n215));
  XNOR2_X1  g0015(.A(KEYINPUT65), .B(G20), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(G50), .B1(G58), .B2(G68), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n208), .A2(G13), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n222), .B(G250), .C1(G257), .C2(G264), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT0), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n221), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  AOI211_X1 g0025(.A(new_n215), .B(new_n225), .C1(new_n224), .C2(new_n223), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT2), .B(G226), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(G264), .B(G270), .Z(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n230), .B(new_n233), .ZN(G358));
  XNOR2_X1  g0034(.A(G87), .B(G97), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT66), .ZN(new_n236));
  XOR2_X1   g0036(.A(G107), .B(G116), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  INV_X1    g0042(.A(KEYINPUT3), .ZN(new_n243));
  INV_X1    g0043(.A(G33), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g0045(.A1(KEYINPUT3), .A2(G33), .ZN(new_n246));
  AOI21_X1  g0046(.A(G1698), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G222), .ZN(new_n248));
  INV_X1    g0048(.A(G77), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n245), .A2(new_n246), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G1698), .ZN(new_n251));
  XOR2_X1   g0051(.A(KEYINPUT68), .B(G223), .Z(new_n252));
  OAI221_X1 g0052(.A(new_n248), .B1(new_n249), .B2(new_n250), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  AND2_X1   g0053(.A1(G1), .A2(G13), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT67), .B(G1), .ZN(new_n259));
  INV_X1    g0059(.A(G41), .ZN(new_n260));
  INV_X1    g0060(.A(G45), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n259), .A2(new_n262), .B1(new_n254), .B2(new_n255), .ZN(new_n263));
  INV_X1    g0063(.A(G274), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n264), .B1(new_n254), .B2(new_n255), .ZN(new_n265));
  AOI21_X1  g0065(.A(G1), .B1(new_n260), .B2(new_n261), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n263), .A2(G226), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  AND2_X1   g0067(.A1(new_n258), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G190), .ZN(new_n269));
  INV_X1    g0069(.A(G200), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n269), .B(KEYINPUT72), .C1(new_n270), .C2(new_n268), .ZN(new_n271));
  NAND3_X1  g0071(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n217), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(KEYINPUT8), .A2(G58), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT69), .B(G58), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n275), .B1(new_n276), .B2(KEYINPUT8), .ZN(new_n277));
  INV_X1    g0077(.A(G20), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT65), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT65), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G20), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(new_n244), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n277), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G50), .A2(G58), .ZN(new_n285));
  INV_X1    g0085(.A(G68), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n278), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OR3_X1    g0087(.A1(KEYINPUT70), .A2(G20), .A3(G33), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT70), .B1(G20), .B2(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n287), .B1(new_n290), .B2(G150), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n274), .B1(new_n284), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n273), .B1(new_n259), .B2(G20), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G50), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n259), .A2(G13), .A3(G20), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n294), .B1(G50), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n297), .B(KEYINPUT9), .ZN(new_n298));
  OR3_X1    g0098(.A1(new_n271), .A2(KEYINPUT10), .A3(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(KEYINPUT10), .B1(new_n271), .B2(new_n298), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n258), .A2(new_n267), .ZN(new_n302));
  INV_X1    g0102(.A(G169), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n297), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n304), .B1(G179), .B2(new_n302), .ZN(new_n305));
  AND2_X1   g0105(.A1(KEYINPUT3), .A2(G33), .ZN(new_n306));
  NOR2_X1   g0106(.A1(KEYINPUT3), .A2(G33), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n247), .A2(G232), .B1(new_n308), .B2(G107), .ZN(new_n309));
  INV_X1    g0109(.A(G238), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n309), .B1(new_n310), .B2(new_n251), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n257), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n263), .A2(G244), .B1(new_n265), .B2(new_n266), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G200), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n293), .A2(G77), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n316), .B1(G77), .B2(new_n295), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT15), .B(G87), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n283), .A2(KEYINPUT71), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT71), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n216), .A2(G33), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n321), .B1(new_n322), .B2(new_n318), .ZN(new_n323));
  XOR2_X1   g0123(.A(KEYINPUT8), .B(G58), .Z(new_n324));
  NAND2_X1  g0124(.A1(new_n290), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n282), .A2(G77), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n320), .A2(new_n323), .A3(new_n325), .A4(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n317), .B1(new_n327), .B2(new_n273), .ZN(new_n328));
  INV_X1    g0128(.A(G190), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n315), .B(new_n328), .C1(new_n329), .C2(new_n314), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n314), .A2(new_n303), .ZN(new_n331));
  INV_X1    g0131(.A(new_n328), .ZN(new_n332));
  INV_X1    g0132(.A(G179), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n312), .A2(new_n333), .A3(new_n313), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n331), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n301), .A2(new_n305), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G1), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT67), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT67), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G1), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n262), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(G232), .A3(new_n256), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT75), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n265), .A2(new_n266), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n344), .B1(new_n343), .B2(new_n345), .ZN(new_n348));
  OR2_X1    g0148(.A1(G223), .A2(G1698), .ZN(new_n349));
  INV_X1    g0149(.A(G226), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(G1698), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n349), .B(new_n351), .C1(new_n306), .C2(new_n307), .ZN(new_n352));
  NAND2_X1  g0152(.A1(G33), .A2(G87), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n256), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NOR4_X1   g0154(.A1(new_n347), .A2(new_n348), .A3(G179), .A4(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n343), .A2(new_n345), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n354), .B1(new_n356), .B2(KEYINPUT75), .ZN(new_n357));
  AOI21_X1  g0157(.A(G169), .B1(new_n357), .B2(new_n346), .ZN(new_n358));
  OAI21_X1  g0158(.A(KEYINPUT76), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n277), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n295), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(new_n360), .B2(new_n293), .ZN(new_n362));
  INV_X1    g0162(.A(G159), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n363), .B1(new_n288), .B2(new_n289), .ZN(new_n364));
  AND2_X1   g0164(.A1(KEYINPUT69), .A2(G58), .ZN(new_n365));
  NOR2_X1   g0165(.A1(KEYINPUT69), .A2(G58), .ZN(new_n366));
  OAI21_X1  g0166(.A(G68), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(G58), .B2(G68), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n364), .B1(new_n368), .B2(G20), .ZN(new_n369));
  OAI21_X1  g0169(.A(KEYINPUT7), .B1(new_n250), .B2(G20), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT7), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n308), .A2(new_n216), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n370), .A2(new_n372), .A3(G68), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n369), .A2(new_n373), .A3(KEYINPUT16), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n273), .ZN(new_n375));
  XNOR2_X1  g0175(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT7), .B1(new_n282), .B2(new_n250), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n308), .A2(new_n371), .A3(new_n278), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n378), .A2(G68), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n377), .B1(new_n369), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n362), .B1(new_n375), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n357), .A2(new_n333), .A3(new_n346), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT76), .ZN(new_n384));
  NOR3_X1   g0184(.A1(new_n347), .A2(new_n348), .A3(new_n354), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n383), .B(new_n384), .C1(new_n385), .C2(G169), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n359), .A2(new_n382), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT18), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT18), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n359), .A2(new_n386), .A3(new_n389), .A4(new_n382), .ZN(new_n390));
  AND3_X1   g0190(.A1(new_n378), .A2(G68), .A3(new_n379), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n290), .A2(G159), .ZN(new_n392));
  NOR2_X1   g0192(.A1(G58), .A2(G68), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(new_n276), .B2(G68), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n392), .B1(new_n394), .B2(new_n278), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n376), .B1(new_n391), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n396), .A2(new_n273), .A3(new_n374), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n357), .A2(new_n346), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(G200), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n357), .A2(G190), .A3(new_n346), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n397), .A2(new_n399), .A3(new_n362), .A4(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT17), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n382), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n404), .A2(KEYINPUT17), .A3(new_n400), .A4(new_n399), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n388), .A2(new_n390), .A3(new_n403), .A4(new_n405), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n263), .A2(G238), .B1(new_n265), .B2(new_n266), .ZN(new_n407));
  OAI211_X1 g0207(.A(G232), .B(G1698), .C1(new_n306), .C2(new_n307), .ZN(new_n408));
  INV_X1    g0208(.A(G1698), .ZN(new_n409));
  OAI211_X1 g0209(.A(G226), .B(new_n409), .C1(new_n306), .C2(new_n307), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G33), .A2(G97), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n408), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n257), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n407), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT73), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n407), .A2(new_n413), .A3(KEYINPUT73), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n416), .A2(KEYINPUT13), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT13), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n407), .A2(new_n413), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n418), .A2(G179), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n411), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n422), .B1(new_n247), .B2(G226), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n256), .B1(new_n423), .B2(new_n408), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n342), .A2(new_n256), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n345), .B1(new_n425), .B2(new_n310), .ZN(new_n426));
  OAI21_X1  g0226(.A(KEYINPUT13), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n420), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT14), .B1(new_n428), .B2(G169), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT14), .ZN(new_n430));
  AOI211_X1 g0230(.A(new_n430), .B(new_n303), .C1(new_n427), .C2(new_n420), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n421), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n216), .A2(G33), .A3(G77), .ZN(new_n433));
  INV_X1    g0233(.A(new_n289), .ZN(new_n434));
  NOR3_X1   g0234(.A1(KEYINPUT70), .A2(G20), .A3(G33), .ZN(new_n435));
  OAI21_X1  g0235(.A(G50), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n286), .A2(G20), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n433), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n273), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT11), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI211_X1 g0241(.A(new_n286), .B(new_n273), .C1(G20), .C2(new_n259), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n339), .A2(new_n341), .ZN(new_n443));
  INV_X1    g0243(.A(G13), .ZN(new_n444));
  NOR3_X1   g0244(.A1(new_n443), .A2(new_n444), .A3(new_n278), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT12), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n445), .A2(new_n446), .A3(new_n286), .ZN(new_n447));
  OAI21_X1  g0247(.A(KEYINPUT12), .B1(new_n295), .B2(G68), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n442), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n438), .A2(KEYINPUT11), .A3(new_n273), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n441), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n432), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n418), .A2(G190), .A3(new_n420), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n451), .B1(new_n428), .B2(G200), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n337), .A2(new_n406), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  OAI211_X1 g0258(.A(G257), .B(G1698), .C1(new_n306), .C2(new_n307), .ZN(new_n459));
  OAI211_X1 g0259(.A(G250), .B(new_n409), .C1(new_n306), .C2(new_n307), .ZN(new_n460));
  INV_X1    g0260(.A(G294), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n459), .B(new_n460), .C1(new_n244), .C2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n257), .ZN(new_n463));
  XNOR2_X1  g0263(.A(KEYINPUT5), .B(G41), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n265), .A2(new_n259), .A3(new_n464), .A4(G45), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n339), .A2(new_n341), .A3(G45), .ZN(new_n466));
  AND2_X1   g0266(.A1(KEYINPUT5), .A2(G41), .ZN(new_n467));
  NOR2_X1   g0267(.A1(KEYINPUT5), .A2(G41), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI211_X1 g0269(.A(G264), .B(new_n256), .C1(new_n466), .C2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n463), .A2(new_n465), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n303), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n463), .A2(new_n333), .A3(new_n465), .A4(new_n470), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n250), .A2(new_n216), .A3(G87), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT22), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT22), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n250), .A2(new_n216), .A3(new_n477), .A4(G87), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(KEYINPUT23), .B1(new_n278), .B2(G107), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n278), .A2(G33), .A3(G116), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT82), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT23), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n282), .A2(new_n483), .A3(new_n484), .A4(new_n203), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n203), .ZN(new_n486));
  OAI21_X1  g0286(.A(KEYINPUT82), .B1(new_n216), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n482), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n479), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT24), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT24), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n479), .A2(new_n491), .A3(new_n488), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n274), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT78), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n494), .B1(new_n443), .B2(new_n244), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n259), .A2(KEYINPUT78), .A3(G33), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n495), .A2(new_n295), .A3(new_n496), .A4(new_n274), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT25), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(new_n295), .B2(G107), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n445), .A2(KEYINPUT25), .A3(new_n203), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n498), .A2(G107), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n474), .B1(new_n493), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n492), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n491), .B1(new_n479), .B2(new_n488), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n273), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n471), .A2(new_n270), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n463), .A2(new_n329), .A3(new_n465), .A4(new_n470), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n507), .A2(new_n510), .A3(new_n502), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n504), .A2(new_n511), .ZN(new_n512));
  AND2_X1   g0312(.A1(KEYINPUT4), .A2(G244), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n409), .B(new_n513), .C1(new_n306), .C2(new_n307), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G33), .A2(G283), .ZN(new_n515));
  INV_X1    g0315(.A(G244), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n516), .B1(new_n245), .B2(new_n246), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n514), .B(new_n515), .C1(new_n517), .C2(KEYINPUT4), .ZN(new_n518));
  OAI21_X1  g0318(.A(G250), .B1(new_n306), .B2(new_n307), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n409), .B1(new_n519), .B2(KEYINPUT4), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n257), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(G257), .B(new_n256), .C1(new_n466), .C2(new_n469), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n522), .A2(new_n465), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n521), .A2(new_n523), .A3(G190), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n270), .B1(new_n521), .B2(new_n523), .ZN(new_n525));
  OAI21_X1  g0325(.A(KEYINPUT79), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n295), .A2(G97), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(new_n497), .B2(new_n202), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n378), .A2(G107), .A3(new_n379), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G97), .A2(G107), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n204), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(KEYINPUT77), .B2(KEYINPUT6), .ZN(new_n533));
  NOR2_X1   g0333(.A1(KEYINPUT77), .A2(KEYINPUT6), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n204), .A2(new_n531), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n202), .A2(KEYINPUT6), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n533), .A2(new_n282), .A3(new_n535), .A4(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n290), .A2(G77), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n530), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n529), .B1(new_n273), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n521), .A2(new_n523), .A3(G190), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT79), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n526), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n529), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n539), .A2(new_n273), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AND3_X1   g0347(.A1(new_n521), .A2(new_n523), .A3(new_n333), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(G169), .B1(new_n521), .B2(new_n523), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n547), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n544), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(G116), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n445), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n244), .A2(G97), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n216), .A2(new_n515), .A3(new_n556), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n272), .A2(new_n217), .B1(G20), .B2(new_n554), .ZN(new_n558));
  AOI21_X1  g0358(.A(KEYINPUT20), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AND3_X1   g0359(.A1(new_n557), .A2(KEYINPUT20), .A3(new_n558), .ZN(new_n560));
  OAI221_X1 g0360(.A(new_n555), .B1(new_n497), .B2(new_n554), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(G264), .B(G1698), .C1(new_n306), .C2(new_n307), .ZN(new_n562));
  OAI211_X1 g0362(.A(G257), .B(new_n409), .C1(new_n306), .C2(new_n307), .ZN(new_n563));
  INV_X1    g0363(.A(G303), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n562), .B(new_n563), .C1(new_n564), .C2(new_n250), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n257), .ZN(new_n566));
  OAI211_X1 g0366(.A(G270), .B(new_n256), .C1(new_n466), .C2(new_n469), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n566), .A2(new_n465), .A3(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n561), .A2(KEYINPUT21), .A3(G169), .A4(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n555), .B1(new_n560), .B2(new_n559), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n497), .A2(new_n554), .ZN(new_n571));
  OAI211_X1 g0371(.A(G169), .B(new_n568), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT21), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n565), .A2(new_n257), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n567), .A2(new_n465), .ZN(new_n576));
  NOR3_X1   g0376(.A1(new_n575), .A2(new_n333), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n561), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n570), .A2(new_n571), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n568), .A2(G200), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n566), .A2(G190), .A3(new_n465), .A4(new_n567), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AND4_X1   g0382(.A1(new_n569), .A2(new_n574), .A3(new_n578), .A4(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT19), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n411), .A2(new_n584), .ZN(new_n585));
  OAI22_X1  g0385(.A1(new_n282), .A2(new_n585), .B1(G87), .B2(new_n204), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n279), .A2(new_n281), .A3(G33), .A4(G97), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n584), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n250), .A2(new_n216), .A3(G68), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT81), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n274), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n586), .A2(new_n588), .A3(KEYINPUT81), .A4(new_n589), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n592), .A2(new_n593), .B1(new_n445), .B2(new_n318), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n498), .A2(G87), .ZN(new_n595));
  INV_X1    g0395(.A(new_n466), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n265), .ZN(new_n597));
  INV_X1    g0397(.A(G250), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n598), .B1(new_n254), .B2(new_n255), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT80), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n466), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n600), .B1(new_n466), .B2(new_n599), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n597), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n247), .A2(G238), .B1(G33), .B2(G116), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n517), .A2(G1698), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n256), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NOR3_X1   g0407(.A1(new_n604), .A2(new_n607), .A3(G190), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n605), .A2(new_n606), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n257), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n466), .A2(new_n599), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT80), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n612), .A2(new_n601), .B1(new_n265), .B2(new_n596), .ZN(new_n613));
  AOI21_X1  g0413(.A(G200), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n594), .B(new_n595), .C1(new_n608), .C2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n590), .A2(new_n591), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n616), .A2(new_n273), .A3(new_n593), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n498), .A2(new_n319), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n445), .A2(new_n318), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n604), .A2(new_n607), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n333), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n303), .B1(new_n604), .B2(new_n607), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n620), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n615), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n512), .A2(new_n553), .A3(new_n583), .A4(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n458), .A2(new_n626), .ZN(G372));
  NAND2_X1  g0427(.A1(new_n405), .A2(new_n403), .ZN(new_n628));
  INV_X1    g0428(.A(new_n335), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n455), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n628), .B1(new_n452), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n388), .A2(new_n390), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n301), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n633), .A2(new_n305), .ZN(new_n634));
  AND4_X1   g0434(.A1(new_n544), .A2(new_n511), .A3(new_n552), .A4(new_n615), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n572), .A2(new_n573), .B1(new_n561), .B2(new_n577), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n504), .A2(new_n636), .A3(new_n569), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n623), .A2(KEYINPUT83), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT83), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n639), .B(new_n303), .C1(new_n604), .C2(new_n607), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n638), .A2(new_n622), .A3(new_n640), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n635), .A2(new_n637), .B1(new_n620), .B2(new_n641), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n540), .A2(new_n548), .A3(new_n550), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n625), .A2(KEYINPUT26), .A3(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n620), .A2(new_n638), .A3(new_n622), .A4(new_n640), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n645), .A2(new_n643), .A3(new_n615), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT26), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n642), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n634), .B1(new_n458), .B2(new_n651), .ZN(G369));
  NOR2_X1   g0452(.A1(new_n282), .A2(new_n444), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n653), .A2(KEYINPUT84), .A3(new_n259), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT84), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n216), .A2(G13), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n655), .B1(new_n656), .B2(new_n443), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT27), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n654), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n659), .A2(G213), .A3(G343), .A4(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n493), .B2(new_n503), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n512), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n472), .A2(new_n473), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n666), .B1(new_n507), .B2(new_n502), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n663), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT85), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n663), .A2(new_n561), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n583), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n569), .A2(new_n574), .A3(new_n578), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n673), .A2(new_n561), .A3(new_n663), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n670), .B1(new_n675), .B2(G330), .ZN(new_n676));
  INV_X1    g0476(.A(G330), .ZN(new_n677));
  AOI211_X1 g0477(.A(KEYINPUT85), .B(new_n677), .C1(new_n672), .C2(new_n674), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n669), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n673), .A2(new_n504), .A3(new_n511), .A4(new_n662), .ZN(new_n680));
  OAI211_X1 g0480(.A(new_n474), .B(new_n662), .C1(new_n493), .C2(new_n503), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n679), .A2(new_n682), .ZN(G399));
  INV_X1    g0483(.A(new_n222), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(G41), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR3_X1   g0486(.A1(new_n204), .A2(G87), .A3(G116), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n686), .A2(G1), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n688), .B1(new_n220), .B2(new_n685), .ZN(new_n689));
  XOR2_X1   g0489(.A(new_n689), .B(KEYINPUT28), .Z(new_n690));
  INV_X1    g0490(.A(KEYINPUT86), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n521), .A2(new_n523), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n463), .A2(new_n470), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n577), .A2(new_n692), .A3(new_n621), .A4(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT30), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AND4_X1   g0496(.A1(new_n470), .A2(new_n610), .A3(new_n613), .A4(new_n463), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n697), .A2(KEYINPUT30), .A3(new_n577), .A4(new_n692), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n333), .B1(new_n575), .B2(new_n576), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(new_n621), .ZN(new_n700));
  AOI22_X1  g0500(.A1(new_n693), .A2(new_n465), .B1(new_n521), .B2(new_n523), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n696), .A2(new_n698), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(KEYINPUT31), .B1(new_n703), .B2(new_n663), .ZN(new_n704));
  OAI22_X1  g0504(.A1(new_n626), .A2(new_n663), .B1(new_n691), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n703), .A2(new_n663), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT31), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n703), .A2(KEYINPUT31), .A3(new_n663), .ZN(new_n709));
  AOI21_X1  g0509(.A(KEYINPUT86), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(G330), .B1(new_n705), .B2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  XOR2_X1   g0512(.A(KEYINPUT88), .B(KEYINPUT29), .Z(new_n713));
  AOI21_X1  g0513(.A(new_n663), .B1(new_n642), .B2(new_n649), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT87), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AOI211_X1 g0516(.A(KEYINPUT87), .B(new_n663), .C1(new_n642), .C2(new_n649), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n713), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n673), .A2(new_n667), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n544), .A2(new_n511), .A3(new_n552), .A4(new_n615), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n645), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n646), .A2(KEYINPUT26), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n643), .A2(new_n615), .A3(new_n624), .A4(new_n647), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n662), .B1(new_n721), .B2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT29), .ZN(new_n726));
  OR2_X1    g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n712), .B1(new_n718), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n690), .B1(new_n728), .B2(G1), .ZN(G364));
  NAND2_X1  g0529(.A1(new_n222), .A2(new_n250), .ZN(new_n730));
  XOR2_X1   g0530(.A(new_n730), .B(KEYINPUT91), .Z(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G355), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n241), .A2(new_n261), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n684), .A2(new_n250), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(G45), .B2(new_n219), .ZN(new_n735));
  OAI221_X1 g0535(.A(new_n732), .B1(G116), .B2(new_n222), .C1(new_n733), .C2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n254), .B1(new_n278), .B2(G169), .ZN(new_n737));
  XOR2_X1   g0537(.A(new_n737), .B(KEYINPUT92), .Z(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(G13), .A2(G33), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(G20), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n736), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n338), .B1(new_n653), .B2(G45), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n685), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n270), .A2(G179), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n282), .A2(new_n329), .A3(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G179), .A2(G200), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n216), .A2(G190), .A3(new_n752), .ZN(new_n753));
  AOI22_X1  g0553(.A1(new_n750), .A2(G283), .B1(new_n753), .B2(G329), .ZN(new_n754));
  XOR2_X1   g0554(.A(new_n754), .B(KEYINPUT96), .Z(new_n755));
  NAND3_X1  g0555(.A1(new_n748), .A2(G20), .A3(G190), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n250), .B1(new_n757), .B2(G303), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n216), .A2(new_n333), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G190), .A2(G200), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(G311), .ZN(new_n762));
  INV_X1    g0562(.A(G326), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n759), .A2(G190), .A3(G200), .ZN(new_n764));
  OAI221_X1 g0564(.A(new_n758), .B1(new_n761), .B2(new_n762), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n282), .B1(new_n329), .B2(new_n752), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT95), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n766), .A2(new_n767), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n765), .B1(G294), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n759), .A2(new_n329), .A3(G200), .ZN(new_n773));
  XOR2_X1   g0573(.A(KEYINPUT33), .B(G317), .Z(new_n774));
  NOR2_X1   g0574(.A1(new_n329), .A2(G200), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n759), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G322), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n773), .A2(new_n774), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT97), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n755), .A2(new_n772), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n753), .A2(G159), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT94), .ZN(new_n782));
  XOR2_X1   g0582(.A(new_n782), .B(KEYINPUT32), .Z(new_n783));
  INV_X1    g0583(.A(G87), .ZN(new_n784));
  INV_X1    g0584(.A(new_n276), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n250), .B1(new_n784), .B2(new_n756), .C1(new_n776), .C2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(G50), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n787), .A2(new_n764), .B1(new_n773), .B2(new_n286), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n749), .A2(new_n203), .ZN(new_n789));
  NOR3_X1   g0589(.A1(new_n786), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n771), .A2(G97), .ZN(new_n791));
  INV_X1    g0591(.A(new_n761), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n792), .A2(KEYINPUT93), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(KEYINPUT93), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n790), .B(new_n791), .C1(new_n249), .C2(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n780), .B1(new_n783), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(new_n739), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n744), .A2(new_n747), .A3(new_n798), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n799), .B(KEYINPUT98), .Z(new_n800));
  INV_X1    g0600(.A(new_n742), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n675), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n675), .A2(G330), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(KEYINPUT85), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n675), .A2(new_n670), .A3(G330), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n805), .A2(KEYINPUT89), .A3(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT89), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n808), .B1(new_n676), .B2(new_n678), .ZN(new_n809));
  INV_X1    g0609(.A(new_n675), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n747), .B1(new_n810), .B2(new_n677), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n807), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n812), .A2(KEYINPUT90), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(KEYINPUT90), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n803), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(G396));
  INV_X1    g0616(.A(KEYINPUT99), .ZN(new_n817));
  NOR3_X1   g0617(.A1(new_n335), .A2(new_n817), .A3(new_n662), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n817), .B1(new_n335), .B2(new_n662), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n663), .A2(new_n332), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n819), .A2(new_n820), .B1(new_n336), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n716), .B2(new_n717), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n330), .A2(new_n335), .A3(new_n821), .ZN(new_n824));
  INV_X1    g0624(.A(new_n820), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n824), .B1(new_n825), .B2(new_n818), .ZN(new_n826));
  AND4_X1   g0626(.A1(KEYINPUT26), .A2(new_n643), .A3(new_n624), .A4(new_n615), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(new_n647), .B2(new_n646), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n662), .B(new_n826), .C1(new_n828), .C2(new_n721), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n823), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n747), .B1(new_n830), .B2(new_n711), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n711), .B2(new_n830), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n308), .B1(new_n757), .B2(G50), .ZN(new_n833));
  INV_X1    g0633(.A(new_n753), .ZN(new_n834));
  INV_X1    g0634(.A(G132), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n833), .B1(new_n286), .B2(new_n749), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n764), .ZN(new_n837));
  INV_X1    g0637(.A(new_n776), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n837), .A2(G137), .B1(new_n838), .B2(G143), .ZN(new_n839));
  INV_X1    g0639(.A(G150), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n839), .B1(new_n840), .B2(new_n773), .C1(new_n795), .C2(new_n363), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n841), .B(KEYINPUT34), .Z(new_n842));
  AOI211_X1 g0642(.A(new_n836), .B(new_n842), .C1(new_n276), .C2(new_n771), .ZN(new_n843));
  INV_X1    g0643(.A(new_n795), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(G116), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n791), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n308), .B1(new_n203), .B2(new_n756), .C1(new_n749), .C2(new_n784), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n834), .A2(new_n762), .B1(new_n776), .B2(new_n461), .ZN(new_n848));
  INV_X1    g0648(.A(G283), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n849), .A2(new_n773), .B1(new_n764), .B2(new_n564), .ZN(new_n850));
  NOR4_X1   g0650(.A1(new_n846), .A2(new_n847), .A3(new_n848), .A4(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n739), .B1(new_n843), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n822), .A2(new_n740), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n739), .A2(new_n740), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n249), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n852), .A2(new_n747), .A3(new_n853), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n832), .A2(new_n856), .ZN(G384));
  AND3_X1   g0657(.A1(new_n659), .A2(G213), .A3(new_n661), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n632), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n629), .A2(new_n662), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n861), .B(KEYINPUT100), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n829), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n451), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n865), .A2(new_n662), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n407), .A2(new_n419), .A3(new_n413), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n419), .B1(new_n407), .B2(new_n413), .ZN(new_n869));
  OAI21_X1  g0669(.A(G169), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n430), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n428), .A2(KEYINPUT14), .A3(G169), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n419), .B1(new_n414), .B2(new_n415), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n868), .B1(new_n873), .B2(new_n417), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n871), .A2(new_n872), .B1(new_n874), .B2(G179), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n455), .B(new_n867), .C1(new_n875), .C2(new_n865), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT101), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n452), .A2(KEYINPUT101), .A3(new_n455), .A4(new_n867), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n453), .A2(new_n454), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n866), .B1(new_n881), .B2(new_n432), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(KEYINPUT102), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT102), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n884), .B(new_n866), .C1(new_n881), .C2(new_n432), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n880), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n864), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n377), .B1(new_n369), .B2(new_n373), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n362), .B1(new_n375), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n858), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n406), .A2(new_n892), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n359), .A2(new_n386), .A3(new_n890), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n891), .A2(new_n401), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT37), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n382), .A2(new_n858), .ZN(new_n897));
  XOR2_X1   g0697(.A(KEYINPUT103), .B(KEYINPUT37), .Z(new_n898));
  NAND4_X1  g0698(.A1(new_n387), .A2(new_n401), .A3(new_n897), .A4(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  AND3_X1   g0700(.A1(new_n893), .A2(KEYINPUT38), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT38), .B1(new_n893), .B2(new_n900), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n860), .B1(new_n888), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n452), .A2(new_n663), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(KEYINPUT39), .B1(new_n901), .B2(new_n902), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n899), .A2(KEYINPUT104), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n897), .A2(new_n401), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT104), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n909), .A2(new_n910), .A3(new_n387), .A4(new_n898), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n387), .A2(new_n401), .A3(new_n897), .ZN(new_n912));
  INV_X1    g0712(.A(new_n898), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n908), .A2(new_n911), .A3(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n897), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n406), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT38), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n406), .A2(new_n892), .B1(new_n896), .B2(new_n899), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT39), .B1(new_n921), .B2(KEYINPUT38), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n906), .B1(new_n907), .B2(new_n923), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n904), .A2(new_n924), .A3(KEYINPUT105), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT105), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n907), .A2(new_n923), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n905), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n878), .A2(new_n879), .B1(new_n883), .B2(new_n885), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(new_n829), .B2(new_n863), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n893), .A2(new_n900), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n919), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n921), .A2(KEYINPUT38), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n930), .A2(new_n934), .B1(new_n632), .B2(new_n859), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n926), .B1(new_n928), .B2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n925), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n718), .A2(new_n457), .A3(new_n727), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n634), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n937), .B(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n708), .A2(new_n709), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n504), .A2(new_n511), .A3(new_n624), .A4(new_n615), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n544), .A2(new_n552), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n569), .A2(new_n574), .A3(new_n578), .A4(new_n582), .ZN(new_n944));
  NOR4_X1   g0744(.A1(new_n942), .A2(new_n943), .A3(new_n944), .A4(new_n663), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n826), .B1(new_n941), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(KEYINPUT106), .B1(new_n929), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n920), .A2(new_n933), .ZN(new_n948));
  AND3_X1   g0748(.A1(new_n703), .A2(KEYINPUT31), .A3(new_n663), .ZN(new_n949));
  AOI21_X1  g0749(.A(KEYINPUT31), .B1(new_n703), .B2(new_n663), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AND4_X1   g0751(.A1(new_n504), .A2(new_n511), .A3(new_n624), .A4(new_n615), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n952), .A2(new_n583), .A3(new_n553), .A4(new_n662), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n822), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT106), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n887), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n947), .A2(new_n948), .A3(new_n956), .A4(KEYINPUT40), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n954), .B(new_n887), .C1(new_n901), .C2(new_n902), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT40), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n951), .A2(new_n953), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n457), .A2(new_n962), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n961), .A2(new_n963), .ZN(new_n965));
  NOR3_X1   g0765(.A1(new_n964), .A2(new_n965), .A3(new_n677), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n940), .A2(new_n967), .B1(new_n443), .B2(new_n656), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n967), .B2(new_n940), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n533), .A2(new_n535), .A3(new_n536), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT35), .ZN(new_n971));
  OAI211_X1 g0771(.A(G116), .B(new_n218), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n972), .B1(new_n971), .B2(new_n970), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n973), .B(KEYINPUT36), .Z(new_n974));
  NAND3_X1  g0774(.A1(new_n367), .A2(G77), .A3(new_n220), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(G50), .B2(new_n286), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n976), .A2(new_n444), .A3(new_n443), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n969), .A2(new_n974), .A3(new_n977), .ZN(G367));
  INV_X1    g0778(.A(new_n734), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n743), .B1(new_n222), .B2(new_n318), .C1(new_n979), .C2(new_n233), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n747), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n844), .A2(G50), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n250), .B1(new_n785), .B2(new_n756), .ZN(new_n983));
  INV_X1    g0783(.A(G137), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n834), .A2(new_n984), .B1(new_n776), .B2(new_n840), .ZN(new_n985));
  AOI211_X1 g0785(.A(new_n983), .B(new_n985), .C1(G77), .C2(new_n750), .ZN(new_n986));
  INV_X1    g0786(.A(new_n773), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G143), .A2(new_n837), .B1(new_n987), .B2(G159), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n771), .A2(G68), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n982), .A2(new_n986), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n749), .A2(new_n202), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n756), .A2(new_n554), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT46), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n991), .B(new_n993), .C1(G303), .C2(new_n838), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n994), .B1(new_n203), .B2(new_n770), .C1(new_n849), .C2(new_n795), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n250), .B1(new_n753), .B2(G317), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n996), .B1(new_n773), .B2(new_n461), .C1(new_n762), .C2(new_n764), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n990), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT47), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n738), .B1(new_n998), .B2(new_n999), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n981), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n662), .B1(new_n594), .B2(new_n595), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(KEYINPUT107), .B1(new_n1004), .B2(new_n645), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT107), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n641), .A2(new_n1006), .A3(new_n620), .A4(new_n1003), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1004), .A2(new_n645), .A3(new_n615), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1002), .B1(new_n801), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT112), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n713), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n650), .A2(new_n662), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(KEYINPUT87), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n714), .A2(new_n715), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1012), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n727), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n711), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n663), .A2(new_n547), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n525), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n542), .B1(new_n1020), .B2(new_n541), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n540), .A2(new_n543), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1019), .B(new_n552), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT110), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n643), .A2(new_n663), .ZN(new_n1025));
  AND3_X1   g0825(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1024), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n682), .B(KEYINPUT45), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(KEYINPUT110), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(KEYINPUT45), .B1(new_n1033), .B2(new_n682), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1029), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n669), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n805), .B2(new_n806), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n680), .A2(new_n681), .ZN(new_n1039));
  XOR2_X1   g0839(.A(KEYINPUT111), .B(KEYINPUT44), .Z(new_n1040));
  NAND3_X1  g0840(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1031), .A2(new_n1039), .A3(new_n1032), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1040), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1041), .A2(new_n1044), .ZN(new_n1045));
  NOR3_X1   g0845(.A1(new_n1035), .A2(new_n1037), .A3(new_n1045), .ZN(new_n1046));
  AND2_X1   g0846(.A1(new_n1041), .A2(new_n1044), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT45), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n1028), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n679), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1046), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n663), .B1(new_n636), .B2(new_n569), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n680), .B1(new_n669), .B2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n807), .A2(new_n809), .A3(new_n1054), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n680), .B1(new_n669), .B2(new_n1053), .C1(new_n676), .C2(new_n678), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1018), .B1(new_n1052), .B2(new_n1058), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n685), .B(KEYINPUT41), .Z(new_n1060));
  OAI21_X1  g0860(.A(new_n745), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1037), .A2(new_n1033), .ZN(new_n1062));
  AOI21_X1  g0862(.A(KEYINPUT43), .B1(new_n1009), .B2(KEYINPUT108), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT108), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1005), .A2(new_n1008), .A3(new_n1007), .A4(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(KEYINPUT109), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT109), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1063), .A2(new_n1068), .A3(new_n1065), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(KEYINPUT42), .B1(new_n1038), .B2(new_n680), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT42), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1033), .A2(new_n1072), .A3(new_n512), .A4(new_n1053), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n643), .B1(new_n1033), .B2(new_n667), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1071), .B(new_n1073), .C1(new_n1074), .C2(new_n663), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1009), .A2(KEYINPUT43), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1070), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1070), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1062), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n667), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n663), .B1(new_n1082), .B2(new_n552), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1076), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1084), .A2(new_n1069), .A3(new_n1067), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1062), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1085), .A2(new_n1086), .A3(new_n1077), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1080), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1011), .B1(new_n1061), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1037), .B1(new_n1035), .B2(new_n1045), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1047), .A2(new_n679), .A3(new_n1050), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n728), .B1(new_n1093), .B2(new_n1057), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1060), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n746), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NOR3_X1   g0896(.A1(new_n1096), .A2(KEYINPUT112), .A3(new_n1088), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1010), .B1(new_n1090), .B2(new_n1097), .ZN(G387));
  NAND2_X1  g0898(.A1(new_n1018), .A2(new_n1057), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1058), .A2(new_n728), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1099), .A2(new_n1100), .A3(new_n685), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n308), .B1(new_n554), .B2(new_n749), .C1(new_n834), .C2(new_n763), .ZN(new_n1102));
  INV_X1    g0902(.A(G317), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n795), .A2(new_n564), .B1(new_n1103), .B2(new_n776), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT114), .ZN(new_n1105));
  OR2_X1    g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(G311), .A2(new_n987), .B1(new_n837), .B2(G322), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT48), .ZN(new_n1110));
  OR2_X1    g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n771), .A2(G283), .B1(G294), .B2(new_n757), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1111), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  OR2_X1    g0914(.A1(new_n1114), .A2(KEYINPUT49), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(KEYINPUT49), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1102), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n308), .B(new_n991), .C1(G77), .C2(new_n757), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n360), .B2(new_n773), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n771), .A2(new_n319), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(G50), .A2(new_n838), .B1(new_n792), .B2(G68), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1120), .B(new_n1121), .C1(new_n840), .C2(new_n834), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n1119), .B(new_n1122), .C1(G159), .C2(new_n837), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n739), .B1(new_n1117), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n747), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n669), .A2(new_n801), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n324), .A2(new_n787), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT50), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n261), .B1(new_n286), .B2(new_n249), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT113), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1129), .B1(new_n687), .B2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n1130), .B2(new_n687), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n734), .B1(new_n1128), .B2(new_n1132), .C1(new_n230), .C2(new_n261), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n731), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n1133), .B1(G107), .B2(new_n222), .C1(new_n1134), .C2(new_n687), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n1125), .B(new_n1126), .C1(new_n743), .C2(new_n1135), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n1124), .A2(new_n1136), .B1(new_n1058), .B2(new_n746), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1101), .A2(new_n1137), .ZN(G393));
  NAND2_X1  g0938(.A1(new_n1052), .A2(new_n746), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1033), .A2(new_n801), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT115), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n979), .A2(new_n238), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n743), .B1(new_n202), .B2(new_n222), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n747), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n250), .B(new_n789), .C1(G283), .C2(new_n757), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n1145), .B1(new_n461), .B2(new_n761), .C1(new_n777), .C2(new_n834), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(G303), .B2(new_n987), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n554), .B2(new_n770), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n764), .A2(new_n1103), .B1(new_n776), .B2(new_n762), .ZN(new_n1149));
  XOR2_X1   g0949(.A(new_n1149), .B(KEYINPUT52), .Z(new_n1150));
  OAI22_X1  g0950(.A1(new_n764), .A2(new_n840), .B1(new_n776), .B2(new_n363), .ZN(new_n1151));
  XOR2_X1   g0951(.A(new_n1151), .B(KEYINPUT116), .Z(new_n1152));
  NOR2_X1   g0952(.A1(new_n1152), .A2(KEYINPUT51), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(KEYINPUT51), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n844), .A2(new_n324), .B1(G77), .B2(new_n771), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n308), .B1(new_n757), .B2(G68), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n753), .A2(G143), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1156), .B(new_n1157), .C1(new_n784), .C2(new_n749), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(G50), .B2(new_n987), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1154), .A2(new_n1155), .A3(new_n1159), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n1148), .A2(new_n1150), .B1(new_n1153), .B2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1144), .B1(new_n1161), .B2(new_n739), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1141), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1139), .A2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1100), .A2(new_n1093), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1165), .A2(new_n686), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1100), .A2(new_n1093), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1164), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(G390));
  AOI22_X1  g0969(.A1(new_n934), .A2(KEYINPUT39), .B1(new_n920), .B2(new_n922), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n740), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n854), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n747), .B1(new_n1172), .B2(new_n277), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n844), .A2(G97), .B1(G77), .B2(new_n771), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n308), .B1(new_n756), .B2(new_n784), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n834), .A2(new_n461), .B1(new_n776), .B2(new_n554), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n1175), .B(new_n1176), .C1(G68), .C2(new_n750), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(G107), .A2(new_n987), .B1(new_n837), .B2(G283), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1174), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n757), .A2(G150), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n308), .B1(new_n1180), .B2(KEYINPUT53), .ZN(new_n1181));
  INV_X1    g0981(.A(G128), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1181), .B1(KEYINPUT53), .B2(new_n1180), .C1(new_n1182), .C2(new_n764), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(G137), .B2(new_n987), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(KEYINPUT54), .B(G143), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n844), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n771), .A2(G159), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n776), .A2(new_n835), .B1(new_n787), .B2(new_n749), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(G125), .B2(new_n753), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1184), .A2(new_n1187), .A3(new_n1188), .A4(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1179), .A2(new_n1191), .ZN(new_n1192));
  OR2_X1    g0992(.A1(new_n1192), .A2(KEYINPUT119), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n738), .B1(new_n1192), .B2(KEYINPUT119), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1173), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1171), .A2(new_n1195), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n826), .B(new_n662), .C1(new_n721), .C2(new_n724), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n863), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n887), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1199), .A2(new_n948), .A3(new_n906), .ZN(new_n1200));
  OAI211_X1 g1000(.A(G330), .B(new_n826), .C1(new_n705), .C2(new_n710), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n887), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n905), .B1(new_n864), .B2(new_n887), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1200), .B(new_n1203), .C1(new_n927), .C2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n862), .B1(new_n714), .B2(new_n826), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n906), .B1(new_n1206), .B2(new_n929), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n905), .B1(new_n920), .B2(new_n933), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n1170), .A2(new_n1207), .B1(new_n1199), .B2(new_n1208), .ZN(new_n1209));
  OAI211_X1 g1009(.A(G330), .B(new_n826), .C1(new_n941), .C2(new_n945), .ZN(new_n1210));
  OAI21_X1  g1010(.A(KEYINPUT117), .B1(new_n1210), .B2(new_n929), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT117), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n887), .A2(new_n954), .A3(new_n1212), .A4(G330), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1211), .A2(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1205), .B1(new_n1209), .B2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1196), .B1(new_n1215), .B2(new_n745), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n457), .A2(G330), .A3(new_n962), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n938), .A2(new_n634), .A3(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1213), .B(new_n1211), .C1(new_n1202), .C2(new_n887), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(new_n864), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1198), .B1(new_n929), .B2(new_n1210), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1203), .A2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1221), .A2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1219), .A2(new_n1224), .A3(KEYINPUT118), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT118), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n1220), .A2(new_n864), .B1(new_n1203), .B2(new_n1222), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1226), .B1(new_n1227), .B2(new_n1218), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1225), .A2(new_n1228), .A3(new_n1215), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1215), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1227), .A2(new_n1218), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n686), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1216), .B1(new_n1229), .B2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(G378));
  AOI21_X1  g1034(.A(new_n677), .B1(new_n958), .B2(new_n959), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n859), .A2(new_n297), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n301), .B2(new_n305), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n305), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n1239), .B(new_n1236), .C1(new_n299), .C2(new_n300), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1238), .A2(new_n1240), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1242), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n1238), .B2(new_n1240), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1243), .A2(new_n1245), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n1235), .A2(new_n957), .A3(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1246), .B1(new_n1235), .B2(new_n957), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n925), .A2(new_n936), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1235), .A2(new_n957), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1246), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n928), .A2(new_n926), .A3(new_n935), .ZN(new_n1253));
  OAI21_X1  g1053(.A(KEYINPUT105), .B1(new_n904), .B2(new_n924), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1235), .A2(new_n957), .A3(new_n1246), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1252), .A2(new_n1253), .A3(new_n1254), .A4(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1249), .A2(new_n746), .A3(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n747), .B1(new_n1172), .B2(G50), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n787), .B1(G33), .B2(G41), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(new_n308), .B2(new_n260), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n749), .A2(new_n785), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n761), .A2(new_n318), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n1261), .B(new_n1262), .C1(G283), .C2(new_n753), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n260), .B(new_n308), .C1(new_n756), .C2(new_n249), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n776), .A2(new_n203), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n1264), .B(new_n1265), .C1(G97), .C2(new_n987), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n837), .A2(G116), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1263), .A2(new_n1266), .A3(new_n989), .A4(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT58), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1260), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  OAI22_X1  g1070(.A1(new_n761), .A2(new_n984), .B1(new_n756), .B2(new_n1185), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1271), .B1(G128), .B2(new_n838), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(G125), .A2(new_n837), .B1(new_n987), .B2(G132), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1272), .B(new_n1273), .C1(new_n840), .C2(new_n770), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(KEYINPUT59), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n750), .A2(G159), .ZN(new_n1276));
  AOI211_X1 g1076(.A(G33), .B(G41), .C1(new_n753), .C2(G124), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1275), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1274), .A2(KEYINPUT59), .ZN(new_n1279));
  OAI221_X1 g1079(.A(new_n1270), .B1(new_n1269), .B2(new_n1268), .C1(new_n1278), .C2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1258), .B1(new_n1280), .B2(new_n739), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1281), .B1(new_n1246), .B2(new_n741), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1257), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1249), .A2(new_n1256), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1219), .B1(new_n1215), .B2(new_n1227), .ZN(new_n1286));
  AOI21_X1  g1086(.A(KEYINPUT57), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1286), .A2(KEYINPUT57), .A3(new_n1256), .A4(new_n1249), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n685), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1284), .B1(new_n1287), .B2(new_n1289), .ZN(G375));
  NAND2_X1  g1090(.A1(new_n1227), .A2(new_n1218), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1225), .A2(new_n1228), .A3(new_n1095), .A4(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n929), .A2(new_n740), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n771), .A2(G50), .ZN(new_n1294));
  OAI22_X1  g1094(.A1(new_n761), .A2(new_n840), .B1(new_n776), .B2(new_n984), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1295), .B1(G128), .B2(new_n753), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n987), .A2(new_n1186), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n250), .B1(new_n756), .B2(new_n363), .ZN(new_n1298));
  AOI211_X1 g1098(.A(new_n1298), .B(new_n1261), .C1(new_n837), .C2(G132), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1294), .A2(new_n1296), .A3(new_n1297), .A4(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1120), .B1(new_n849), .B2(new_n776), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1301), .B(KEYINPUT120), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n250), .B1(new_n757), .B2(G97), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1303), .B1(new_n249), .B2(new_n749), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1304), .B1(G303), .B2(new_n753), .ZN(new_n1305));
  AOI22_X1  g1105(.A1(G116), .A2(new_n987), .B1(new_n837), .B2(G294), .ZN(new_n1306));
  OAI211_X1 g1106(.A(new_n1305), .B(new_n1306), .C1(new_n795), .C2(new_n203), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1300), .B1(new_n1302), .B2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT121), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n738), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1310), .B1(new_n1309), .B2(new_n1308), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1125), .B1(new_n286), .B2(new_n854), .ZN(new_n1312));
  AND2_X1   g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  AOI22_X1  g1113(.A1(new_n1224), .A2(new_n746), .B1(new_n1293), .B2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1292), .A2(new_n1314), .ZN(G381));
  OAI211_X1 g1115(.A(new_n1010), .B(new_n1168), .C1(new_n1090), .C2(new_n1097), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1101), .A2(new_n815), .A3(new_n1137), .ZN(new_n1317));
  NOR4_X1   g1117(.A1(new_n1316), .A2(G384), .A3(G381), .A4(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1229), .A2(new_n1232), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1216), .ZN(new_n1320));
  AND2_X1   g1120(.A1(new_n1288), .A2(new_n685), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT57), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1286), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1249), .A2(new_n1256), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1322), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1283), .B1(new_n1321), .B2(new_n1325), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1318), .A2(new_n1319), .A3(new_n1320), .A4(new_n1326), .ZN(G407));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1233), .ZN(new_n1328));
  OAI211_X1 g1128(.A(G407), .B(G213), .C1(G343), .C2(new_n1328), .ZN(G409));
  INV_X1    g1129(.A(G213), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1330), .A2(G343), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT122), .ZN(new_n1332));
  AND3_X1   g1132(.A1(new_n1257), .A2(new_n1332), .A3(new_n1282), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1332), .B1(new_n1257), .B2(new_n1282), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1286), .A2(new_n1095), .A3(new_n1256), .A4(new_n1249), .ZN(new_n1336));
  AND3_X1   g1136(.A1(new_n1319), .A2(new_n1320), .A3(new_n1336), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1331), .B1(new_n1335), .B2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(G375), .A2(G378), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1291), .A2(KEYINPUT60), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT60), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1227), .A2(new_n1341), .A3(new_n1218), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1340), .A2(new_n1342), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n685), .B1(new_n1227), .B2(new_n1218), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1343), .A2(new_n1345), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1346), .A2(G384), .A3(new_n1314), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1344), .B1(new_n1340), .B2(new_n1342), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1314), .ZN(new_n1349));
  OAI211_X1 g1149(.A(new_n832), .B(new_n856), .C1(new_n1348), .C2(new_n1349), .ZN(new_n1350));
  AND3_X1   g1150(.A1(new_n1347), .A2(new_n1350), .A3(KEYINPUT63), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1338), .A2(new_n1339), .A3(new_n1351), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT127), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1352), .A2(new_n1353), .ZN(new_n1354));
  NAND4_X1  g1154(.A1(new_n1338), .A2(new_n1339), .A3(KEYINPUT127), .A4(new_n1351), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1354), .A2(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1347), .A2(new_n1350), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1331), .A2(G2897), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1357), .A2(new_n1358), .ZN(new_n1359));
  NAND4_X1  g1159(.A1(new_n1350), .A2(new_n1347), .A3(G2897), .A4(new_n1331), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1359), .A2(new_n1360), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1361), .A2(KEYINPUT124), .ZN(new_n1362));
  INV_X1    g1162(.A(new_n1331), .ZN(new_n1363));
  INV_X1    g1163(.A(new_n1334), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1257), .A2(new_n1332), .A3(new_n1282), .ZN(new_n1365));
  NAND4_X1  g1165(.A1(new_n1364), .A2(new_n1233), .A3(new_n1336), .A4(new_n1365), .ZN(new_n1366));
  OAI211_X1 g1166(.A(new_n1363), .B(new_n1366), .C1(new_n1326), .C2(new_n1233), .ZN(new_n1367));
  INV_X1    g1167(.A(KEYINPUT124), .ZN(new_n1368));
  NAND3_X1  g1168(.A1(new_n1359), .A2(new_n1368), .A3(new_n1360), .ZN(new_n1369));
  NAND3_X1  g1169(.A1(new_n1362), .A2(new_n1367), .A3(new_n1369), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(G387), .A2(G390), .ZN(new_n1371));
  INV_X1    g1171(.A(KEYINPUT125), .ZN(new_n1372));
  INV_X1    g1172(.A(new_n1317), .ZN(new_n1373));
  AOI21_X1  g1173(.A(new_n815), .B1(new_n1101), .B2(new_n1137), .ZN(new_n1374));
  OAI21_X1  g1174(.A(new_n1372), .B1(new_n1373), .B2(new_n1374), .ZN(new_n1375));
  INV_X1    g1175(.A(new_n1374), .ZN(new_n1376));
  NAND3_X1  g1176(.A1(new_n1376), .A2(KEYINPUT125), .A3(new_n1317), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(new_n1375), .A2(new_n1377), .ZN(new_n1378));
  NAND3_X1  g1178(.A1(new_n1371), .A2(new_n1378), .A3(new_n1316), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(new_n1379), .A2(KEYINPUT126), .ZN(new_n1380));
  INV_X1    g1180(.A(KEYINPUT126), .ZN(new_n1381));
  NAND4_X1  g1181(.A1(new_n1371), .A2(new_n1378), .A3(new_n1381), .A4(new_n1316), .ZN(new_n1382));
  NAND2_X1  g1182(.A1(new_n1371), .A2(new_n1316), .ZN(new_n1383));
  NAND2_X1  g1183(.A1(new_n1376), .A2(new_n1317), .ZN(new_n1384));
  NAND2_X1  g1184(.A1(new_n1383), .A2(new_n1384), .ZN(new_n1385));
  NAND3_X1  g1185(.A1(new_n1380), .A2(new_n1382), .A3(new_n1385), .ZN(new_n1386));
  INV_X1    g1186(.A(new_n1357), .ZN(new_n1387));
  NAND3_X1  g1187(.A1(new_n1338), .A2(new_n1339), .A3(new_n1387), .ZN(new_n1388));
  XOR2_X1   g1188(.A(KEYINPUT123), .B(KEYINPUT63), .Z(new_n1389));
  AOI21_X1  g1189(.A(KEYINPUT61), .B1(new_n1388), .B2(new_n1389), .ZN(new_n1390));
  NAND4_X1  g1190(.A1(new_n1356), .A2(new_n1370), .A3(new_n1386), .A4(new_n1390), .ZN(new_n1391));
  AOI21_X1  g1191(.A(KEYINPUT61), .B1(new_n1367), .B2(new_n1361), .ZN(new_n1392));
  NAND2_X1  g1192(.A1(new_n1388), .A2(KEYINPUT62), .ZN(new_n1393));
  INV_X1    g1193(.A(KEYINPUT62), .ZN(new_n1394));
  NAND4_X1  g1194(.A1(new_n1338), .A2(new_n1339), .A3(new_n1387), .A4(new_n1394), .ZN(new_n1395));
  NAND3_X1  g1195(.A1(new_n1392), .A2(new_n1393), .A3(new_n1395), .ZN(new_n1396));
  INV_X1    g1196(.A(new_n1386), .ZN(new_n1397));
  NAND2_X1  g1197(.A1(new_n1396), .A2(new_n1397), .ZN(new_n1398));
  NAND2_X1  g1198(.A1(new_n1391), .A2(new_n1398), .ZN(G405));
  NAND2_X1  g1199(.A1(new_n1328), .A2(new_n1339), .ZN(new_n1400));
  AOI22_X1  g1200(.A1(new_n1379), .A2(KEYINPUT126), .B1(new_n1383), .B2(new_n1384), .ZN(new_n1401));
  AOI21_X1  g1201(.A(new_n1357), .B1(new_n1401), .B2(new_n1382), .ZN(new_n1402));
  AND4_X1   g1202(.A1(new_n1382), .A2(new_n1380), .A3(new_n1385), .A4(new_n1357), .ZN(new_n1403));
  OAI21_X1  g1203(.A(new_n1400), .B1(new_n1402), .B2(new_n1403), .ZN(new_n1404));
  NAND2_X1  g1204(.A1(new_n1386), .A2(new_n1387), .ZN(new_n1405));
  NAND3_X1  g1205(.A1(new_n1401), .A2(new_n1382), .A3(new_n1357), .ZN(new_n1406));
  NAND4_X1  g1206(.A1(new_n1405), .A2(new_n1406), .A3(new_n1328), .A4(new_n1339), .ZN(new_n1407));
  NAND2_X1  g1207(.A1(new_n1404), .A2(new_n1407), .ZN(G402));
endmodule


