//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 1 1 0 1 1 0 0 1 0 1 0 1 0 1 1 1 1 0 1 1 0 0 1 1 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n530, new_n531, new_n532, new_n533, new_n534, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n545, new_n546,
    new_n547, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n600, new_n601, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1155, new_n1156;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT64), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(G125), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n466), .A2(G2105), .B1(G101), .B2(new_n468), .ZN(new_n469));
  OAI211_X1 g044(.A(G137), .B(new_n467), .C1(new_n462), .C2(new_n463), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT65), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n473), .A2(KEYINPUT65), .A3(G137), .A4(new_n467), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n469), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G112), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(G2105), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n462), .A2(new_n463), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(new_n467), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT66), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n481), .A2(G2105), .ZN(new_n485));
  AOI211_X1 g060(.A(new_n480), .B(new_n484), .C1(G136), .C2(new_n485), .ZN(G162));
  OAI211_X1 g061(.A(G138), .B(new_n467), .C1(new_n462), .C2(new_n463), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n489), .A2(new_n467), .A3(G138), .ZN(new_n490));
  OAI21_X1  g065(.A(KEYINPUT67), .B1(new_n481), .B2(new_n490), .ZN(new_n491));
  AND3_X1   g066(.A1(new_n489), .A2(new_n467), .A3(G138), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT67), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n473), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n488), .A2(new_n491), .A3(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(G2105), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n498), .B1(new_n482), .B2(G126), .ZN(new_n499));
  AND3_X1   g074(.A1(new_n495), .A2(KEYINPUT68), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g075(.A(KEYINPUT68), .B1(new_n495), .B2(new_n499), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(G164));
  AND2_X1   g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G50), .ZN(new_n508));
  INV_X1    g083(.A(G88), .ZN(new_n509));
  INV_X1    g084(.A(new_n505), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT5), .B(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n508), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n513), .A2(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n510), .A2(G543), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT69), .B(G51), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n511), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n510), .A2(G89), .ZN(new_n525));
  NAND2_X1  g100(.A1(G63), .A2(G651), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n523), .A2(new_n527), .ZN(G286));
  INV_X1    g103(.A(G286), .ZN(G168));
  NOR2_X1   g104(.A1(new_n524), .A2(new_n505), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n530), .A2(G90), .B1(new_n507), .B2(G52), .ZN(new_n531));
  XOR2_X1   g106(.A(new_n531), .B(KEYINPUT70), .Z(new_n532));
  AOI22_X1  g107(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n533), .A2(new_n515), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(new_n534), .ZN(G301));
  INV_X1    g110(.A(G301), .ZN(G171));
  NAND2_X1  g111(.A1(new_n507), .A2(G43), .ZN(new_n537));
  INV_X1    g112(.A(G81), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n538), .B2(new_n512), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n515), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  NAND4_X1  g118(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND4_X1  g121(.A1(G319), .A2(G483), .A3(G661), .A4(new_n546), .ZN(new_n547));
  XOR2_X1   g122(.A(new_n547), .B(KEYINPUT71), .Z(G188));
  XOR2_X1   g123(.A(KEYINPUT72), .B(KEYINPUT9), .Z(new_n549));
  INV_X1    g124(.A(G53), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n521), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT9), .ZN(new_n552));
  OAI211_X1 g127(.A(new_n507), .B(G53), .C1(KEYINPUT72), .C2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(G78), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G65), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n524), .B2(new_n556), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n557), .A2(G651), .B1(new_n530), .B2(G91), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n554), .A2(new_n558), .ZN(G299));
  NAND2_X1  g134(.A1(new_n530), .A2(G87), .ZN(new_n560));
  OAI21_X1  g135(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n507), .A2(G49), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  OR2_X1    g138(.A1(new_n563), .A2(KEYINPUT73), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(KEYINPUT73), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(G288));
  NAND2_X1  g142(.A1(new_n507), .A2(G48), .ZN(new_n568));
  INV_X1    g143(.A(G86), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n569), .B2(new_n512), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n511), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n571), .A2(new_n515), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n570), .A2(new_n572), .ZN(G305));
  NAND2_X1  g148(.A1(G72), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G60), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n524), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT74), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n515), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n578), .B1(new_n577), .B2(new_n576), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n530), .A2(G85), .B1(new_n507), .B2(G47), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(G290));
  NAND2_X1  g156(.A1(G301), .A2(G868), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n530), .A2(G92), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n583), .B(KEYINPUT75), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT10), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n584), .A2(new_n585), .ZN(new_n587));
  NAND2_X1  g162(.A1(G79), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G66), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n524), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(G651), .B1(new_n507), .B2(G54), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n586), .A2(new_n587), .A3(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n582), .B1(new_n593), .B2(G868), .ZN(G284));
  OAI21_X1  g169(.A(new_n582), .B1(new_n593), .B2(G868), .ZN(G321));
  NAND2_X1  g170(.A1(G286), .A2(G868), .ZN(new_n596));
  INV_X1    g171(.A(G299), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(G868), .ZN(G297));
  OAI21_X1  g173(.A(new_n596), .B1(new_n597), .B2(G868), .ZN(G280));
  XNOR2_X1  g174(.A(KEYINPUT76), .B(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n593), .B1(G860), .B2(new_n600), .ZN(new_n601));
  XOR2_X1   g176(.A(new_n601), .B(KEYINPUT77), .Z(G148));
  NAND2_X1  g177(.A1(new_n593), .A2(new_n600), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G868), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(G868), .B2(new_n542), .ZN(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g181(.A1(new_n473), .A2(new_n468), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT12), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT13), .ZN(new_n609));
  INV_X1    g184(.A(G2100), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n609), .A2(new_n610), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n485), .A2(G135), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n482), .A2(G123), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n467), .A2(G111), .ZN(new_n615));
  OAI21_X1  g190(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n613), .B(new_n614), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(G2096), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n611), .A2(new_n612), .A3(new_n619), .ZN(G156));
  XNOR2_X1  g195(.A(G2427), .B(G2438), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2430), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT15), .B(G2435), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n624), .A2(KEYINPUT14), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2451), .B(G2454), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT16), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n626), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(G2443), .B(G2446), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(G1341), .B(G1348), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT78), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT79), .ZN(new_n635));
  OAI21_X1  g210(.A(G14), .B1(new_n631), .B2(new_n633), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n635), .A2(new_n636), .ZN(G401));
  INV_X1    g212(.A(KEYINPUT18), .ZN(new_n638));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  XNOR2_X1  g214(.A(G2067), .B(G2678), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(KEYINPUT17), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n639), .A2(new_n640), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n638), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT80), .B(G2100), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2072), .B(G2078), .Z(new_n647));
  AOI21_X1  g222(.A(new_n647), .B1(new_n641), .B2(KEYINPUT18), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(new_n618), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n646), .B(new_n649), .ZN(G227));
  XOR2_X1   g225(.A(G1971), .B(G1976), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT19), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1956), .B(G2474), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1961), .B(G1966), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT20), .ZN(new_n657));
  AND2_X1   g232(.A1(new_n653), .A2(new_n654), .ZN(new_n658));
  NOR3_X1   g233(.A1(new_n652), .A2(new_n655), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n659), .B1(new_n652), .B2(new_n658), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT81), .ZN(new_n662));
  XOR2_X1   g237(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1991), .B(G1996), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1981), .B(G1986), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(G229));
  MUX2_X1   g243(.A(G24), .B(G290), .S(G16), .Z(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT83), .Z(new_n670));
  NOR2_X1   g245(.A1(new_n670), .A2(G1986), .ZN(new_n671));
  NOR2_X1   g246(.A1(G25), .A2(G29), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n485), .A2(G131), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n482), .A2(G119), .ZN(new_n674));
  OR2_X1    g249(.A1(G95), .A2(G2105), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n675), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n673), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n672), .B1(new_n678), .B2(G29), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT35), .B(G1991), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT82), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n679), .B(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n671), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n670), .A2(G1986), .ZN(new_n684));
  INV_X1    g259(.A(G16), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(G23), .ZN(new_n686));
  INV_X1    g261(.A(new_n563), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n686), .B1(new_n687), .B2(new_n685), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT33), .B(G1976), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n685), .A2(G22), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT84), .Z(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(G303), .B2(G16), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT85), .Z(new_n694));
  AOI21_X1  g269(.A(new_n690), .B1(new_n694), .B2(G1971), .ZN(new_n695));
  NOR2_X1   g270(.A1(G6), .A2(G16), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n570), .A2(new_n572), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(G16), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT32), .ZN(new_n699));
  INV_X1    g274(.A(G1981), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n695), .B(new_n701), .C1(G1971), .C2(new_n694), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n683), .B(new_n684), .C1(KEYINPUT34), .C2(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT86), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(KEYINPUT34), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT36), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n473), .A2(G127), .ZN(new_n708));
  AND2_X1   g283(.A1(G115), .A2(G2104), .ZN(new_n709));
  OAI21_X1  g284(.A(G2105), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT88), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT25), .ZN(new_n714));
  NAND2_X1  g289(.A1(G103), .A2(G2104), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(G2105), .ZN(new_n716));
  NAND4_X1  g291(.A1(new_n467), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n717));
  AOI22_X1  g292(.A1(new_n485), .A2(G139), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n712), .A2(new_n713), .A3(new_n718), .ZN(new_n719));
  MUX2_X1   g294(.A(G33), .B(new_n719), .S(G29), .Z(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G2072), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT89), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n720), .A2(G2072), .ZN(new_n723));
  INV_X1    g298(.A(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G32), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n485), .A2(G141), .B1(G105), .B2(new_n468), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n482), .A2(G129), .ZN(new_n727));
  NAND3_X1  g302(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT26), .Z(new_n729));
  AND3_X1   g304(.A1(new_n726), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n725), .B1(new_n730), .B2(new_n724), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT27), .B(G1996), .Z(new_n732));
  INV_X1    g307(.A(G34), .ZN(new_n733));
  AOI21_X1  g308(.A(G29), .B1(new_n733), .B2(KEYINPUT24), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(KEYINPUT24), .B2(new_n733), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n476), .B2(new_n724), .ZN(new_n736));
  INV_X1    g311(.A(G2084), .ZN(new_n737));
  OAI22_X1  g312(.A1(new_n731), .A2(new_n732), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NOR3_X1   g313(.A1(new_n722), .A2(new_n723), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT90), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n724), .A2(G35), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G162), .B2(new_n724), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT29), .Z(new_n743));
  INV_X1    g318(.A(G2090), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT92), .ZN(new_n746));
  NOR2_X1   g321(.A1(G168), .A2(new_n685), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n685), .B2(G21), .ZN(new_n748));
  INV_X1    g323(.A(G1966), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT31), .B(G11), .Z(new_n751));
  NOR2_X1   g326(.A1(new_n617), .A2(new_n724), .ZN(new_n752));
  INV_X1    g327(.A(G28), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n753), .A2(KEYINPUT30), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT91), .Z(new_n755));
  AOI21_X1  g330(.A(G29), .B1(new_n753), .B2(KEYINPUT30), .ZN(new_n756));
  AOI211_X1 g331(.A(new_n751), .B(new_n752), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n748), .A2(new_n749), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n731), .A2(new_n732), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n750), .A2(new_n757), .A3(new_n758), .A4(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n685), .A2(G19), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n542), .B2(new_n685), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G1341), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n736), .A2(new_n737), .ZN(new_n764));
  NOR3_X1   g339(.A1(new_n760), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(G4), .A2(G16), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n593), .B2(G16), .ZN(new_n767));
  INV_X1    g342(.A(G1348), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n685), .A2(G20), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT93), .Z(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT23), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G299), .B2(G16), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1956), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n724), .A2(G27), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G164), .B2(new_n724), .ZN(new_n776));
  INV_X1    g351(.A(G2078), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n765), .A2(new_n769), .A3(new_n774), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n685), .A2(G5), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G171), .B2(new_n685), .ZN(new_n781));
  INV_X1    g356(.A(G1961), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n724), .A2(G26), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT28), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n485), .A2(G140), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n482), .A2(G128), .ZN(new_n787));
  OR2_X1    g362(.A1(G104), .A2(G2105), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n788), .B(G2104), .C1(G116), .C2(new_n467), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n786), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n785), .B1(new_n791), .B2(new_n724), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT87), .ZN(new_n793));
  INV_X1    g368(.A(G2067), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n783), .B(new_n795), .C1(new_n743), .C2(new_n744), .ZN(new_n796));
  NOR4_X1   g371(.A1(new_n740), .A2(new_n746), .A3(new_n779), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n707), .A2(new_n797), .ZN(G150));
  INV_X1    g373(.A(G150), .ZN(G311));
  NAND2_X1  g374(.A1(new_n507), .A2(G55), .ZN(new_n800));
  INV_X1    g375(.A(G93), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n800), .B1(new_n801), .B2(new_n512), .ZN(new_n802));
  AOI22_X1  g377(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n803), .A2(new_n515), .ZN(new_n804));
  OAI21_X1  g379(.A(G860), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT96), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT95), .B(KEYINPUT37), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n593), .A2(G559), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT38), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n802), .A2(new_n804), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n542), .B(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n810), .B(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n814), .A2(KEYINPUT39), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT94), .ZN(new_n816));
  AOI21_X1  g391(.A(G860), .B1(new_n814), .B2(KEYINPUT39), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n808), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT97), .Z(G145));
  XNOR2_X1  g394(.A(new_n719), .B(new_n730), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n482), .A2(G130), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n467), .A2(G118), .ZN(new_n822));
  OAI21_X1  g397(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(G142), .B2(new_n485), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(new_n608), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n820), .B(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n495), .A2(new_n499), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(new_n790), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(new_n677), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n827), .B(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n617), .B(KEYINPUT98), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(G160), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(G162), .ZN(new_n834));
  AOI21_X1  g409(.A(G37), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n834), .B2(new_n831), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT99), .ZN(new_n837));
  XNOR2_X1  g412(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(G395));
  XNOR2_X1  g414(.A(new_n603), .B(new_n812), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n592), .B(new_n597), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(KEYINPUT41), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n842), .B1(new_n843), .B2(new_n840), .ZN(new_n844));
  XNOR2_X1  g419(.A(G290), .B(G305), .ZN(new_n845));
  XNOR2_X1  g420(.A(G303), .B(new_n687), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT42), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n844), .B(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(G868), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(G868), .B2(new_n811), .ZN(G331));
  XOR2_X1   g426(.A(G331), .B(KEYINPUT101), .Z(G295));
  XNOR2_X1  g427(.A(G301), .B(G286), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n853), .A2(new_n812), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n812), .ZN(new_n855));
  AND3_X1   g430(.A1(new_n854), .A2(new_n841), .A3(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(KEYINPUT102), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(new_n854), .ZN(new_n858));
  INV_X1    g433(.A(new_n843), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n856), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n847), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OR3_X1    g437(.A1(new_n862), .A2(KEYINPUT103), .A3(G37), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT43), .ZN(new_n864));
  OAI21_X1  g439(.A(KEYINPUT103), .B1(new_n862), .B2(G37), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n860), .A2(new_n861), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n863), .A2(new_n864), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT44), .ZN(new_n868));
  AND3_X1   g443(.A1(new_n857), .A2(new_n841), .A3(new_n854), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n843), .B1(new_n854), .B2(new_n855), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n847), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(G37), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n866), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n868), .B1(new_n873), .B2(KEYINPUT43), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n867), .A2(KEYINPUT104), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(KEYINPUT104), .B1(new_n867), .B2(new_n874), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n873), .A2(KEYINPUT43), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n863), .A2(new_n865), .A3(new_n866), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n877), .B1(new_n878), .B2(KEYINPUT43), .ZN(new_n879));
  OAI22_X1  g454(.A1(new_n875), .A2(new_n876), .B1(KEYINPUT44), .B2(new_n879), .ZN(G397));
  XOR2_X1   g455(.A(KEYINPUT105), .B(G1384), .Z(new_n881));
  AOI21_X1  g456(.A(new_n881), .B1(new_n495), .B2(new_n499), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n882), .A2(KEYINPUT45), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n469), .A2(G40), .A3(new_n475), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  OR3_X1    g461(.A1(new_n886), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n887));
  OAI21_X1  g462(.A(KEYINPUT46), .B1(new_n886), .B2(G1996), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n790), .B(new_n794), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(new_n730), .ZN(new_n890));
  AOI22_X1  g465(.A1(new_n887), .A2(new_n888), .B1(new_n885), .B2(new_n890), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n891), .B(KEYINPUT47), .Z(new_n892));
  XNOR2_X1  g467(.A(new_n730), .B(G1996), .ZN(new_n893));
  AND2_X1   g468(.A1(new_n893), .A2(new_n889), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n678), .A2(new_n680), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT125), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n791), .A2(new_n794), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n886), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OR3_X1    g474(.A1(new_n886), .A2(G1986), .A3(G290), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n901), .A2(KEYINPUT48), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n678), .A2(new_n680), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n894), .A2(new_n895), .A3(new_n903), .ZN(new_n904));
  AOI22_X1  g479(.A1(new_n901), .A2(KEYINPUT48), .B1(new_n885), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n899), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n892), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(KEYINPUT126), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT124), .ZN(new_n909));
  XNOR2_X1  g484(.A(G290), .B(G1986), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n885), .B1(new_n904), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT123), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT108), .ZN(new_n913));
  INV_X1    g488(.A(G8), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n884), .B1(new_n882), .B2(KEYINPUT45), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT68), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n828), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n495), .A2(new_n499), .A3(KEYINPUT68), .ZN(new_n918));
  AOI21_X1  g493(.A(G1384), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n915), .B1(new_n919), .B2(KEYINPUT45), .ZN(new_n920));
  INV_X1    g495(.A(G1971), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT50), .ZN(new_n923));
  INV_X1    g498(.A(G1384), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n923), .B(new_n924), .C1(new_n500), .C2(new_n501), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n828), .A2(new_n924), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n884), .B1(new_n926), .B2(KEYINPUT50), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n925), .A2(new_n927), .A3(new_n744), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n914), .B1(new_n922), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(G303), .A2(G8), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n930), .B(KEYINPUT55), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n913), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n881), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n828), .A2(KEYINPUT45), .A3(new_n934), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n469), .A2(G40), .A3(new_n475), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT45), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n924), .B1(new_n500), .B2(new_n501), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n928), .B1(new_n940), .B2(G1971), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(G8), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n942), .A2(KEYINPUT108), .A3(new_n931), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n933), .A2(new_n943), .ZN(new_n944));
  AOI211_X1 g519(.A(KEYINPUT50), .B(G1384), .C1(new_n495), .C2(new_n499), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n946), .B(new_n936), .C1(new_n919), .C2(new_n923), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n922), .B1(G2090), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT106), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n922), .B(KEYINPUT106), .C1(G2090), .C2(new_n947), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n950), .A2(new_n951), .A3(G8), .A4(new_n932), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT49), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n697), .A2(new_n700), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n697), .A2(new_n700), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n953), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n956), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n958), .A2(KEYINPUT49), .A3(new_n954), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n926), .A2(new_n884), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n961), .A2(new_n914), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G1976), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n962), .B1(new_n964), .B2(new_n563), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT52), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n966), .B1(new_n566), .B2(G1976), .ZN(new_n967));
  OAI22_X1  g542(.A1(new_n960), .A2(new_n963), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n965), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT107), .B1(new_n969), .B2(new_n966), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT107), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n965), .A2(new_n971), .A3(KEYINPUT52), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n968), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n944), .A2(new_n952), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n947), .A2(new_n782), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n777), .B(new_n915), .C1(new_n919), .C2(KEYINPUT45), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT53), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI211_X1 g553(.A(KEYINPUT45), .B(new_n924), .C1(new_n500), .C2(new_n501), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n884), .B1(new_n926), .B2(new_n938), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n979), .A2(new_n980), .A3(KEYINPUT53), .A4(new_n777), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n975), .A2(new_n978), .A3(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT120), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n982), .A2(new_n983), .A3(G171), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n983), .B1(new_n982), .B2(G171), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n974), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n945), .B1(new_n939), .B2(KEYINPUT50), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n936), .A2(new_n737), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n979), .A2(new_n980), .ZN(new_n991));
  AOI22_X1  g566(.A1(new_n988), .A2(new_n990), .B1(new_n991), .B2(new_n749), .ZN(new_n992));
  NAND2_X1  g567(.A1(G286), .A2(G8), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n993), .B(KEYINPUT116), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n992), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n991), .A2(new_n749), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n990), .B(new_n946), .C1(new_n919), .C2(new_n923), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(G8), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n997), .B1(new_n1001), .B2(new_n995), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT117), .B1(new_n992), .B2(new_n914), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT117), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1000), .A2(new_n1004), .A3(G8), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n994), .A2(KEYINPUT51), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1003), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT118), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1002), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1003), .A2(new_n1005), .A3(KEYINPUT118), .A4(new_n1006), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n996), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT62), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n987), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AOI211_X1 g588(.A(KEYINPUT62), .B(new_n996), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n912), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1002), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1016), .A2(new_n1010), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n996), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT62), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1021), .A2(new_n1022), .A3(KEYINPUT123), .A4(new_n987), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1015), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT112), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n554), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n551), .A2(new_n553), .A3(KEYINPUT112), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1026), .A2(new_n558), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT57), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT113), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n597), .A2(KEYINPUT57), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1028), .A2(new_n1033), .A3(new_n1029), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1031), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT111), .ZN(new_n1036));
  AOI21_X1  g611(.A(G1384), .B1(new_n495), .B2(new_n499), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n936), .B1(new_n1037), .B2(new_n923), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1038), .B1(new_n919), .B2(new_n923), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1036), .B1(new_n1039), .B2(G1956), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n925), .A2(new_n927), .ZN(new_n1041));
  INV_X1    g616(.A(G1956), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(KEYINPUT111), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g619(.A(KEYINPUT56), .B(G2072), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n915), .B(new_n1045), .C1(new_n919), .C2(KEYINPUT45), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT114), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n939), .A2(new_n938), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1049), .A2(KEYINPUT114), .A3(new_n915), .A4(new_n1045), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1044), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1035), .B1(new_n1052), .B2(KEYINPUT115), .ZN(new_n1053));
  AOI22_X1  g628(.A1(new_n1040), .A2(new_n1043), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT115), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1044), .A2(new_n1051), .A3(new_n1035), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n947), .A2(new_n768), .ZN(new_n1058));
  INV_X1    g633(.A(new_n961), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1059), .A2(G2067), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n592), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1062));
  AOI22_X1  g637(.A1(new_n1053), .A2(new_n1056), .B1(new_n1057), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT60), .ZN(new_n1064));
  AOI21_X1  g639(.A(G1348), .B1(new_n988), .B2(new_n936), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1064), .B1(new_n1065), .B2(new_n1060), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1058), .A2(KEYINPUT60), .A3(new_n1061), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n1066), .A2(new_n1067), .A3(new_n593), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n1069));
  INV_X1    g644(.A(G1996), .ZN(new_n1070));
  XOR2_X1   g645(.A(KEYINPUT58), .B(G1341), .Z(new_n1071));
  AOI22_X1  g646(.A1(new_n940), .A2(new_n1070), .B1(new_n1059), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n542), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1069), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1058), .A2(new_n1061), .A3(KEYINPUT60), .A4(new_n592), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1059), .A2(new_n1071), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1076), .B1(new_n920), .B2(G1996), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1077), .A2(KEYINPUT59), .A3(new_n542), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1074), .A2(new_n1075), .A3(new_n1078), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1068), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT61), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1044), .A2(new_n1051), .A3(new_n1035), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1035), .B1(new_n1044), .B2(new_n1051), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1081), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1080), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1057), .A2(KEYINPUT61), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1086), .B1(new_n1053), .B2(new_n1056), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1063), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n974), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT54), .B1(new_n982), .B2(G171), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n883), .A2(new_n915), .A3(KEYINPUT53), .A4(new_n777), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n975), .A2(new_n978), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT122), .ZN(new_n1093));
  OR2_X1    g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(G301), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1090), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n985), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n975), .A2(new_n978), .A3(G301), .A4(new_n1091), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT121), .ZN(new_n1099));
  OR2_X1    g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n982), .A2(new_n983), .A3(G171), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1097), .A2(new_n1100), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  XOR2_X1   g678(.A(KEYINPUT119), .B(KEYINPUT54), .Z(new_n1104));
  AOI21_X1  g679(.A(new_n1096), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1088), .A2(new_n1089), .A3(new_n1105), .A4(new_n1020), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n950), .A2(G8), .A3(new_n951), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n931), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT63), .ZN(new_n1109));
  AOI211_X1 g684(.A(new_n945), .B(new_n989), .C1(new_n939), .C2(KEYINPUT50), .ZN(new_n1110));
  AOI21_X1  g685(.A(G1966), .B1(new_n979), .B2(new_n980), .ZN(new_n1111));
  OAI211_X1 g686(.A(G8), .B(G168), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(KEYINPUT109), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n914), .B1(new_n998), .B2(new_n999), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT109), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1114), .A2(new_n1115), .A3(G168), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1109), .B1(new_n1113), .B2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1108), .A2(new_n1117), .A3(new_n952), .A4(new_n973), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n944), .A2(new_n952), .A3(new_n1119), .A4(new_n973), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT110), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1109), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1118), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n952), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n973), .ZN(new_n1126));
  INV_X1    g701(.A(new_n960), .ZN(new_n1127));
  AOI211_X1 g702(.A(G1976), .B(G288), .C1(new_n1127), .C2(new_n962), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n962), .B1(new_n1128), .B2(new_n955), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1106), .A2(new_n1124), .A3(new_n1131), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n909), .B(new_n911), .C1(new_n1024), .C2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1081), .B1(new_n1054), .B2(new_n1035), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1035), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1136), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1052), .A2(KEYINPUT115), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1135), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1139), .A2(new_n1084), .A3(new_n1080), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1011), .B1(new_n1140), .B2(new_n1063), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1104), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n1098), .B(KEYINPUT121), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1142), .B1(new_n986), .B2(new_n1143), .ZN(new_n1144));
  NOR3_X1   g719(.A1(new_n1144), .A2(new_n974), .A3(new_n1096), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1130), .B1(new_n1141), .B2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1146), .A2(new_n1015), .A3(new_n1124), .A4(new_n1023), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n909), .B1(new_n1147), .B2(new_n911), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n908), .B1(new_n1134), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(KEYINPUT127), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT127), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n1151), .B(new_n908), .C1(new_n1134), .C2(new_n1148), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1150), .A2(new_n1152), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g728(.A1(G229), .A2(new_n460), .A3(G401), .A4(G227), .ZN(new_n1155));
  NAND2_X1  g729(.A1(new_n1155), .A2(new_n837), .ZN(new_n1156));
  NOR2_X1   g730(.A1(new_n879), .A2(new_n1156), .ZN(G308));
  INV_X1    g731(.A(G308), .ZN(G225));
endmodule


