//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 1 1 1 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 0 1 0 0 1 1 0 0 0 1 1 1 0 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n636, new_n637, new_n638,
    new_n639, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n837, new_n838, new_n839, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957;
  INV_X1    g000(.A(KEYINPUT74), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT24), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n203), .A2(G183gat), .A3(G190gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  INV_X1    g004(.A(G183gat), .ZN(new_n206));
  INV_X1    g005(.A(G190gat), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT24), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NOR2_X1   g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209));
  OAI221_X1 g008(.A(new_n204), .B1(KEYINPUT23), .B2(new_n205), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  INV_X1    g010(.A(new_n205), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT23), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n210), .B1(KEYINPUT65), .B2(new_n214), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n214), .A2(KEYINPUT65), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT25), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n217), .B1(new_n210), .B2(new_n214), .ZN(new_n219));
  AOI22_X1  g018(.A1(new_n215), .A2(new_n218), .B1(new_n219), .B2(KEYINPUT64), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(KEYINPUT64), .B2(new_n219), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT26), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n212), .A2(new_n222), .A3(new_n211), .ZN(new_n223));
  OAI221_X1 g022(.A(new_n223), .B1(new_n222), .B2(new_n212), .C1(new_n206), .C2(new_n207), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT66), .ZN(new_n225));
  OR2_X1    g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n225), .ZN(new_n227));
  XNOR2_X1  g026(.A(KEYINPUT27), .B(G183gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(new_n207), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n229), .A2(KEYINPUT28), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(KEYINPUT28), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n226), .A2(new_n227), .A3(new_n230), .A4(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n221), .A2(new_n232), .ZN(new_n233));
  AND3_X1   g032(.A1(new_n233), .A2(G226gat), .A3(G233gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT29), .ZN(new_n235));
  AOI22_X1  g034(.A1(new_n233), .A2(new_n235), .B1(G226gat), .B2(G233gat), .ZN(new_n236));
  OR2_X1    g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT73), .B(G218gat), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT22), .B1(new_n238), .B2(G211gat), .ZN(new_n239));
  XOR2_X1   g038(.A(G197gat), .B(G204gat), .Z(new_n240));
  NOR2_X1   g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G211gat), .B(G218gat), .ZN(new_n242));
  XOR2_X1   g041(.A(new_n241), .B(new_n242), .Z(new_n243));
  NAND2_X1  g042(.A1(new_n237), .A2(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n234), .A2(new_n236), .ZN(new_n245));
  INV_X1    g044(.A(new_n243), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G8gat), .B(G36gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(G64gat), .B(G92gat), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n249), .B(new_n250), .Z(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n202), .B1(new_n248), .B2(new_n252), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n244), .A2(KEYINPUT74), .A3(new_n247), .A4(new_n251), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT37), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n256), .B1(new_n244), .B2(new_n247), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n257), .A2(KEYINPUT85), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n252), .B1(new_n248), .B2(KEYINPUT37), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT38), .B1(new_n257), .B2(KEYINPUT85), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n255), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(G141gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(G148gat), .ZN(new_n264));
  INV_X1    g063(.A(G148gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G141gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G155gat), .ZN(new_n268));
  INV_X1    g067(.A(G162gat), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT2), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(G155gat), .B(G162gat), .ZN(new_n272));
  OR2_X1    g071(.A1(new_n272), .A2(KEYINPUT75), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(KEYINPUT75), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n271), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AND2_X1   g074(.A1(new_n267), .A2(new_n270), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT76), .B1(new_n276), .B2(new_n272), .ZN(new_n277));
  OR2_X1    g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT76), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT3), .ZN(new_n283));
  INV_X1    g082(.A(G113gat), .ZN(new_n284));
  INV_X1    g083(.A(G120gat), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT1), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n286), .B1(new_n284), .B2(new_n285), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G127gat), .B(G134gat), .ZN(new_n289));
  OR2_X1    g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  XOR2_X1   g089(.A(KEYINPUT67), .B(G113gat), .Z(new_n291));
  OAI211_X1 g090(.A(new_n286), .B(new_n289), .C1(new_n291), .C2(new_n285), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT3), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n281), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n283), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(G225gat), .A2(G233gat), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NOR3_X1   g098(.A1(new_n297), .A2(KEYINPUT5), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n281), .A2(new_n290), .A3(new_n292), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n301), .B(KEYINPUT4), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n302), .A2(KEYINPUT80), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT4), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n301), .B(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT80), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n300), .B1(new_n303), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n302), .A2(new_n298), .A3(new_n296), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT5), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n282), .A2(new_n293), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(new_n301), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n310), .B1(new_n312), .B2(new_n299), .ZN(new_n313));
  AND3_X1   g112(.A1(new_n309), .A2(KEYINPUT77), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(KEYINPUT77), .B1(new_n309), .B2(new_n313), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n308), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  XOR2_X1   g115(.A(G1gat), .B(G29gat), .Z(new_n317));
  XNOR2_X1  g116(.A(new_n317), .B(KEYINPUT79), .ZN(new_n318));
  XOR2_X1   g117(.A(G57gat), .B(G85gat), .Z(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n321));
  XOR2_X1   g120(.A(new_n320), .B(new_n321), .Z(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT81), .B1(new_n316), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n313), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT77), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n309), .A2(new_n313), .A3(KEYINPUT77), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT81), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n329), .A2(new_n330), .A3(new_n322), .A4(new_n308), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n323), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT6), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n324), .A2(new_n331), .A3(new_n332), .A4(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n316), .A2(KEYINPUT6), .A3(new_n323), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT38), .B1(new_n259), .B2(new_n257), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n262), .A2(new_n334), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n311), .A2(new_n298), .A3(new_n301), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n305), .A2(new_n306), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n302), .A2(KEYINPUT80), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n297), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  OAI211_X1 g140(.A(KEYINPUT39), .B(new_n338), .C1(new_n341), .C2(new_n298), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n296), .B1(new_n303), .B2(new_n307), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT39), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n343), .A2(new_n344), .A3(new_n299), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n342), .A2(new_n345), .A3(new_n322), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT40), .ZN(new_n347));
  OR2_X1    g146(.A1(new_n347), .A2(KEYINPUT84), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(KEYINPUT84), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT30), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n253), .A2(new_n352), .A3(new_n254), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n251), .B1(new_n244), .B2(new_n247), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n248), .A2(new_n252), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n354), .B1(new_n355), .B2(KEYINPUT30), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n346), .A2(KEYINPUT84), .A3(new_n347), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n351), .A2(new_n357), .A3(new_n332), .A4(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G78gat), .B(G106gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(G22gat), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n246), .B1(new_n295), .B2(new_n235), .ZN(new_n363));
  OR2_X1    g162(.A1(new_n363), .A2(KEYINPUT83), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n241), .A2(new_n242), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT82), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n242), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT29), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n368), .B1(new_n246), .B2(KEYINPUT82), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(new_n294), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(new_n282), .ZN(new_n371));
  NAND2_X1  g170(.A1(G228gat), .A2(G233gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n363), .A2(KEYINPUT83), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n364), .A2(new_n371), .A3(new_n372), .A4(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n246), .A2(new_n235), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n281), .B1(new_n375), .B2(new_n294), .ZN(new_n376));
  OAI211_X1 g175(.A(G228gat), .B(G233gat), .C1(new_n376), .C2(new_n363), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT31), .B(G50gat), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n374), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n379), .B1(new_n374), .B2(new_n377), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n362), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n382), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n384), .A2(new_n361), .A3(new_n380), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  AND3_X1   g186(.A1(new_n337), .A2(new_n359), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n357), .B1(new_n334), .B2(new_n335), .ZN(new_n389));
  XOR2_X1   g188(.A(G71gat), .B(G99gat), .Z(new_n390));
  XNOR2_X1  g189(.A(G15gat), .B(G43gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n390), .B(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n233), .B(new_n293), .ZN(new_n393));
  NAND2_X1  g192(.A1(G227gat), .A2(G233gat), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT32), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT69), .ZN(new_n398));
  XOR2_X1   g197(.A(KEYINPUT68), .B(KEYINPUT33), .Z(new_n399));
  AOI21_X1  g198(.A(new_n398), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n399), .ZN(new_n401));
  AOI211_X1 g200(.A(KEYINPUT69), .B(new_n401), .C1(new_n393), .C2(new_n395), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n392), .B(new_n397), .C1(new_n400), .C2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n392), .A2(new_n401), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n396), .A2(KEYINPUT32), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT70), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT70), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n396), .A2(new_n407), .A3(KEYINPUT32), .A4(new_n404), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n403), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n393), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT34), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n411), .A2(new_n412), .A3(new_n394), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT72), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n411), .A2(KEYINPUT72), .A3(new_n412), .A4(new_n394), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT34), .B1(new_n393), .B2(new_n395), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n410), .A2(new_n418), .ZN(new_n419));
  AND3_X1   g218(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n420), .A2(new_n409), .A3(new_n403), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT36), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT36), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n418), .A2(KEYINPUT71), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n410), .A2(new_n424), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n418), .A2(new_n403), .A3(new_n409), .A4(KEYINPUT71), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n423), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  OAI22_X1  g226(.A1(new_n389), .A2(new_n387), .B1(new_n422), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n421), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n420), .B1(new_n403), .B2(new_n409), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n386), .A2(KEYINPUT35), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n389), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT35), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n386), .B1(new_n425), .B2(new_n426), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n434), .B1(new_n389), .B2(new_n435), .ZN(new_n436));
  OAI22_X1  g235(.A1(new_n388), .A2(new_n428), .B1(new_n433), .B2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G113gat), .B(G141gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(KEYINPUT86), .B(G197gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n438), .B(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(KEYINPUT11), .B(G169gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n440), .B(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n442), .B(KEYINPUT12), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT87), .ZN(new_n444));
  INV_X1    g243(.A(G50gat), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n444), .B1(new_n445), .B2(G43gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(G43gat), .ZN(new_n447));
  INV_X1    g246(.A(G43gat), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n448), .A2(KEYINPUT87), .A3(G50gat), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n446), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT15), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT15), .B1(new_n445), .B2(G43gat), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n448), .A2(G50gat), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(G29gat), .ZN(new_n457));
  INV_X1    g256(.A(G36gat), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n457), .A2(new_n458), .A3(KEYINPUT14), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT14), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n460), .B1(G29gat), .B2(G36gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(G29gat), .A2(G36gat), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n459), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n452), .A2(new_n456), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n463), .A2(new_n455), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT88), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n463), .A2(new_n455), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n469), .A2(KEYINPUT88), .A3(new_n452), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(G15gat), .B(G22gat), .ZN(new_n472));
  INV_X1    g271(.A(G1gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT16), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n475), .B1(G1gat), .B2(new_n472), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n476), .B(G8gat), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n471), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(G229gat), .A2(G233gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT89), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n469), .A2(KEYINPUT88), .A3(new_n452), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n469), .A2(new_n452), .B1(new_n466), .B2(KEYINPUT88), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT17), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT17), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n468), .A2(new_n486), .A3(new_n470), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n477), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n482), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AOI211_X1 g289(.A(KEYINPUT89), .B(new_n477), .C1(new_n485), .C2(new_n487), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n481), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT90), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT18), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT90), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n495), .B(new_n481), .C1(new_n490), .C2(new_n491), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n493), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  OAI211_X1 g296(.A(KEYINPUT18), .B(new_n481), .C1(new_n490), .C2(new_n491), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n471), .B(new_n477), .ZN(new_n499));
  XOR2_X1   g298(.A(new_n479), .B(KEYINPUT13), .Z(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n443), .B1(new_n497), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT91), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n493), .A2(new_n504), .A3(new_n494), .A4(new_n496), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n498), .A2(new_n501), .A3(new_n443), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AND3_X1   g306(.A1(new_n468), .A2(new_n486), .A3(new_n470), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n486), .B1(new_n468), .B2(new_n470), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n489), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT89), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n488), .A2(new_n482), .A3(new_n489), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n480), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n494), .B1(new_n513), .B2(new_n495), .ZN(new_n514));
  INV_X1    g313(.A(new_n496), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT91), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n503), .B1(new_n507), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n437), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n334), .A2(new_n335), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n520), .A2(KEYINPUT96), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n520), .A2(KEYINPUT96), .ZN(new_n522));
  OR2_X1    g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(G85gat), .A2(G92gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  INV_X1    g325(.A(G99gat), .ZN(new_n527));
  INV_X1    g326(.A(G106gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(G99gat), .A2(G106gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(G85gat), .ZN(new_n532));
  INV_X1    g331(.A(G92gat), .ZN(new_n533));
  AOI22_X1  g332(.A1(KEYINPUT8), .A2(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n526), .A2(new_n531), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n531), .B1(new_n526), .B2(new_n534), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AND2_X1   g337(.A1(G232gat), .A2(G233gat), .ZN(new_n539));
  AOI22_X1  g338(.A1(new_n471), .A2(new_n538), .B1(KEYINPUT41), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n488), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n540), .B1(new_n541), .B2(new_n538), .ZN(new_n542));
  XOR2_X1   g341(.A(G190gat), .B(G218gat), .Z(new_n543));
  XOR2_X1   g342(.A(new_n542), .B(new_n543), .Z(new_n544));
  NOR2_X1   g343(.A1(new_n539), .A2(KEYINPUT41), .ZN(new_n545));
  XNOR2_X1  g344(.A(G134gat), .B(G162gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n544), .B(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(G71gat), .A2(G78gat), .ZN(new_n550));
  OR2_X1    g349(.A1(G71gat), .A2(G78gat), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT9), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT92), .ZN(new_n554));
  INV_X1    g353(.A(G57gat), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n554), .B1(new_n555), .B2(G64gat), .ZN(new_n556));
  INV_X1    g355(.A(G64gat), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n557), .A2(KEYINPUT92), .A3(G57gat), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n556), .B(new_n558), .C1(G57gat), .C2(new_n557), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n555), .A2(G64gat), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n557), .A2(G57gat), .ZN(new_n561));
  OAI21_X1  g360(.A(KEYINPUT9), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n551), .A2(new_n550), .ZN(new_n563));
  AOI22_X1  g362(.A1(new_n553), .A2(new_n559), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n564), .A2(KEYINPUT21), .ZN(new_n565));
  NAND2_X1  g364(.A1(G231gat), .A2(G233gat), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n565), .B(new_n566), .Z(new_n567));
  XNOR2_X1  g366(.A(G127gat), .B(G155gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT20), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n567), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G183gat), .B(G211gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n477), .B1(KEYINPUT21), .B2(new_n564), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  OR2_X1    g374(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n572), .A2(new_n575), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n549), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n559), .A2(new_n553), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n562), .A2(new_n563), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT94), .B1(new_n526), .B2(new_n534), .ZN(new_n583));
  OAI22_X1  g382(.A1(new_n582), .A2(new_n583), .B1(new_n536), .B2(new_n537), .ZN(new_n584));
  INV_X1    g383(.A(new_n537), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n526), .A2(new_n534), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT94), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n585), .A2(new_n564), .A3(new_n588), .A4(new_n535), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT10), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n584), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n538), .A2(KEYINPUT10), .A3(new_n564), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G230gat), .A2(G233gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n584), .A2(new_n589), .ZN(new_n596));
  INV_X1    g395(.A(new_n594), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G120gat), .B(G148gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT95), .ZN(new_n601));
  XNOR2_X1  g400(.A(G176gat), .B(G204gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n599), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n599), .A2(new_n604), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n579), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n524), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(G1gat), .ZN(G1324gat));
  INV_X1    g412(.A(new_n519), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n614), .A2(new_n611), .A3(new_n357), .ZN(new_n615));
  XOR2_X1   g414(.A(KEYINPUT16), .B(G8gat), .Z(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  AOI22_X1  g417(.A1(new_n618), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n615), .ZN(new_n619));
  INV_X1    g418(.A(new_n618), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT97), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT42), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n621), .B1(new_n620), .B2(new_n622), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n619), .B1(new_n624), .B2(new_n625), .ZN(G1325gat));
  NOR2_X1   g425(.A1(new_n427), .A2(new_n422), .ZN(new_n627));
  AND4_X1   g426(.A1(G15gat), .A2(new_n614), .A3(new_n611), .A4(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n431), .ZN(new_n629));
  NOR3_X1   g428(.A1(new_n519), .A2(new_n610), .A3(new_n629), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n630), .A2(G15gat), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT98), .ZN(new_n632));
  OR2_X1    g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n628), .B1(new_n633), .B2(new_n634), .ZN(G1326gat));
  NOR2_X1   g434(.A1(new_n519), .A2(new_n387), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n611), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT99), .ZN(new_n638));
  XNOR2_X1  g437(.A(KEYINPUT43), .B(G22gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(G1327gat));
  INV_X1    g439(.A(new_n578), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n641), .A2(new_n608), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n643), .A2(new_n548), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n524), .A2(new_n457), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT45), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n643), .A2(new_n517), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(KEYINPUT100), .B(KEYINPUT44), .Z(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n337), .A2(new_n359), .A3(new_n387), .ZN(new_n651));
  INV_X1    g450(.A(new_n357), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n520), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n427), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n423), .B1(new_n429), .B2(new_n430), .ZN(new_n655));
  AOI22_X1  g454(.A1(new_n653), .A2(new_n386), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n435), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT35), .B1(new_n653), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n389), .A2(new_n431), .A3(new_n432), .ZN(new_n659));
  AOI22_X1  g458(.A1(new_n651), .A2(new_n656), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n650), .B1(new_n660), .B2(new_n548), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT100), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n437), .A2(new_n549), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n648), .B1(new_n661), .B2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n521), .A2(new_n522), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n646), .B1(new_n457), .B2(new_n669), .ZN(G1328gat));
  NAND4_X1  g469(.A1(new_n614), .A2(new_n458), .A3(new_n357), .A4(new_n644), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n671), .B(KEYINPUT46), .Z(new_n672));
  AOI21_X1  g471(.A(new_n458), .B1(new_n667), .B2(new_n357), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n672), .A2(KEYINPUT101), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT101), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n671), .B(KEYINPUT46), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n676), .B1(new_n677), .B2(new_n673), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n675), .A2(new_n678), .ZN(G1329gat));
  AND4_X1   g478(.A1(new_n448), .A2(new_n614), .A3(new_n431), .A4(new_n644), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n667), .A2(new_n627), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n680), .B1(new_n681), .B2(G43gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g482(.A(G50gat), .B1(new_n636), .B2(new_n644), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n684), .B1(KEYINPUT102), .B2(KEYINPUT48), .ZN(new_n685));
  OR2_X1    g484(.A1(KEYINPUT102), .A2(KEYINPUT48), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n667), .A2(G50gat), .A3(new_n386), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n686), .B1(new_n685), .B2(new_n687), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n688), .A2(new_n689), .ZN(G1331gat));
  NOR4_X1   g489(.A1(new_n518), .A2(new_n578), .A3(new_n549), .A4(new_n609), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n437), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n523), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(new_n555), .ZN(G1332gat));
  INV_X1    g493(.A(new_n692), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT103), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n357), .B(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n698), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT104), .ZN(new_n701));
  NOR2_X1   g500(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1333gat));
  NOR3_X1   g502(.A1(new_n692), .A2(G71gat), .A3(new_n629), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n695), .A2(new_n627), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n704), .B1(G71gat), .B2(new_n705), .ZN(new_n706));
  XOR2_X1   g505(.A(KEYINPUT105), .B(KEYINPUT50), .Z(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1334gat));
  NAND2_X1  g507(.A1(new_n695), .A2(new_n386), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g509(.A1(new_n641), .A2(new_n518), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(new_n609), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n656), .A2(new_n651), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n658), .A2(new_n659), .ZN(new_n715));
  AOI211_X1 g514(.A(new_n548), .B(new_n664), .C1(new_n714), .C2(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n649), .B1(new_n437), .B2(new_n549), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n713), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(G85gat), .B1(new_n718), .B2(new_n523), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n437), .A2(new_n549), .A3(new_n711), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT51), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n548), .B1(new_n714), .B2(new_n715), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT51), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n722), .A2(new_n723), .A3(new_n711), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n668), .A2(new_n532), .A3(new_n608), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n719), .B1(new_n725), .B2(new_n726), .ZN(G1336gat));
  NAND2_X1  g526(.A1(new_n608), .A2(new_n533), .ZN(new_n728));
  OAI21_X1  g527(.A(KEYINPUT106), .B1(new_n698), .B2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT107), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT106), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n697), .A2(new_n731), .A3(new_n533), .A4(new_n608), .ZN(new_n732));
  AND3_X1   g531(.A1(new_n729), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n730), .B1(new_n729), .B2(new_n732), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n723), .A2(KEYINPUT108), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n736), .B1(new_n722), .B2(new_n711), .ZN(new_n737));
  AND4_X1   g536(.A1(new_n549), .A2(new_n437), .A3(new_n711), .A4(new_n736), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n735), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(KEYINPUT52), .ZN(new_n740));
  INV_X1    g539(.A(new_n713), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n741), .B1(new_n661), .B2(new_n666), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n533), .B1(new_n742), .B2(new_n357), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n697), .B(new_n713), .C1(new_n716), .C2(new_n717), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G92gat), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n729), .A2(new_n732), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n721), .A2(new_n724), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT52), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(KEYINPUT109), .B1(new_n744), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(G92gat), .B1(new_n718), .B2(new_n652), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT52), .ZN(new_n752));
  INV_X1    g551(.A(new_n736), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n720), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n722), .A2(new_n711), .A3(new_n736), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n752), .B1(new_n756), .B2(new_n735), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n751), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT109), .ZN(new_n759));
  INV_X1    g558(.A(new_n725), .ZN(new_n760));
  AOI22_X1  g559(.A1(new_n760), .A2(new_n747), .B1(new_n745), .B2(G92gat), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n758), .B(new_n759), .C1(new_n761), .C2(KEYINPUT52), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n750), .A2(new_n762), .ZN(G1337gat));
  INV_X1    g562(.A(new_n627), .ZN(new_n764));
  OAI21_X1  g563(.A(G99gat), .B1(new_n718), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n431), .A2(new_n527), .A3(new_n608), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n765), .B1(new_n725), .B2(new_n766), .ZN(G1338gat));
  INV_X1    g566(.A(KEYINPUT53), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n386), .B(new_n713), .C1(new_n716), .C2(new_n717), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(G106gat), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n386), .A2(new_n528), .A3(new_n608), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(KEYINPUT110), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT111), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n756), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n768), .B1(new_n770), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n528), .B1(new_n742), .B2(new_n386), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n721), .A2(new_n724), .A3(new_n772), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n768), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(KEYINPUT112), .B1(new_n775), .B2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT112), .ZN(new_n781));
  AOI22_X1  g580(.A1(new_n769), .A2(G106gat), .B1(new_n756), .B2(new_n773), .ZN(new_n782));
  OAI221_X1 g581(.A(new_n781), .B1(new_n776), .B2(new_n778), .C1(new_n782), .C2(new_n768), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n780), .A2(new_n783), .ZN(G1339gat));
  NOR2_X1   g583(.A1(new_n499), .A2(new_n500), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT114), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n511), .A2(new_n512), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n479), .B1(new_n788), .B2(new_n478), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n442), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n505), .A2(new_n506), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT18), .B1(new_n492), .B2(KEYINPUT90), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n504), .B1(new_n792), .B2(new_n496), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n608), .B(new_n790), .C1(new_n791), .C2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n591), .A2(new_n597), .A3(new_n592), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n595), .A2(KEYINPUT54), .A3(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n597), .B1(new_n591), .B2(new_n592), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n603), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(KEYINPUT55), .B1(new_n797), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n801), .A2(new_n605), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n797), .A2(KEYINPUT55), .A3(new_n800), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT113), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n803), .A2(new_n804), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n802), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n516), .A2(new_n505), .A3(new_n506), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n502), .B1(new_n514), .B2(new_n515), .ZN(new_n809));
  INV_X1    g608(.A(new_n443), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n807), .B1(new_n808), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(KEYINPUT115), .B1(new_n795), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT115), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n814), .B(new_n794), .C1(new_n517), .C2(new_n807), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n813), .A2(new_n548), .A3(new_n815), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n548), .A2(new_n807), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n817), .A2(new_n808), .A3(new_n790), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT116), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n641), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n816), .A2(KEYINPUT116), .A3(new_n818), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n610), .A2(new_n518), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n523), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n629), .A2(new_n386), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n826), .A2(new_n698), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(G113gat), .B1(new_n828), .B2(new_n517), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n824), .B1(new_n821), .B2(new_n822), .ZN(new_n830));
  NOR4_X1   g629(.A1(new_n830), .A2(new_n523), .A3(new_n657), .A4(new_n697), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(new_n291), .A3(new_n518), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n829), .A2(new_n832), .ZN(G1340gat));
  NOR3_X1   g632(.A1(new_n828), .A2(new_n285), .A3(new_n609), .ZN(new_n834));
  AOI21_X1  g633(.A(G120gat), .B1(new_n831), .B2(new_n608), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n834), .A2(new_n835), .ZN(G1341gat));
  OAI21_X1  g635(.A(G127gat), .B1(new_n828), .B2(new_n578), .ZN(new_n837));
  INV_X1    g636(.A(G127gat), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n831), .A2(new_n838), .A3(new_n641), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n839), .ZN(G1342gat));
  INV_X1    g639(.A(G134gat), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n357), .A2(new_n548), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n826), .A2(new_n841), .A3(new_n435), .A4(new_n842), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n843), .A2(KEYINPUT56), .ZN(new_n844));
  OAI21_X1  g643(.A(G134gat), .B1(new_n828), .B2(new_n548), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(KEYINPUT56), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(G1343gat));
  NAND3_X1  g646(.A1(new_n668), .A2(new_n764), .A3(new_n698), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n849), .B1(new_n830), .B2(new_n387), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n548), .B1(new_n795), .B2(new_n812), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n853), .A2(new_n818), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n851), .A2(new_n852), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n641), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI211_X1 g655(.A(KEYINPUT57), .B(new_n386), .C1(new_n856), .C2(new_n824), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n848), .B1(new_n850), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n263), .B1(new_n858), .B2(new_n518), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n860), .B1(new_n830), .B2(new_n523), .ZN(new_n861));
  AND3_X1   g660(.A1(new_n816), .A2(KEYINPUT116), .A3(new_n818), .ZN(new_n862));
  AOI21_X1  g661(.A(KEYINPUT116), .B1(new_n816), .B2(new_n818), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n862), .A2(new_n863), .A3(new_n641), .ZN(new_n864));
  OAI211_X1 g663(.A(KEYINPUT119), .B(new_n668), .C1(new_n864), .C2(new_n824), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n627), .A2(new_n387), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n861), .A2(new_n865), .A3(new_n698), .A4(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n517), .A2(G141gat), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT120), .B1(new_n859), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT58), .ZN(new_n872));
  INV_X1    g671(.A(new_n866), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n873), .B1(new_n826), .B2(KEYINPUT119), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n874), .A2(new_n698), .A3(new_n861), .A4(new_n868), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT118), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n872), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n878));
  AOI211_X1 g677(.A(new_n517), .B(new_n848), .C1(new_n850), .C2(new_n857), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n875), .B(new_n878), .C1(new_n879), .C2(new_n263), .ZN(new_n880));
  AND3_X1   g679(.A1(new_n871), .A2(new_n877), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n877), .B1(new_n871), .B2(new_n880), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n881), .A2(new_n882), .ZN(G1344gat));
  OAI21_X1  g682(.A(KEYINPUT59), .B1(new_n867), .B2(new_n609), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n265), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n858), .A2(new_n886), .A3(new_n608), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n830), .A2(new_n849), .A3(new_n387), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n641), .B1(new_n851), .B2(new_n818), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n386), .B1(new_n824), .B2(new_n889), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n890), .A2(new_n849), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  OR2_X1    g691(.A1(new_n848), .A2(new_n609), .ZN(new_n893));
  OAI211_X1 g692(.A(KEYINPUT59), .B(G148gat), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n885), .A2(new_n887), .A3(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT121), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n885), .A2(KEYINPUT121), .A3(new_n887), .A4(new_n894), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1345gat));
  AND2_X1   g698(.A1(new_n858), .A2(new_n641), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n641), .A2(new_n268), .ZN(new_n901));
  OAI22_X1  g700(.A1(new_n900), .A2(new_n268), .B1(new_n867), .B2(new_n901), .ZN(G1346gat));
  NAND4_X1  g701(.A1(new_n874), .A2(new_n269), .A3(new_n842), .A4(new_n861), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n858), .A2(new_n549), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n903), .B1(new_n904), .B2(new_n269), .ZN(G1347gat));
  NOR3_X1   g704(.A1(new_n830), .A2(new_n668), .A3(new_n698), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n906), .A2(new_n435), .ZN(new_n907));
  INV_X1    g706(.A(G169gat), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n907), .A2(new_n908), .A3(new_n518), .ZN(new_n909));
  XOR2_X1   g708(.A(new_n909), .B(KEYINPUT122), .Z(new_n910));
  NAND3_X1  g709(.A1(new_n523), .A2(new_n357), .A3(new_n827), .ZN(new_n911));
  OR2_X1    g710(.A1(new_n911), .A2(new_n830), .ZN(new_n912));
  OAI21_X1  g711(.A(G169gat), .B1(new_n912), .B2(new_n517), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n910), .A2(new_n913), .ZN(G1348gat));
  INV_X1    g713(.A(new_n912), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n915), .A2(G176gat), .A3(new_n608), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT123), .ZN(new_n917));
  AOI21_X1  g716(.A(G176gat), .B1(new_n907), .B2(new_n608), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n917), .A2(new_n918), .ZN(G1349gat));
  NAND3_X1  g718(.A1(new_n907), .A2(new_n641), .A3(new_n228), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT124), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n921), .B1(new_n912), .B2(new_n578), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(G183gat), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n912), .A2(new_n921), .A3(new_n578), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n920), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g725(.A(G190gat), .B1(new_n912), .B2(new_n548), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT61), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n907), .A2(new_n207), .A3(new_n549), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(G1351gat));
  NAND2_X1  g729(.A1(new_n906), .A2(new_n866), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n931), .A2(G197gat), .A3(new_n517), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n523), .A2(new_n357), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n933), .A2(new_n627), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n518), .B(new_n934), .C1(new_n888), .C2(new_n891), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n932), .B1(G197gat), .B2(new_n935), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n936), .B(KEYINPUT125), .ZN(G1352gat));
  INV_X1    g736(.A(new_n931), .ZN(new_n938));
  INV_X1    g737(.A(G204gat), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n938), .A2(new_n939), .A3(new_n608), .ZN(new_n940));
  OR3_X1    g739(.A1(new_n940), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n941));
  OAI21_X1  g740(.A(KEYINPUT126), .B1(new_n940), .B2(KEYINPUT62), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n892), .A2(new_n627), .A3(new_n933), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n939), .B1(new_n944), .B2(new_n608), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n945), .B1(KEYINPUT62), .B2(new_n940), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n943), .A2(new_n946), .ZN(G1353gat));
  NOR3_X1   g746(.A1(new_n931), .A2(G211gat), .A3(new_n578), .ZN(new_n948));
  OAI211_X1 g747(.A(new_n641), .B(new_n934), .C1(new_n888), .C2(new_n891), .ZN(new_n949));
  AOI21_X1  g748(.A(KEYINPUT63), .B1(new_n949), .B2(G211gat), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n950), .A2(new_n951), .ZN(new_n953));
  AND3_X1   g752(.A1(new_n949), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(G1354gat));
  AOI21_X1  g754(.A(G218gat), .B1(new_n938), .B2(new_n549), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n549), .A2(new_n238), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n956), .B1(new_n944), .B2(new_n957), .ZN(G1355gat));
endmodule


