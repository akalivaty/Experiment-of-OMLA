//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 1 1 0 1 1 1 1 0 1 0 0 1 1 0 1 1 0 0 1 1 0 1 0 1 1 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 1 0 1 1 1 0 1 0 1 0 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  INV_X1    g005(.A(G125), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT74), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT74), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G125), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  NOR3_X1   g010(.A1(new_n196), .A2(KEYINPUT16), .A3(G140), .ZN(new_n197));
  NOR2_X1   g011(.A1(G125), .A2(G140), .ZN(new_n198));
  XNOR2_X1  g012(.A(KEYINPUT74), .B(G125), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(G140), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT16), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT75), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n193), .A2(new_n195), .A3(G140), .ZN(new_n203));
  INV_X1    g017(.A(new_n198), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT75), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(KEYINPUT16), .ZN(new_n207));
  AOI211_X1 g021(.A(new_n191), .B(new_n197), .C1(new_n202), .C2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT64), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(new_n191), .ZN(new_n210));
  NAND2_X1  g024(.A1(KEYINPUT64), .A2(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AND2_X1   g026(.A1(G125), .A2(G140), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n212), .B1(new_n198), .B2(new_n213), .ZN(new_n214));
  XOR2_X1   g028(.A(KEYINPUT24), .B(G110), .Z(new_n215));
  INV_X1    g029(.A(G119), .ZN(new_n216));
  OR2_X1    g030(.A1(KEYINPUT67), .A2(G128), .ZN(new_n217));
  NAND2_X1  g031(.A1(KEYINPUT67), .A2(G128), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G128), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n220), .A2(G119), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT73), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  AND2_X1   g036(.A1(KEYINPUT67), .A2(G128), .ZN(new_n223));
  NOR2_X1   g037(.A1(KEYINPUT67), .A2(G128), .ZN(new_n224));
  OAI21_X1  g038(.A(G119), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT73), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n225), .B(new_n226), .C1(G119), .C2(new_n220), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n215), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n225), .B(KEYINPUT23), .C1(G119), .C2(new_n220), .ZN(new_n229));
  OR3_X1    g043(.A1(new_n216), .A2(KEYINPUT23), .A3(G128), .ZN(new_n230));
  AOI21_X1  g044(.A(G110), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n214), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n208), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n222), .A2(new_n227), .A3(new_n215), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n197), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n206), .B1(new_n205), .B2(KEYINPUT16), .ZN(new_n237));
  AOI211_X1 g051(.A(KEYINPUT75), .B(new_n201), .C1(new_n203), .C2(new_n204), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(new_n191), .ZN(new_n240));
  OAI211_X1 g054(.A(G146), .B(new_n236), .C1(new_n237), .C2(new_n238), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n235), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n229), .A2(G110), .A3(new_n230), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n233), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G953), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT70), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G953), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n249), .A2(G221), .A3(G234), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT22), .B(G137), .ZN(new_n253));
  XOR2_X1   g067(.A(new_n252), .B(new_n253), .Z(new_n254));
  OAI21_X1  g068(.A(KEYINPUT78), .B1(new_n244), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n202), .A2(new_n207), .ZN(new_n256));
  AOI21_X1  g070(.A(G146), .B1(new_n256), .B2(new_n236), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n243), .B(new_n234), .C1(new_n257), .C2(new_n208), .ZN(new_n258));
  OR2_X1    g072(.A1(new_n208), .A2(new_n232), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT78), .ZN(new_n261));
  INV_X1    g075(.A(new_n254), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n255), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n258), .A2(new_n259), .A3(new_n254), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT79), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n258), .A2(new_n259), .A3(new_n254), .A4(KEYINPUT79), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n264), .A2(new_n188), .A3(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT25), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n255), .A2(new_n263), .B1(new_n267), .B2(new_n268), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n273), .A2(KEYINPUT25), .A3(new_n188), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n190), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n189), .A2(G902), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n276), .B(KEYINPUT80), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n275), .B1(new_n278), .B2(new_n273), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n257), .A2(new_n208), .ZN(new_n280));
  AOI21_X1  g094(.A(G237), .B1(new_n246), .B2(new_n248), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n281), .A2(G143), .A3(G214), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(G143), .B1(new_n281), .B2(G214), .ZN(new_n284));
  OAI211_X1 g098(.A(KEYINPUT17), .B(G131), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(G131), .B1(new_n283), .B2(new_n284), .ZN(new_n286));
  INV_X1    g100(.A(G237), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n249), .A2(G214), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G143), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G131), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n290), .A2(new_n291), .A3(new_n282), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n286), .A2(new_n292), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n280), .B(new_n285), .C1(KEYINPUT17), .C2(new_n293), .ZN(new_n294));
  XNOR2_X1  g108(.A(G113), .B(G122), .ZN(new_n295));
  INV_X1    g109(.A(G104), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n295), .B(new_n296), .ZN(new_n297));
  OAI211_X1 g111(.A(KEYINPUT18), .B(G131), .C1(new_n283), .C2(new_n284), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n200), .A2(G146), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n214), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT18), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n290), .B(new_n282), .C1(new_n302), .C2(new_n291), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT93), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n303), .A2(KEYINPUT93), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n301), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n294), .A2(new_n297), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n297), .B1(new_n294), .B2(new_n307), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n188), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G475), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT94), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n298), .A2(new_n300), .ZN(new_n314));
  OR2_X1    g128(.A1(new_n303), .A2(KEYINPUT93), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n314), .B1(new_n315), .B2(new_n304), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n213), .A2(new_n198), .ZN(new_n317));
  MUX2_X1   g131(.A(new_n317), .B(new_n205), .S(KEYINPUT19), .Z(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n212), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n293), .A2(new_n241), .A3(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n313), .B1(new_n316), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n293), .A2(new_n241), .A3(new_n319), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n307), .A2(KEYINPUT94), .A3(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n297), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n321), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n308), .ZN(new_n326));
  INV_X1    g140(.A(G475), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n327), .A3(new_n188), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n328), .A2(KEYINPUT20), .ZN(new_n329));
  XOR2_X1   g143(.A(KEYINPUT92), .B(KEYINPUT20), .Z(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(G475), .B1(new_n325), .B2(new_n308), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n331), .B1(new_n332), .B2(new_n188), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n312), .B1(new_n329), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(G134), .ZN(new_n335));
  OAI21_X1  g149(.A(G143), .B1(new_n223), .B2(new_n224), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT13), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n335), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT96), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n339), .B1(new_n220), .B2(G143), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n289), .A2(KEYINPUT96), .A3(G128), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n336), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n338), .B(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G122), .ZN(new_n344));
  OAI21_X1  g158(.A(KEYINPUT95), .B1(new_n344), .B2(G116), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT95), .ZN(new_n346));
  INV_X1    g160(.A(G116), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n347), .A3(G122), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n349), .B1(new_n347), .B2(G122), .ZN(new_n350));
  INV_X1    g164(.A(G107), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n350), .B(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n343), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n342), .A2(new_n335), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n354), .B1(G107), .B2(new_n350), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n347), .A2(G122), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n356), .B1(new_n349), .B2(KEYINPUT14), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT97), .ZN(new_n358));
  OR2_X1    g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n358), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n359), .B(new_n360), .C1(KEYINPUT14), .C2(new_n349), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n355), .B1(new_n361), .B2(G107), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n342), .A2(new_n335), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n353), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  XOR2_X1   g179(.A(KEYINPUT9), .B(G234), .Z(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NOR3_X1   g181(.A1(new_n367), .A2(new_n187), .A3(G953), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n368), .ZN(new_n370));
  AOI211_X1 g184(.A(new_n363), .B(new_n355), .C1(new_n361), .C2(G107), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n370), .B1(new_n371), .B2(new_n353), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n188), .ZN(new_n374));
  INV_X1    g188(.A(G478), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n375), .A2(KEYINPUT15), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n374), .A2(new_n376), .ZN(new_n379));
  INV_X1    g193(.A(G952), .ZN(new_n380));
  AOI211_X1 g194(.A(G953), .B(new_n380), .C1(G234), .C2(G237), .ZN(new_n381));
  AOI211_X1 g195(.A(new_n188), .B(new_n249), .C1(G234), .C2(G237), .ZN(new_n382));
  XOR2_X1   g196(.A(KEYINPUT21), .B(G898), .Z(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n381), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n378), .A2(new_n379), .A3(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n334), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n335), .A2(G137), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(KEYINPUT11), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n335), .A2(G137), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT11), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n392), .B1(new_n335), .B2(G137), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n390), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(KEYINPUT66), .B1(new_n335), .B2(G137), .ZN(new_n395));
  MUX2_X1   g209(.A(new_n395), .B(KEYINPUT66), .S(new_n389), .Z(new_n396));
  MUX2_X1   g210(.A(new_n394), .B(new_n396), .S(G131), .Z(new_n397));
  NAND3_X1  g211(.A1(new_n210), .A2(new_n289), .A3(new_n211), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT65), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n289), .A2(G146), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT65), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n210), .A2(new_n402), .A3(new_n289), .A4(new_n211), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n399), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n289), .B1(new_n210), .B2(new_n211), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT1), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n217), .B(new_n218), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT69), .ZN(new_n409));
  AND2_X1   g223(.A1(KEYINPUT64), .A2(G146), .ZN(new_n410));
  NOR2_X1   g224(.A1(KEYINPUT64), .A2(G146), .ZN(new_n411));
  OAI21_X1  g225(.A(G143), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n191), .A2(G143), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n412), .A2(new_n406), .A3(G128), .A4(new_n414), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n408), .A2(new_n409), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n409), .B1(new_n408), .B2(new_n415), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n397), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  XOR2_X1   g232(.A(KEYINPUT0), .B(G128), .Z(new_n419));
  NAND2_X1  g233(.A1(new_n404), .A2(new_n419), .ZN(new_n420));
  NOR3_X1   g234(.A1(new_n405), .A2(new_n220), .A3(new_n413), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT0), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n394), .B(new_n291), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n418), .A2(KEYINPUT30), .A3(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(KEYINPUT2), .B(G113), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n216), .A2(G116), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n347), .A2(G119), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT68), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n429), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n432), .A2(new_n428), .A3(KEYINPUT68), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT30), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n408), .A2(new_n415), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n397), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n438), .B1(new_n440), .B2(new_n425), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n427), .A2(new_n437), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n437), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n418), .A2(new_n443), .A3(new_n426), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n281), .A2(G210), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n445), .B(G101), .ZN(new_n446));
  XNOR2_X1  g260(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n446), .B(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n442), .A2(new_n444), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(KEYINPUT31), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT31), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n442), .A2(new_n451), .A3(new_n444), .A4(new_n448), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n440), .A2(new_n425), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n453), .A2(new_n443), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n444), .A2(KEYINPUT28), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT28), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n418), .A2(new_n456), .A3(new_n426), .A4(new_n443), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n454), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n450), .B(new_n452), .C1(new_n458), .C2(new_n448), .ZN(new_n459));
  NOR2_X1   g273(.A1(G472), .A2(G902), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n459), .A2(KEYINPUT32), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(KEYINPUT32), .B1(new_n459), .B2(new_n460), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n448), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n442), .A2(new_n444), .A3(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n465), .B1(new_n458), .B2(new_n464), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT29), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n443), .B1(new_n418), .B2(new_n426), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n448), .A2(KEYINPUT29), .ZN(new_n470));
  AOI211_X1 g284(.A(new_n469), .B(new_n470), .C1(new_n455), .C2(new_n457), .ZN(new_n471));
  OAI21_X1  g285(.A(KEYINPUT71), .B1(new_n471), .B2(G902), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n455), .A2(new_n457), .ZN(new_n473));
  INV_X1    g287(.A(new_n469), .ZN(new_n474));
  INV_X1    g288(.A(new_n470), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT71), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(new_n477), .A3(new_n188), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n468), .A2(new_n472), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G472), .ZN(new_n480));
  AOI21_X1  g294(.A(KEYINPUT72), .B1(new_n463), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n450), .A2(new_n452), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n458), .A2(new_n448), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n460), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT32), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n459), .A2(KEYINPUT32), .A3(new_n460), .ZN(new_n487));
  AND4_X1   g301(.A1(KEYINPUT72), .A2(new_n480), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n279), .B(new_n388), .C1(new_n481), .C2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT91), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT90), .ZN(new_n491));
  OAI21_X1  g305(.A(G210), .B1(G237), .B2(G902), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n430), .A2(new_n431), .A3(KEYINPUT5), .ZN(new_n493));
  OAI21_X1  g307(.A(G113), .B1(new_n430), .B2(KEYINPUT5), .ZN(new_n494));
  OAI21_X1  g308(.A(KEYINPUT86), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n430), .A2(new_n431), .A3(KEYINPUT5), .ZN(new_n496));
  OR3_X1    g310(.A1(new_n347), .A2(KEYINPUT5), .A3(G119), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT86), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n496), .A2(new_n497), .A3(new_n498), .A4(G113), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n433), .A2(new_n429), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n495), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n351), .A2(KEYINPUT81), .A3(G104), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT3), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n351), .A2(G104), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(G101), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT3), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n507), .A2(new_n351), .A3(KEYINPUT81), .A4(G104), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n503), .A2(new_n505), .A3(new_n506), .A4(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n296), .A2(G107), .ZN(new_n510));
  OAI21_X1  g324(.A(G101), .B1(new_n504), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(KEYINPUT87), .B1(new_n501), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n503), .A2(new_n505), .A3(new_n508), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(G101), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n515), .A2(KEYINPUT4), .A3(new_n509), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT4), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(new_n517), .A3(G101), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n516), .A2(new_n518), .A3(new_n437), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n509), .A2(new_n511), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n496), .A2(new_n497), .A3(G113), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n521), .A2(KEYINPUT86), .B1(new_n433), .B2(new_n429), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT87), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n520), .A2(new_n522), .A3(new_n523), .A4(new_n499), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n513), .A2(new_n519), .A3(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(G110), .B(G122), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT88), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n513), .A2(new_n519), .A3(new_n524), .A4(new_n526), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n528), .A2(new_n529), .A3(KEYINPUT6), .A4(new_n530), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n528), .A2(KEYINPUT6), .A3(new_n530), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT6), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n525), .A2(new_n533), .A3(new_n527), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT88), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n531), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n196), .B1(new_n420), .B2(new_n422), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n408), .A2(new_n415), .A3(new_n196), .ZN(new_n539));
  INV_X1    g353(.A(G224), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n540), .A2(G953), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n538), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n408), .A2(new_n415), .A3(new_n196), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n541), .B1(new_n544), .B2(new_n537), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n536), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n500), .A2(new_n521), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n520), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n526), .B(KEYINPUT8), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n549), .B(new_n550), .C1(new_n520), .C2(new_n501), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT89), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n544), .A2(new_n537), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n542), .A2(KEYINPUT7), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n554), .B1(new_n539), .B2(KEYINPUT89), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n551), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n538), .A2(KEYINPUT7), .A3(new_n539), .A4(new_n542), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n530), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n188), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n492), .B1(new_n547), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n492), .ZN(new_n562));
  AOI211_X1 g376(.A(new_n562), .B(new_n559), .C1(new_n536), .C2(new_n546), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n491), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n547), .A2(new_n492), .A3(new_n560), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT90), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(G214), .B1(G237), .B2(G902), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n490), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n546), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n528), .A2(KEYINPUT6), .A3(new_n530), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n571), .A2(KEYINPUT88), .A3(new_n534), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n570), .B1(new_n572), .B2(new_n531), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n562), .B1(new_n573), .B2(new_n559), .ZN(new_n574));
  AOI21_X1  g388(.A(KEYINPUT90), .B1(new_n565), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n563), .A2(new_n491), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n490), .B(new_n568), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n569), .A2(new_n578), .ZN(new_n579));
  OAI211_X1 g393(.A(KEYINPUT10), .B(new_n520), .C1(new_n416), .C2(new_n417), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT10), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT82), .ZN(new_n582));
  OAI21_X1  g396(.A(G128), .B1(new_n400), .B2(new_n406), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n583), .B1(new_n405), .B2(new_n413), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n415), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n520), .A2(new_n582), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n582), .B1(new_n520), .B2(new_n585), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n581), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n516), .A2(new_n420), .A3(new_n422), .A4(new_n518), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n580), .A2(new_n424), .A3(new_n588), .A4(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n520), .A2(new_n585), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT82), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n520), .A2(new_n585), .A3(new_n582), .ZN(new_n593));
  AOI22_X1  g407(.A1(new_n404), .A2(new_n407), .B1(new_n421), .B2(new_n406), .ZN(new_n594));
  AOI22_X1  g408(.A1(new_n592), .A2(new_n593), .B1(new_n512), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT12), .ZN(new_n596));
  NOR3_X1   g410(.A1(new_n595), .A2(new_n596), .A3(new_n424), .ZN(new_n597));
  OAI22_X1  g411(.A1(new_n586), .A2(new_n587), .B1(new_n439), .B2(new_n520), .ZN(new_n598));
  INV_X1    g412(.A(new_n424), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT12), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n590), .B1(new_n597), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n249), .A2(G227), .ZN(new_n602));
  XNOR2_X1  g416(.A(G110), .B(G140), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n580), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n588), .A2(new_n589), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n599), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n609), .A2(new_n590), .A3(new_n604), .ZN(new_n610));
  AOI21_X1  g424(.A(G902), .B1(new_n606), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(G469), .ZN(new_n612));
  OAI21_X1  g426(.A(KEYINPUT83), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n590), .A2(new_n604), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n588), .A2(new_n589), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n424), .B1(new_n615), .B2(new_n580), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n596), .B1(new_n595), .B2(new_n424), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n598), .A2(KEYINPUT12), .A3(new_n599), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n604), .B1(new_n620), .B2(new_n590), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n188), .B1(new_n617), .B2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT83), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n622), .A2(new_n623), .A3(G469), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT84), .B(G469), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n620), .A2(new_n590), .A3(new_n604), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n604), .B1(new_n609), .B2(new_n590), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n188), .B(new_n626), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n613), .A2(new_n624), .A3(new_n630), .ZN(new_n631));
  OAI21_X1  g445(.A(G221), .B1(new_n367), .B2(G902), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT85), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n631), .A2(KEYINPUT85), .A3(new_n632), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n579), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n489), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(new_n506), .ZN(G3));
  NAND2_X1  g454(.A1(new_n459), .A2(new_n188), .ZN(new_n641));
  AOI22_X1  g455(.A1(new_n641), .A2(G472), .B1(new_n460), .B2(new_n459), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  AND4_X1   g457(.A1(KEYINPUT25), .A2(new_n264), .A3(new_n188), .A4(new_n269), .ZN(new_n644));
  AOI21_X1  g458(.A(KEYINPUT25), .B1(new_n273), .B2(new_n188), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n189), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n273), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n646), .B1(new_n277), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n643), .A2(new_n648), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n637), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT98), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n372), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n373), .A2(new_n652), .A3(KEYINPUT33), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT33), .ZN(new_n654));
  OAI211_X1 g468(.A(new_n369), .B(new_n372), .C1(new_n651), .C2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n653), .A2(G478), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n373), .A2(new_n375), .A3(new_n188), .ZN(new_n657));
  NAND2_X1  g471(.A1(G478), .A2(G902), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n334), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n568), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n661), .B1(new_n565), .B2(new_n574), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n660), .A2(new_n385), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n650), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT34), .B(G104), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G6));
  NOR2_X1   g481(.A1(new_n663), .A2(new_n385), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n328), .A2(new_n330), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n333), .ZN(new_n670));
  INV_X1    g484(.A(new_n379), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n671), .A2(new_n377), .ZN(new_n672));
  INV_X1    g486(.A(new_n312), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n670), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n650), .A2(new_n668), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G107), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT99), .B(KEYINPUT35), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G9));
  INV_X1    g492(.A(KEYINPUT100), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n262), .A2(KEYINPUT36), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(new_n260), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n278), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n679), .B1(new_n275), .B2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n646), .A2(KEYINPUT100), .A3(new_n682), .ZN(new_n685));
  AND4_X1   g499(.A1(new_n388), .A2(new_n684), .A3(new_n685), .A4(new_n642), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n579), .A2(new_n686), .A3(new_n637), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT37), .B(G110), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G12));
  INV_X1    g503(.A(G900), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n381), .B1(new_n382), .B2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n674), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT72), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n486), .A2(new_n487), .ZN(new_n695));
  INV_X1    g509(.A(G472), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n471), .A2(KEYINPUT71), .A3(G902), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n477), .B1(new_n476), .B2(new_n188), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n696), .B1(new_n699), .B2(new_n468), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n694), .B1(new_n695), .B2(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n480), .A2(new_n486), .A3(KEYINPUT72), .A4(new_n487), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n693), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n684), .A2(new_n685), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n704), .B1(new_n635), .B2(new_n636), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n703), .A2(new_n705), .A3(new_n662), .ZN(new_n706));
  XOR2_X1   g520(.A(KEYINPUT101), .B(G128), .Z(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G30));
  INV_X1    g522(.A(new_n334), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n691), .B(KEYINPUT39), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n710), .B1(new_n635), .B2(new_n636), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT40), .ZN(new_n712));
  AOI211_X1 g526(.A(new_n709), .B(new_n672), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n442), .A2(new_n444), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n448), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n474), .A2(new_n444), .A3(new_n464), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT102), .ZN(new_n718));
  AOI21_X1  g532(.A(G902), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n719), .B1(new_n718), .B2(new_n717), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(G472), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n463), .ZN(new_n722));
  OR2_X1    g536(.A1(new_n711), .A2(new_n712), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n575), .A2(new_n576), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(KEYINPUT38), .ZN(new_n725));
  INV_X1    g539(.A(new_n704), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n725), .A2(new_n726), .A3(new_n661), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n713), .A2(new_n722), .A3(new_n723), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G143), .ZN(G45));
  NAND3_X1  g543(.A1(new_n334), .A2(new_n659), .A3(new_n692), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n730), .B1(new_n701), .B2(new_n702), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(new_n705), .A3(new_n662), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G146), .ZN(G48));
  NAND2_X1  g547(.A1(new_n701), .A2(new_n702), .ZN(new_n734));
  INV_X1    g548(.A(new_n630), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n188), .B1(new_n628), .B2(new_n629), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n735), .B1(G469), .B2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n632), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n734), .A2(new_n279), .A3(new_n664), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(KEYINPUT41), .B(G113), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(G15));
  NOR3_X1   g557(.A1(new_n738), .A2(new_n739), .A3(new_n663), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n279), .A2(new_n674), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n734), .A2(new_n386), .A3(new_n744), .A4(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G116), .ZN(G18));
  INV_X1    g561(.A(new_n388), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n704), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n734), .A2(new_n749), .A3(new_n744), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G119), .ZN(G21));
  AOI21_X1  g565(.A(new_n469), .B1(new_n455), .B2(new_n457), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n450), .B(new_n452), .C1(new_n448), .C2(new_n752), .ZN(new_n753));
  AOI22_X1  g567(.A1(new_n641), .A2(G472), .B1(new_n460), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n279), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n709), .A2(new_n672), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n756), .A2(new_n668), .A3(new_n740), .A4(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G122), .ZN(G24));
  NAND3_X1  g573(.A1(new_n684), .A2(new_n685), .A3(new_n754), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(KEYINPUT103), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT103), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n684), .A2(new_n685), .A3(new_n754), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NOR4_X1   g578(.A1(new_n738), .A2(new_n730), .A3(new_n739), .A4(new_n663), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G125), .ZN(G27));
  OAI21_X1  g581(.A(new_n630), .B1(new_n612), .B2(new_n611), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n739), .A2(new_n661), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n564), .A2(new_n566), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n770), .A2(new_n730), .A3(KEYINPUT42), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n734), .A2(new_n279), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n770), .ZN(new_n773));
  INV_X1    g587(.A(new_n730), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n480), .A2(new_n486), .A3(new_n487), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n279), .ZN(new_n777));
  OAI21_X1  g591(.A(KEYINPUT42), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n772), .A2(new_n778), .ZN(new_n779));
  XOR2_X1   g593(.A(KEYINPUT104), .B(G131), .Z(new_n780));
  XNOR2_X1  g594(.A(new_n779), .B(new_n780), .ZN(G33));
  INV_X1    g595(.A(new_n693), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n734), .A2(new_n279), .A3(new_n782), .A4(new_n773), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G134), .ZN(G36));
  NAND2_X1  g598(.A1(new_n606), .A2(new_n610), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(KEYINPUT45), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(G469), .ZN(new_n787));
  NAND2_X1  g601(.A1(G469), .A2(G902), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n787), .A2(KEYINPUT46), .A3(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT46), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n790), .B(G469), .C1(new_n786), .C2(G902), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n789), .A2(new_n630), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n632), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT105), .ZN(new_n794));
  OR3_X1    g608(.A1(new_n793), .A2(new_n794), .A3(new_n710), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n794), .B1(new_n793), .B2(new_n710), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT44), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n726), .A2(KEYINPUT106), .A3(new_n643), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT106), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n800), .B1(new_n704), .B2(new_n642), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n709), .A2(new_n659), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(KEYINPUT43), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n798), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n567), .A2(new_n661), .ZN(new_n806));
  INV_X1    g620(.A(new_n804), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n807), .A2(KEYINPUT44), .A3(new_n801), .A4(new_n799), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n797), .A2(new_n805), .A3(new_n806), .A4(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G137), .ZN(G39));
  NOR2_X1   g624(.A1(new_n481), .A2(new_n488), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n811), .A2(new_n648), .A3(new_n774), .A4(new_n806), .ZN(new_n812));
  OR2_X1    g626(.A1(new_n812), .A2(KEYINPUT107), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(KEYINPUT107), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT47), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n793), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n792), .A2(KEYINPUT47), .A3(new_n632), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n813), .A2(new_n814), .A3(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G140), .ZN(G42));
  NOR2_X1   g634(.A1(new_n380), .A2(G953), .ZN(new_n821));
  XOR2_X1   g635(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n822));
  OAI211_X1 g636(.A(new_n816), .B(new_n817), .C1(new_n632), .C2(new_n738), .ZN(new_n823));
  INV_X1    g637(.A(new_n381), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n804), .A2(new_n824), .A3(new_n755), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n823), .A2(new_n806), .A3(new_n825), .ZN(new_n826));
  XOR2_X1   g640(.A(new_n826), .B(KEYINPUT114), .Z(new_n827));
  AND4_X1   g641(.A1(new_n724), .A2(new_n737), .A3(new_n381), .A4(new_n769), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n807), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n764), .ZN(new_n830));
  AND4_X1   g644(.A1(new_n279), .A2(new_n828), .A3(new_n463), .A4(new_n721), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n334), .A2(new_n659), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n825), .A2(new_n661), .A3(new_n725), .A4(new_n740), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT50), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n834), .A2(new_n835), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n830), .B(new_n833), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n822), .B1(new_n827), .B2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n777), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n829), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT48), .ZN(new_n843));
  INV_X1    g657(.A(new_n838), .ZN(new_n844));
  AOI22_X1  g658(.A1(new_n844), .A2(new_n836), .B1(new_n831), .B2(new_n832), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n845), .A2(KEYINPUT51), .A3(new_n830), .A4(new_n826), .ZN(new_n846));
  AND4_X1   g660(.A1(new_n821), .A2(new_n840), .A3(new_n843), .A4(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n831), .A2(new_n334), .A3(new_n659), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n783), .A2(new_n778), .A3(new_n772), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n811), .A2(new_n673), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n378), .A2(new_n379), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n670), .A2(new_n851), .A3(new_n691), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n850), .A2(new_n705), .A3(new_n806), .A4(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n775), .B1(new_n761), .B2(new_n763), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n854), .A2(KEYINPUT111), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n854), .A2(KEYINPUT111), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n849), .B(new_n853), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n741), .A2(new_n750), .A3(new_n758), .ZN(new_n858));
  INV_X1    g672(.A(new_n638), .ZN(new_n859));
  AOI211_X1 g673(.A(new_n648), .B(new_n748), .C1(new_n701), .C2(new_n702), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n859), .B1(new_n860), .B2(new_n686), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n851), .B(new_n312), .C1(new_n333), .C2(new_n329), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n385), .B1(new_n862), .B2(new_n660), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n579), .A2(new_n637), .A3(new_n649), .A4(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n858), .A2(new_n746), .A3(new_n861), .A4(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n857), .A2(new_n865), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n709), .A2(new_n663), .A3(new_n672), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n646), .A2(new_n682), .A3(new_n768), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n691), .A2(new_n739), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n722), .A2(new_n867), .A3(new_n868), .A4(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n706), .A2(new_n766), .A3(new_n732), .A4(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT52), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n662), .B(new_n705), .C1(new_n703), .C2(new_n731), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT52), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n873), .A2(new_n874), .A3(new_n766), .A4(new_n870), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n866), .A2(new_n876), .A3(KEYINPUT53), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT53), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n783), .A2(new_n778), .A3(new_n772), .ZN(new_n879));
  OR2_X1    g693(.A1(new_n854), .A2(KEYINPUT111), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n854), .A2(KEYINPUT111), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n741), .A2(new_n746), .A3(new_n750), .A4(new_n758), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n864), .B(new_n687), .C1(new_n638), .C2(new_n489), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n882), .A2(new_n885), .A3(new_n853), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n872), .A2(new_n875), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n878), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n877), .A2(new_n888), .A3(KEYINPUT112), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT112), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n890), .B(new_n878), .C1(new_n886), .C2(new_n887), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n889), .A2(KEYINPUT54), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n877), .A2(new_n888), .ZN(new_n893));
  OR2_X1    g707(.A1(new_n893), .A2(KEYINPUT54), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n847), .A2(new_n848), .A3(new_n892), .A4(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n825), .A2(new_n744), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT115), .ZN(new_n897));
  OAI22_X1  g711(.A1(new_n895), .A2(new_n897), .B1(G952), .B2(G953), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n738), .A2(KEYINPUT49), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(KEYINPUT110), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(new_n725), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n279), .A2(new_n769), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT108), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n803), .B1(new_n738), .B2(KEYINPUT49), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  AOI211_X1 g720(.A(new_n722), .B(new_n901), .C1(new_n906), .C2(KEYINPUT109), .ZN(new_n907));
  OAI221_X1 g721(.A(new_n907), .B1(KEYINPUT109), .B2(new_n906), .C1(KEYINPUT110), .C2(new_n899), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n898), .A2(new_n908), .ZN(G75));
  XNOR2_X1  g723(.A(new_n536), .B(new_n570), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT55), .Z(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n188), .B1(new_n877), .B2(new_n888), .ZN(new_n913));
  AOI21_X1  g727(.A(KEYINPUT56), .B1(new_n913), .B2(G210), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT116), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n912), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n249), .A2(G952), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT117), .Z(new_n918));
  AOI21_X1  g732(.A(new_n918), .B1(new_n914), .B2(new_n915), .ZN(new_n919));
  INV_X1    g733(.A(G210), .ZN(new_n920));
  AOI211_X1 g734(.A(new_n920), .B(new_n188), .C1(new_n877), .C2(new_n888), .ZN(new_n921));
  OAI211_X1 g735(.A(KEYINPUT116), .B(new_n911), .C1(new_n921), .C2(KEYINPUT56), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n916), .A2(new_n919), .A3(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT118), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n916), .A2(new_n919), .A3(KEYINPUT118), .A4(new_n922), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(G51));
  XNOR2_X1  g741(.A(new_n893), .B(KEYINPUT54), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n788), .A2(KEYINPUT57), .ZN(new_n929));
  OR2_X1    g743(.A1(new_n788), .A2(KEYINPUT57), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n931), .B1(new_n629), .B2(new_n628), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n913), .A2(G469), .A3(new_n786), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n917), .B1(new_n932), .B2(new_n933), .ZN(G54));
  AND3_X1   g748(.A1(new_n913), .A2(KEYINPUT58), .A3(G475), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n935), .A2(new_n326), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n935), .A2(new_n326), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n936), .A2(new_n937), .A3(new_n917), .ZN(G60));
  NAND2_X1  g752(.A1(new_n653), .A2(new_n655), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n658), .B(KEYINPUT59), .Z(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n928), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n918), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n940), .B1(new_n894), .B2(new_n892), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n942), .B(new_n943), .C1(new_n939), .C2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(G63));
  OAI21_X1  g760(.A(KEYINPUT60), .B1(new_n187), .B2(new_n188), .ZN(new_n947));
  OR3_X1    g761(.A1(new_n187), .A2(new_n188), .A3(KEYINPUT60), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n893), .A2(new_n681), .A3(new_n947), .A4(new_n948), .ZN(new_n949));
  OR2_X1    g763(.A1(new_n949), .A2(KEYINPUT119), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n893), .A2(new_n947), .A3(new_n948), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n918), .B1(new_n951), .B2(new_n647), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n949), .A2(KEYINPUT119), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n950), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT61), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n950), .A2(KEYINPUT61), .A3(new_n952), .A4(new_n953), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(G66));
  NAND2_X1  g772(.A1(new_n865), .A2(new_n249), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT120), .ZN(new_n960));
  OAI21_X1  g774(.A(G953), .B1(new_n384), .B2(new_n540), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n572), .B(new_n531), .C1(G898), .C2(new_n249), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(G69));
  AOI21_X1  g778(.A(new_n249), .B1(G227), .B2(G900), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n427), .A2(new_n441), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(new_n318), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n862), .A2(new_n660), .ZN(new_n970));
  AOI211_X1 g784(.A(new_n648), .B(new_n811), .C1(KEYINPUT123), .C2(new_n970), .ZN(new_n971));
  OR2_X1    g785(.A1(new_n970), .A2(KEYINPUT123), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n971), .A2(new_n711), .A3(new_n806), .A4(new_n972), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n809), .A2(new_n819), .A3(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT121), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n706), .A2(new_n732), .ZN(new_n976));
  INV_X1    g790(.A(new_n766), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n975), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n873), .A2(KEYINPUT121), .A3(new_n766), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n978), .A2(new_n728), .A3(new_n979), .ZN(new_n980));
  XOR2_X1   g794(.A(KEYINPUT122), .B(KEYINPUT62), .Z(new_n981));
  OR2_X1    g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n980), .B1(KEYINPUT122), .B2(KEYINPUT62), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n974), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n969), .B1(new_n984), .B2(new_n249), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n795), .A2(new_n841), .A3(new_n796), .A4(new_n867), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n987), .A2(KEYINPUT124), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n987), .A2(KEYINPUT124), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n849), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n809), .A2(new_n819), .A3(new_n978), .A4(new_n979), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n249), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n246), .A2(new_n248), .A3(new_n690), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(KEYINPUT125), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT125), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n992), .A2(new_n996), .A3(new_n993), .ZN(new_n997));
  AND2_X1   g811(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  OAI211_X1 g812(.A(new_n966), .B(new_n986), .C1(new_n998), .C2(new_n968), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n968), .B1(new_n995), .B2(new_n997), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n965), .B1(new_n1000), .B2(new_n985), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n999), .A2(new_n1001), .ZN(G72));
  XNOR2_X1  g816(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n696), .A2(new_n188), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1003), .B(new_n1004), .Z(new_n1005));
  OR2_X1    g819(.A1(new_n990), .A2(new_n991), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1005), .B1(new_n1006), .B2(new_n865), .ZN(new_n1007));
  INV_X1    g821(.A(new_n465), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n917), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1005), .B1(new_n984), .B2(new_n865), .ZN(new_n1010));
  INV_X1    g824(.A(new_n715), .ZN(new_n1011));
  AND3_X1   g825(.A1(new_n1010), .A2(KEYINPUT127), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(KEYINPUT127), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1009), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n889), .A2(new_n715), .A3(new_n891), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n1015), .A2(new_n1008), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1014), .B1(new_n1005), .B2(new_n1016), .ZN(G57));
endmodule


