

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588;

  NOR2_X1 U322 ( .A1(n578), .A2(n384), .ZN(n385) );
  XNOR2_X1 U323 ( .A(n367), .B(G127GAT), .ZN(n368) );
  XNOR2_X1 U324 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U325 ( .A(n389), .B(KEYINPUT64), .ZN(n390) );
  XNOR2_X1 U326 ( .A(n391), .B(n390), .ZN(n539) );
  INV_X1 U327 ( .A(KEYINPUT58), .ZN(n451) );
  XOR2_X1 U328 ( .A(n377), .B(n376), .Z(n582) );
  XNOR2_X1 U329 ( .A(n451), .B(G190GAT), .ZN(n452) );
  XNOR2_X1 U330 ( .A(n453), .B(n452), .ZN(G1351GAT) );
  XOR2_X1 U331 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n291) );
  XNOR2_X1 U332 ( .A(G183GAT), .B(KEYINPUT18), .ZN(n290) );
  XNOR2_X1 U333 ( .A(n291), .B(n290), .ZN(n441) );
  XOR2_X1 U334 ( .A(G197GAT), .B(KEYINPUT21), .Z(n293) );
  XNOR2_X1 U335 ( .A(G218GAT), .B(G211GAT), .ZN(n292) );
  XNOR2_X1 U336 ( .A(n293), .B(n292), .ZN(n416) );
  XNOR2_X1 U337 ( .A(n441), .B(n416), .ZN(n303) );
  XOR2_X1 U338 ( .A(G8GAT), .B(G169GAT), .Z(n305) );
  XOR2_X1 U339 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n298) );
  XNOR2_X1 U340 ( .A(G36GAT), .B(KEYINPUT75), .ZN(n294) );
  XNOR2_X1 U341 ( .A(n294), .B(G190GAT), .ZN(n353) );
  XOR2_X1 U342 ( .A(G204GAT), .B(G176GAT), .Z(n296) );
  XNOR2_X1 U343 ( .A(G92GAT), .B(G64GAT), .ZN(n295) );
  XNOR2_X1 U344 ( .A(n296), .B(n295), .ZN(n322) );
  XNOR2_X1 U345 ( .A(n353), .B(n322), .ZN(n297) );
  XNOR2_X1 U346 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U347 ( .A(n305), .B(n299), .Z(n301) );
  NAND2_X1 U348 ( .A1(G226GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U349 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U350 ( .A(n303), .B(n302), .Z(n516) );
  INV_X1 U351 ( .A(n516), .ZN(n492) );
  XNOR2_X1 U352 ( .A(G1GAT), .B(G15GAT), .ZN(n304) );
  XNOR2_X1 U353 ( .A(n304), .B(G22GAT), .ZN(n373) );
  XOR2_X1 U354 ( .A(n305), .B(n373), .Z(n307) );
  XNOR2_X1 U355 ( .A(G36GAT), .B(G50GAT), .ZN(n306) );
  XNOR2_X1 U356 ( .A(n307), .B(n306), .ZN(n311) );
  XOR2_X1 U357 ( .A(KEYINPUT67), .B(KEYINPUT68), .Z(n309) );
  NAND2_X1 U358 ( .A1(G229GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U359 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U360 ( .A(n311), .B(n310), .Z(n316) );
  XOR2_X1 U361 ( .A(KEYINPUT29), .B(G197GAT), .Z(n313) );
  XNOR2_X1 U362 ( .A(G113GAT), .B(G141GAT), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U364 ( .A(n314), .B(KEYINPUT30), .ZN(n315) );
  XNOR2_X1 U365 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U366 ( .A(KEYINPUT8), .B(KEYINPUT69), .Z(n318) );
  XNOR2_X1 U367 ( .A(KEYINPUT7), .B(G43GAT), .ZN(n317) );
  XNOR2_X1 U368 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U369 ( .A(G29GAT), .B(n319), .ZN(n357) );
  XOR2_X1 U370 ( .A(n320), .B(n357), .Z(n542) );
  INV_X1 U371 ( .A(n542), .ZN(n571) );
  XNOR2_X1 U372 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n321) );
  XNOR2_X1 U373 ( .A(n321), .B(KEYINPUT70), .ZN(n366) );
  XNOR2_X1 U374 ( .A(n366), .B(n322), .ZN(n337) );
  XOR2_X1 U375 ( .A(G85GAT), .B(G99GAT), .Z(n351) );
  XOR2_X1 U376 ( .A(G120GAT), .B(G57GAT), .Z(n399) );
  XNOR2_X1 U377 ( .A(n399), .B(KEYINPUT33), .ZN(n323) );
  XNOR2_X1 U378 ( .A(n323), .B(KEYINPUT32), .ZN(n324) );
  NAND2_X1 U379 ( .A1(n351), .A2(n324), .ZN(n328) );
  INV_X1 U380 ( .A(n324), .ZN(n326) );
  INV_X1 U381 ( .A(n351), .ZN(n325) );
  NAND2_X1 U382 ( .A1(n326), .A2(n325), .ZN(n327) );
  NAND2_X1 U383 ( .A1(n328), .A2(n327), .ZN(n330) );
  AND2_X1 U384 ( .A1(G230GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U385 ( .A(n330), .B(n329), .ZN(n332) );
  INV_X1 U386 ( .A(KEYINPUT31), .ZN(n331) );
  XNOR2_X1 U387 ( .A(n332), .B(n331), .ZN(n335) );
  XNOR2_X1 U388 ( .A(G148GAT), .B(G106GAT), .ZN(n333) );
  XNOR2_X1 U389 ( .A(n333), .B(G78GAT), .ZN(n427) );
  XNOR2_X1 U390 ( .A(n427), .B(KEYINPUT71), .ZN(n334) );
  XNOR2_X1 U391 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U392 ( .A(n337), .B(n336), .ZN(n578) );
  XOR2_X1 U393 ( .A(n578), .B(KEYINPUT41), .Z(n338) );
  XNOR2_X1 U394 ( .A(KEYINPUT65), .B(n338), .ZN(n545) );
  NOR2_X1 U395 ( .A1(n571), .A2(n545), .ZN(n339) );
  XNOR2_X1 U396 ( .A(KEYINPUT46), .B(n339), .ZN(n379) );
  XOR2_X1 U397 ( .A(G92GAT), .B(G106GAT), .Z(n341) );
  XNOR2_X1 U398 ( .A(G134GAT), .B(G218GAT), .ZN(n340) );
  XNOR2_X1 U399 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U400 ( .A(KEYINPUT10), .B(KEYINPUT74), .Z(n343) );
  XNOR2_X1 U401 ( .A(KEYINPUT72), .B(KEYINPUT9), .ZN(n342) );
  XNOR2_X1 U402 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U403 ( .A(n345), .B(n344), .Z(n350) );
  XOR2_X1 U404 ( .A(KEYINPUT11), .B(KEYINPUT66), .Z(n347) );
  NAND2_X1 U405 ( .A1(G232GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U406 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U407 ( .A(KEYINPUT73), .B(n348), .ZN(n349) );
  XNOR2_X1 U408 ( .A(n350), .B(n349), .ZN(n352) );
  XOR2_X1 U409 ( .A(n352), .B(n351), .Z(n355) );
  XOR2_X1 U410 ( .A(G162GAT), .B(G50GAT), .Z(n420) );
  XNOR2_X1 U411 ( .A(n353), .B(n420), .ZN(n354) );
  XNOR2_X1 U412 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U413 ( .A(n357), .B(n356), .Z(n552) );
  XOR2_X1 U414 ( .A(KEYINPUT14), .B(KEYINPUT76), .Z(n359) );
  XNOR2_X1 U415 ( .A(KEYINPUT77), .B(KEYINPUT15), .ZN(n358) );
  XNOR2_X1 U416 ( .A(n359), .B(n358), .ZN(n377) );
  XOR2_X1 U417 ( .A(G78GAT), .B(G211GAT), .Z(n361) );
  XNOR2_X1 U418 ( .A(G155GAT), .B(G57GAT), .ZN(n360) );
  XNOR2_X1 U419 ( .A(n361), .B(n360), .ZN(n365) );
  XOR2_X1 U420 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n363) );
  XNOR2_X1 U421 ( .A(G8GAT), .B(G64GAT), .ZN(n362) );
  XNOR2_X1 U422 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U423 ( .A(n365), .B(n364), .Z(n371) );
  XOR2_X1 U424 ( .A(n366), .B(G183GAT), .Z(n369) );
  NAND2_X1 U425 ( .A1(G231GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U426 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U427 ( .A(n372), .B(KEYINPUT80), .Z(n375) );
  XNOR2_X1 U428 ( .A(n373), .B(KEYINPUT12), .ZN(n374) );
  XNOR2_X1 U429 ( .A(n375), .B(n374), .ZN(n376) );
  OR2_X1 U430 ( .A1(n552), .A2(n582), .ZN(n378) );
  NOR2_X1 U431 ( .A1(n379), .A2(n378), .ZN(n380) );
  XNOR2_X1 U432 ( .A(KEYINPUT47), .B(n380), .ZN(n388) );
  XNOR2_X1 U433 ( .A(KEYINPUT104), .B(KEYINPUT36), .ZN(n382) );
  INV_X1 U434 ( .A(n552), .ZN(n381) );
  XOR2_X1 U435 ( .A(n382), .B(n381), .Z(n584) );
  NAND2_X1 U436 ( .A1(n582), .A2(n584), .ZN(n383) );
  XNOR2_X1 U437 ( .A(KEYINPUT45), .B(n383), .ZN(n384) );
  XNOR2_X1 U438 ( .A(KEYINPUT114), .B(n385), .ZN(n386) );
  NAND2_X1 U439 ( .A1(n386), .A2(n571), .ZN(n387) );
  NAND2_X1 U440 ( .A1(n388), .A2(n387), .ZN(n391) );
  XOR2_X1 U441 ( .A(KEYINPUT115), .B(KEYINPUT48), .Z(n389) );
  AND2_X1 U442 ( .A1(n492), .A2(n539), .ZN(n393) );
  INV_X1 U443 ( .A(KEYINPUT54), .ZN(n392) );
  XNOR2_X1 U444 ( .A(n393), .B(n392), .ZN(n567) );
  XOR2_X1 U445 ( .A(KEYINPUT81), .B(G134GAT), .Z(n395) );
  XNOR2_X1 U446 ( .A(G127GAT), .B(G113GAT), .ZN(n394) );
  XNOR2_X1 U447 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U448 ( .A(KEYINPUT0), .B(n396), .Z(n445) );
  XOR2_X1 U449 ( .A(G141GAT), .B(G155GAT), .Z(n398) );
  XNOR2_X1 U450 ( .A(KEYINPUT3), .B(KEYINPUT2), .ZN(n397) );
  XNOR2_X1 U451 ( .A(n398), .B(n397), .ZN(n428) );
  XOR2_X1 U452 ( .A(n399), .B(n428), .Z(n401) );
  XNOR2_X1 U453 ( .A(G29GAT), .B(G162GAT), .ZN(n400) );
  XNOR2_X1 U454 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U455 ( .A(n445), .B(n402), .ZN(n415) );
  XOR2_X1 U456 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n404) );
  XNOR2_X1 U457 ( .A(G85GAT), .B(G148GAT), .ZN(n403) );
  XNOR2_X1 U458 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U459 ( .A(KEYINPUT91), .B(G1GAT), .Z(n406) );
  XNOR2_X1 U460 ( .A(KEYINPUT4), .B(KEYINPUT6), .ZN(n405) );
  XNOR2_X1 U461 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U462 ( .A(n408), .B(n407), .Z(n413) );
  XOR2_X1 U463 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n410) );
  NAND2_X1 U464 ( .A1(G225GAT), .A2(G233GAT), .ZN(n409) );
  XNOR2_X1 U465 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U466 ( .A(KEYINPUT90), .B(n411), .ZN(n412) );
  XNOR2_X1 U467 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U468 ( .A(n415), .B(n414), .Z(n514) );
  XOR2_X1 U469 ( .A(KEYINPUT24), .B(n416), .Z(n418) );
  NAND2_X1 U470 ( .A1(G228GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U471 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U472 ( .A(n419), .B(KEYINPUT23), .Z(n422) );
  XNOR2_X1 U473 ( .A(n420), .B(KEYINPUT87), .ZN(n421) );
  XNOR2_X1 U474 ( .A(n422), .B(n421), .ZN(n426) );
  XOR2_X1 U475 ( .A(KEYINPUT86), .B(KEYINPUT22), .Z(n424) );
  XNOR2_X1 U476 ( .A(G22GAT), .B(G204GAT), .ZN(n423) );
  XNOR2_X1 U477 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U478 ( .A(n426), .B(n425), .Z(n430) );
  XNOR2_X1 U479 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U480 ( .A(n430), .B(n429), .Z(n459) );
  NAND2_X1 U481 ( .A1(n514), .A2(n459), .ZN(n431) );
  OR2_X1 U482 ( .A1(n567), .A2(n431), .ZN(n432) );
  XNOR2_X1 U483 ( .A(n432), .B(KEYINPUT55), .ZN(n556) );
  XOR2_X1 U484 ( .A(KEYINPUT82), .B(KEYINPUT83), .Z(n434) );
  XNOR2_X1 U485 ( .A(KEYINPUT85), .B(KEYINPUT84), .ZN(n433) );
  XNOR2_X1 U486 ( .A(n434), .B(n433), .ZN(n449) );
  XOR2_X1 U487 ( .A(G169GAT), .B(G99GAT), .Z(n436) );
  XNOR2_X1 U488 ( .A(G43GAT), .B(G190GAT), .ZN(n435) );
  XNOR2_X1 U489 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U490 ( .A(KEYINPUT20), .B(G176GAT), .Z(n438) );
  XNOR2_X1 U491 ( .A(G120GAT), .B(G15GAT), .ZN(n437) );
  XNOR2_X1 U492 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U493 ( .A(n440), .B(n439), .Z(n447) );
  XOR2_X1 U494 ( .A(n441), .B(G71GAT), .Z(n443) );
  NAND2_X1 U495 ( .A1(G227GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U496 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U497 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U498 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U499 ( .A(n449), .B(n448), .ZN(n555) );
  AND2_X1 U500 ( .A1(n555), .A2(n552), .ZN(n450) );
  AND2_X1 U501 ( .A1(n556), .A2(n450), .ZN(n453) );
  NOR2_X1 U502 ( .A1(n571), .A2(n578), .ZN(n486) );
  INV_X1 U503 ( .A(n582), .ZN(n565) );
  NOR2_X1 U504 ( .A1(n552), .A2(n565), .ZN(n454) );
  XNOR2_X1 U505 ( .A(n454), .B(KEYINPUT16), .ZN(n469) );
  INV_X1 U506 ( .A(n555), .ZN(n526) );
  INV_X1 U507 ( .A(n514), .ZN(n568) );
  XOR2_X1 U508 ( .A(n516), .B(KEYINPUT27), .Z(n462) );
  NAND2_X1 U509 ( .A1(n568), .A2(n462), .ZN(n541) );
  XOR2_X1 U510 ( .A(n459), .B(KEYINPUT28), .Z(n496) );
  NOR2_X1 U511 ( .A1(n541), .A2(n496), .ZN(n524) );
  NAND2_X1 U512 ( .A1(n526), .A2(n524), .ZN(n455) );
  XNOR2_X1 U513 ( .A(n455), .B(KEYINPUT94), .ZN(n468) );
  NAND2_X1 U514 ( .A1(n492), .A2(n555), .ZN(n456) );
  XNOR2_X1 U515 ( .A(n456), .B(KEYINPUT96), .ZN(n457) );
  NAND2_X1 U516 ( .A1(n457), .A2(n459), .ZN(n458) );
  XNOR2_X1 U517 ( .A(n458), .B(KEYINPUT25), .ZN(n464) );
  NOR2_X1 U518 ( .A1(n555), .A2(n459), .ZN(n461) );
  XNOR2_X1 U519 ( .A(KEYINPUT95), .B(KEYINPUT26), .ZN(n460) );
  XOR2_X1 U520 ( .A(n461), .B(n460), .Z(n569) );
  AND2_X1 U521 ( .A1(n569), .A2(n462), .ZN(n463) );
  NOR2_X1 U522 ( .A1(n464), .A2(n463), .ZN(n465) );
  XNOR2_X1 U523 ( .A(n465), .B(KEYINPUT97), .ZN(n466) );
  NAND2_X1 U524 ( .A1(n466), .A2(n514), .ZN(n467) );
  NAND2_X1 U525 ( .A1(n468), .A2(n467), .ZN(n482) );
  NAND2_X1 U526 ( .A1(n469), .A2(n482), .ZN(n470) );
  XOR2_X1 U527 ( .A(KEYINPUT98), .B(n470), .Z(n500) );
  NAND2_X1 U528 ( .A1(n486), .A2(n500), .ZN(n478) );
  NOR2_X1 U529 ( .A1(n514), .A2(n478), .ZN(n471) );
  XOR2_X1 U530 ( .A(G1GAT), .B(n471), .Z(n472) );
  XNOR2_X1 U531 ( .A(KEYINPUT34), .B(n472), .ZN(G1324GAT) );
  NOR2_X1 U532 ( .A1(n516), .A2(n478), .ZN(n474) );
  XNOR2_X1 U533 ( .A(G8GAT), .B(KEYINPUT99), .ZN(n473) );
  XNOR2_X1 U534 ( .A(n474), .B(n473), .ZN(G1325GAT) );
  NOR2_X1 U535 ( .A1(n526), .A2(n478), .ZN(n476) );
  XNOR2_X1 U536 ( .A(KEYINPUT100), .B(KEYINPUT35), .ZN(n475) );
  XNOR2_X1 U537 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U538 ( .A(G15GAT), .B(n477), .ZN(G1326GAT) );
  INV_X1 U539 ( .A(n496), .ZN(n521) );
  NOR2_X1 U540 ( .A1(n521), .A2(n478), .ZN(n480) );
  XNOR2_X1 U541 ( .A(KEYINPUT101), .B(KEYINPUT102), .ZN(n479) );
  XNOR2_X1 U542 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U543 ( .A(G22GAT), .B(n481), .ZN(G1327GAT) );
  XNOR2_X1 U544 ( .A(G29GAT), .B(KEYINPUT103), .ZN(n491) );
  XOR2_X1 U545 ( .A(KEYINPUT106), .B(KEYINPUT38), .Z(n488) );
  NAND2_X1 U546 ( .A1(n565), .A2(n482), .ZN(n483) );
  XNOR2_X1 U547 ( .A(n483), .B(KEYINPUT105), .ZN(n484) );
  NAND2_X1 U548 ( .A1(n484), .A2(n584), .ZN(n485) );
  XNOR2_X1 U549 ( .A(KEYINPUT37), .B(n485), .ZN(n513) );
  NAND2_X1 U550 ( .A1(n486), .A2(n513), .ZN(n487) );
  XNOR2_X1 U551 ( .A(n488), .B(n487), .ZN(n497) );
  NAND2_X1 U552 ( .A1(n497), .A2(n568), .ZN(n489) );
  XNOR2_X1 U553 ( .A(n489), .B(KEYINPUT39), .ZN(n490) );
  XNOR2_X1 U554 ( .A(n491), .B(n490), .ZN(G1328GAT) );
  NAND2_X1 U555 ( .A1(n497), .A2(n492), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n493), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U557 ( .A1(n555), .A2(n497), .ZN(n494) );
  XNOR2_X1 U558 ( .A(n494), .B(KEYINPUT40), .ZN(n495) );
  XNOR2_X1 U559 ( .A(G43GAT), .B(n495), .ZN(G1330GAT) );
  XOR2_X1 U560 ( .A(G50GAT), .B(KEYINPUT107), .Z(n499) );
  NAND2_X1 U561 ( .A1(n497), .A2(n496), .ZN(n498) );
  XNOR2_X1 U562 ( .A(n499), .B(n498), .ZN(G1331GAT) );
  XNOR2_X1 U563 ( .A(KEYINPUT108), .B(n545), .ZN(n558) );
  NOR2_X1 U564 ( .A1(n558), .A2(n542), .ZN(n512) );
  NAND2_X1 U565 ( .A1(n512), .A2(n500), .ZN(n508) );
  NOR2_X1 U566 ( .A1(n514), .A2(n508), .ZN(n502) );
  XNOR2_X1 U567 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n501) );
  XNOR2_X1 U568 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(n503), .ZN(G1332GAT) );
  NOR2_X1 U570 ( .A1(n516), .A2(n508), .ZN(n504) );
  XOR2_X1 U571 ( .A(KEYINPUT110), .B(n504), .Z(n505) );
  XNOR2_X1 U572 ( .A(G64GAT), .B(n505), .ZN(G1333GAT) );
  NOR2_X1 U573 ( .A1(n526), .A2(n508), .ZN(n507) );
  XNOR2_X1 U574 ( .A(G71GAT), .B(KEYINPUT111), .ZN(n506) );
  XNOR2_X1 U575 ( .A(n507), .B(n506), .ZN(G1334GAT) );
  NOR2_X1 U576 ( .A1(n521), .A2(n508), .ZN(n510) );
  XNOR2_X1 U577 ( .A(KEYINPUT112), .B(KEYINPUT43), .ZN(n509) );
  XNOR2_X1 U578 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U579 ( .A(G78GAT), .B(n511), .ZN(G1335GAT) );
  NAND2_X1 U580 ( .A1(n513), .A2(n512), .ZN(n520) );
  NOR2_X1 U581 ( .A1(n514), .A2(n520), .ZN(n515) );
  XOR2_X1 U582 ( .A(G85GAT), .B(n515), .Z(G1336GAT) );
  NOR2_X1 U583 ( .A1(n516), .A2(n520), .ZN(n518) );
  XNOR2_X1 U584 ( .A(G92GAT), .B(KEYINPUT113), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(G1337GAT) );
  NOR2_X1 U586 ( .A1(n526), .A2(n520), .ZN(n519) );
  XOR2_X1 U587 ( .A(G99GAT), .B(n519), .Z(G1338GAT) );
  NOR2_X1 U588 ( .A1(n521), .A2(n520), .ZN(n522) );
  XOR2_X1 U589 ( .A(KEYINPUT44), .B(n522), .Z(n523) );
  XNOR2_X1 U590 ( .A(G106GAT), .B(n523), .ZN(G1339GAT) );
  NAND2_X1 U591 ( .A1(n524), .A2(n539), .ZN(n525) );
  NOR2_X1 U592 ( .A1(n526), .A2(n525), .ZN(n535) );
  NAND2_X1 U593 ( .A1(n542), .A2(n535), .ZN(n527) );
  XNOR2_X1 U594 ( .A(n527), .B(G113GAT), .ZN(G1340GAT) );
  INV_X1 U595 ( .A(n535), .ZN(n528) );
  NOR2_X1 U596 ( .A1(n558), .A2(n528), .ZN(n530) );
  XNOR2_X1 U597 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n529) );
  XNOR2_X1 U598 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U599 ( .A(G120GAT), .B(n531), .ZN(G1341GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n533) );
  NAND2_X1 U601 ( .A1(n535), .A2(n582), .ZN(n532) );
  XNOR2_X1 U602 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(n534), .ZN(G1342GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n537) );
  NAND2_X1 U605 ( .A1(n535), .A2(n552), .ZN(n536) );
  XNOR2_X1 U606 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U607 ( .A(G134GAT), .B(n538), .ZN(G1343GAT) );
  NAND2_X1 U608 ( .A1(n569), .A2(n539), .ZN(n540) );
  NOR2_X1 U609 ( .A1(n541), .A2(n540), .ZN(n551) );
  NAND2_X1 U610 ( .A1(n542), .A2(n551), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n543), .B(G141GAT), .ZN(G1344GAT) );
  INV_X1 U612 ( .A(n551), .ZN(n544) );
  NOR2_X1 U613 ( .A1(n545), .A2(n544), .ZN(n547) );
  XNOR2_X1 U614 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(n548), .ZN(G1345GAT) );
  XOR2_X1 U617 ( .A(G155GAT), .B(KEYINPUT119), .Z(n550) );
  NAND2_X1 U618 ( .A1(n551), .A2(n582), .ZN(n549) );
  XNOR2_X1 U619 ( .A(n550), .B(n549), .ZN(G1346GAT) );
  NAND2_X1 U620 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n553), .B(KEYINPUT120), .ZN(n554) );
  XNOR2_X1 U622 ( .A(G162GAT), .B(n554), .ZN(G1347GAT) );
  NAND2_X1 U623 ( .A1(n556), .A2(n555), .ZN(n564) );
  NOR2_X1 U624 ( .A1(n571), .A2(n564), .ZN(n557) );
  XOR2_X1 U625 ( .A(G169GAT), .B(n557), .Z(G1348GAT) );
  NOR2_X1 U626 ( .A1(n558), .A2(n564), .ZN(n563) );
  XOR2_X1 U627 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n560) );
  XNOR2_X1 U628 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n559) );
  XNOR2_X1 U629 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U630 ( .A(KEYINPUT121), .B(n561), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n563), .B(n562), .ZN(G1349GAT) );
  NOR2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U633 ( .A(G183GAT), .B(n566), .Z(G1350GAT) );
  NOR2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n570) );
  NAND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n577) );
  NOR2_X1 U636 ( .A1(n571), .A2(n577), .ZN(n576) );
  XOR2_X1 U637 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n573) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(KEYINPUT60), .B(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n580) );
  INV_X1 U643 ( .A(n577), .ZN(n585) );
  NAND2_X1 U644 ( .A1(n585), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XOR2_X1 U646 ( .A(G204GAT), .B(n581), .Z(G1353GAT) );
  NAND2_X1 U647 ( .A1(n585), .A2(n582), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n583), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U649 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n587) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(n588) );
  XOR2_X1 U652 ( .A(G218GAT), .B(n588), .Z(G1355GAT) );
endmodule

