

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788;

  XNOR2_X1 U372 ( .A(n423), .B(n564), .ZN(n714) );
  NOR2_X1 U373 ( .A1(n601), .A2(n620), .ZN(n587) );
  AND2_X1 U374 ( .A1(n723), .A2(n724), .ZN(n720) );
  BUF_X1 U375 ( .A(G107), .Z(n704) );
  XNOR2_X1 U376 ( .A(n456), .B(n488), .ZN(n479) );
  XOR2_X1 U377 ( .A(KEYINPUT23), .B(KEYINPUT97), .Z(n491) );
  XNOR2_X2 U378 ( .A(n392), .B(n408), .ZN(n407) );
  XNOR2_X1 U379 ( .A(n348), .B(n495), .ZN(n496) );
  XNOR2_X1 U380 ( .A(n349), .B(n493), .ZN(n348) );
  OR2_X2 U381 ( .A1(n380), .A2(n373), .ZN(n437) );
  NOR2_X4 U382 ( .A1(n643), .A2(n646), .ZN(n753) );
  XOR2_X2 U383 ( .A(n465), .B(n464), .Z(n379) );
  NOR2_X1 U384 ( .A1(G237), .A2(G953), .ZN(n508) );
  INV_X1 U385 ( .A(G953), .ZN(n780) );
  BUF_X1 U386 ( .A(G122), .Z(n663) );
  BUF_X1 U387 ( .A(G143), .Z(n654) );
  XOR2_X1 U388 ( .A(n491), .B(n490), .Z(n349) );
  AND2_X2 U389 ( .A1(n354), .A2(n430), .ZN(n429) );
  XNOR2_X1 U390 ( .A(n352), .B(n350), .ZN(n688) );
  XNOR2_X2 U391 ( .A(G119), .B(G113), .ZN(n358) );
  XNOR2_X2 U392 ( .A(G110), .B(G107), .ZN(n356) );
  XNOR2_X1 U393 ( .A(n645), .B(KEYINPUT86), .ZN(n646) );
  AND2_X1 U394 ( .A1(n440), .A2(n435), .ZN(n434) );
  AND2_X1 U395 ( .A1(n659), .A2(n658), .ZN(n574) );
  NOR2_X1 U396 ( .A1(n380), .A2(KEYINPUT89), .ZN(n433) );
  XNOR2_X1 U397 ( .A(n607), .B(n606), .ZN(n657) );
  AND2_X1 U398 ( .A1(n381), .A2(n555), .ZN(n570) );
  XNOR2_X1 U399 ( .A(n553), .B(n552), .ZN(n381) );
  NOR2_X1 U400 ( .A1(n758), .A2(n418), .ZN(n360) );
  XNOR2_X1 U401 ( .A(n769), .B(n484), .ZN(n352) );
  XNOR2_X1 U402 ( .A(n461), .B(n351), .ZN(n350) );
  XNOR2_X1 U403 ( .A(n357), .B(n356), .ZN(n770) );
  XNOR2_X1 U404 ( .A(n477), .B(n479), .ZN(n351) );
  XNOR2_X1 U405 ( .A(n770), .B(KEYINPUT75), .ZN(n484) );
  XNOR2_X2 U406 ( .A(n353), .B(n511), .ZN(n769) );
  XNOR2_X2 U407 ( .A(n455), .B(n454), .ZN(n477) );
  XNOR2_X2 U408 ( .A(n529), .B(KEYINPUT16), .ZN(n353) );
  XNOR2_X2 U409 ( .A(n358), .B(n359), .ZN(n511) );
  NAND2_X1 U410 ( .A1(n591), .A2(n431), .ZN(n354) );
  XNOR2_X2 U411 ( .A(n355), .B(n579), .ZN(n642) );
  NAND2_X1 U412 ( .A1(n578), .A2(n577), .ZN(n355) );
  XNOR2_X2 U413 ( .A(G104), .B(G101), .ZN(n357) );
  XNOR2_X2 U414 ( .A(KEYINPUT74), .B(KEYINPUT3), .ZN(n359) );
  XNOR2_X2 U415 ( .A(n425), .B(G116), .ZN(n529) );
  NAND2_X1 U416 ( .A1(n416), .A2(n360), .ZN(n361) );
  XNOR2_X2 U417 ( .A(n513), .B(KEYINPUT33), .ZN(n758) );
  XNOR2_X2 U418 ( .A(n549), .B(KEYINPUT96), .ZN(n416) );
  XNOR2_X2 U419 ( .A(n476), .B(n368), .ZN(n549) );
  NAND2_X1 U420 ( .A1(n361), .A2(n417), .ZN(n384) );
  BUF_X1 U421 ( .A(n770), .Z(n362) );
  XNOR2_X1 U422 ( .A(n378), .B(n379), .ZN(n363) );
  XNOR2_X1 U423 ( .A(n378), .B(n379), .ZN(n591) );
  XNOR2_X1 U424 ( .A(n388), .B(KEYINPUT10), .ZN(n778) );
  XNOR2_X1 U425 ( .A(G125), .B(G140), .ZN(n388) );
  XNOR2_X1 U426 ( .A(n565), .B(KEYINPUT109), .ZN(n601) );
  INV_X1 U427 ( .A(n511), .ZN(n421) );
  NOR2_X1 U428 ( .A1(n657), .A2(n788), .ZN(n419) );
  NAND2_X1 U429 ( .A1(n375), .A2(n433), .ZN(n432) );
  INV_X1 U430 ( .A(G469), .ZN(n411) );
  NAND2_X1 U431 ( .A1(G902), .A2(G469), .ZN(n413) );
  INV_X1 U432 ( .A(G146), .ZN(n488) );
  INV_X1 U433 ( .A(G128), .ZN(n454) );
  NAND2_X1 U434 ( .A1(n462), .A2(n448), .ZN(n447) );
  NAND2_X1 U435 ( .A1(KEYINPUT65), .A2(KEYINPUT2), .ZN(n448) );
  XNOR2_X1 U436 ( .A(G131), .B(KEYINPUT103), .ZN(n519) );
  XOR2_X1 U437 ( .A(G104), .B(KEYINPUT102), .Z(n520) );
  XNOR2_X1 U438 ( .A(n588), .B(n487), .ZN(n554) );
  INV_X1 U439 ( .A(n778), .ZN(n389) );
  XNOR2_X1 U440 ( .A(n778), .B(n488), .ZN(n518) );
  AND2_X1 U441 ( .A1(n407), .A2(n622), .ZN(n513) );
  XNOR2_X1 U442 ( .A(n593), .B(n393), .ZN(n757) );
  XNOR2_X1 U443 ( .A(n394), .B(KEYINPUT41), .ZN(n393) );
  INV_X1 U444 ( .A(KEYINPUT115), .ZN(n394) );
  XNOR2_X1 U445 ( .A(n605), .B(KEYINPUT39), .ZN(n405) );
  NAND2_X1 U446 ( .A1(n428), .A2(n427), .ZN(n426) );
  NOR2_X1 U447 ( .A1(n600), .A2(n431), .ZN(n427) );
  OR2_X1 U448 ( .A1(n601), .A2(KEYINPUT67), .ZN(n398) );
  AND2_X1 U449 ( .A1(n399), .A2(n555), .ZN(n385) );
  XNOR2_X1 U450 ( .A(n528), .B(n527), .ZN(n568) );
  OR2_X1 U451 ( .A1(n666), .A2(G902), .ZN(n406) );
  INV_X1 U452 ( .A(n563), .ZN(n439) );
  INV_X1 U453 ( .A(G237), .ZN(n463) );
  XNOR2_X1 U454 ( .A(KEYINPUT79), .B(KEYINPUT5), .ZN(n506) );
  XNOR2_X1 U455 ( .A(G101), .B(G116), .ZN(n507) );
  XNOR2_X1 U456 ( .A(G125), .B(KEYINPUT17), .ZN(n459) );
  NAND2_X1 U457 ( .A1(G234), .A2(G237), .ZN(n468) );
  XNOR2_X1 U458 ( .A(n387), .B(KEYINPUT107), .ZN(n738) );
  NOR2_X1 U459 ( .A1(n568), .A2(n566), .ZN(n387) );
  XNOR2_X1 U460 ( .A(n592), .B(KEYINPUT38), .ZN(n736) );
  INV_X1 U461 ( .A(KEYINPUT91), .ZN(n431) );
  NAND2_X1 U462 ( .A1(n600), .A2(n431), .ZN(n430) );
  INV_X1 U463 ( .A(n612), .ZN(n418) );
  NOR2_X1 U464 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X2 U465 ( .A1(n412), .A2(n409), .ZN(n588) );
  AND2_X1 U466 ( .A1(n414), .A2(n413), .ZN(n412) );
  NAND2_X1 U467 ( .A1(n411), .A2(n537), .ZN(n410) );
  XNOR2_X1 U468 ( .A(KEYINPUT24), .B(KEYINPUT98), .ZN(n490) );
  XNOR2_X1 U469 ( .A(G119), .B(G128), .ZN(n492) );
  INV_X1 U470 ( .A(KEYINPUT105), .ZN(n402) );
  NAND2_X1 U471 ( .A1(n449), .A2(n447), .ZN(n446) );
  NAND2_X1 U472 ( .A1(n641), .A2(KEYINPUT65), .ZN(n449) );
  INV_X1 U473 ( .A(KEYINPUT2), .ZN(n444) );
  XNOR2_X1 U474 ( .A(n526), .B(n525), .ZN(n647) );
  XNOR2_X1 U475 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U476 ( .A(G137), .B(G131), .ZN(n478) );
  XOR2_X1 U477 ( .A(G140), .B(KEYINPUT81), .Z(n482) );
  BUF_X1 U478 ( .A(n554), .Z(n719) );
  INV_X1 U479 ( .A(KEYINPUT19), .ZN(n467) );
  INV_X1 U480 ( .A(KEYINPUT6), .ZN(n391) );
  XOR2_X1 U481 ( .A(KEYINPUT62), .B(n666), .Z(n667) );
  XOR2_X1 U482 ( .A(n647), .B(KEYINPUT59), .Z(n648) );
  NAND2_X1 U483 ( .A1(n405), .A2(n403), .ZN(n607) );
  INV_X1 U484 ( .A(n619), .ZN(n403) );
  NAND2_X1 U485 ( .A1(n424), .A2(n549), .ZN(n423) );
  NAND2_X1 U486 ( .A1(n397), .A2(n395), .ZN(n659) );
  AND2_X1 U487 ( .A1(n386), .A2(n367), .ZN(n397) );
  NAND2_X1 U488 ( .A1(n396), .A2(n556), .ZN(n395) );
  NOR2_X1 U489 ( .A1(n762), .A2(G953), .ZN(n763) );
  AND2_X1 U490 ( .A1(n407), .A2(n565), .ZN(n364) );
  INV_X1 U491 ( .A(KEYINPUT65), .ZN(n451) );
  XOR2_X1 U492 ( .A(G110), .B(G137), .Z(n365) );
  NOR2_X1 U493 ( .A1(n597), .A2(n565), .ZN(n366) );
  AND2_X1 U494 ( .A1(n398), .A2(n586), .ZN(n367) );
  XOR2_X1 U495 ( .A(n475), .B(KEYINPUT0), .Z(n368) );
  INV_X1 U496 ( .A(n715), .ZN(n404) );
  XNOR2_X1 U497 ( .A(G902), .B(KEYINPUT15), .ZN(n641) );
  XOR2_X1 U498 ( .A(n608), .B(KEYINPUT46), .Z(n369) );
  AND2_X1 U499 ( .A1(n462), .A2(KEYINPUT65), .ZN(n370) );
  NAND2_X1 U500 ( .A1(n451), .A2(n444), .ZN(n371) );
  AND2_X1 U501 ( .A1(n563), .A2(KEYINPUT89), .ZN(n372) );
  AND2_X1 U502 ( .A1(n439), .A2(n438), .ZN(n373) );
  INV_X1 U503 ( .A(KEYINPUT89), .ZN(n438) );
  XNOR2_X1 U504 ( .A(n689), .B(n690), .ZN(n691) );
  NAND2_X1 U505 ( .A1(n445), .A2(n443), .ZN(n374) );
  NAND2_X1 U506 ( .A1(n445), .A2(n443), .ZN(n450) );
  OR2_X1 U507 ( .A1(n750), .A2(n371), .ZN(n443) );
  NOR2_X2 U508 ( .A1(n753), .A2(n374), .ZN(n687) );
  AND2_X1 U509 ( .A1(n562), .A2(n574), .ZN(n375) );
  NOR2_X2 U510 ( .A1(n753), .A2(n450), .ZN(n376) );
  NOR2_X1 U511 ( .A1(n753), .A2(n374), .ZN(n377) );
  XNOR2_X1 U512 ( .A(n420), .B(n390), .ZN(n666) );
  XNOR2_X1 U513 ( .A(n623), .B(n467), .ZN(n609) );
  NAND2_X1 U514 ( .A1(n429), .A2(n426), .ZN(n623) );
  BUF_X1 U515 ( .A(n363), .Z(n592) );
  NAND2_X1 U516 ( .A1(n714), .A2(n700), .ZN(n422) );
  XNOR2_X1 U517 ( .A(n565), .B(n391), .ZN(n622) );
  NOR2_X2 U518 ( .A1(n688), .A2(n462), .ZN(n378) );
  NAND2_X1 U519 ( .A1(n612), .A2(n514), .ZN(n417) );
  NAND2_X1 U520 ( .A1(n380), .A2(n438), .ZN(n436) );
  NAND2_X1 U521 ( .A1(n571), .A2(n698), .ZN(n380) );
  NAND2_X1 U522 ( .A1(n381), .A2(n453), .ZN(n561) );
  NAND2_X1 U523 ( .A1(n381), .A2(n385), .ZN(n386) );
  XNOR2_X2 U524 ( .A(n382), .B(n542), .ZN(n661) );
  NAND2_X1 U525 ( .A1(n384), .A2(n383), .ZN(n382) );
  NAND2_X1 U526 ( .A1(n415), .A2(n416), .ZN(n383) );
  NOR2_X1 U527 ( .A1(n738), .A2(n547), .ZN(n548) );
  XNOR2_X1 U528 ( .A(n485), .B(n390), .ZN(n682) );
  XNOR2_X1 U529 ( .A(n390), .B(n389), .ZN(n782) );
  XNOR2_X2 U530 ( .A(n535), .B(n480), .ZN(n390) );
  INV_X1 U531 ( .A(n565), .ZN(n726) );
  NAND2_X1 U532 ( .A1(n554), .A2(n720), .ZN(n392) );
  NAND2_X1 U533 ( .A1(n416), .A2(n366), .ZN(n700) );
  INV_X1 U534 ( .A(n570), .ZN(n396) );
  AND2_X1 U535 ( .A1(n601), .A2(KEYINPUT67), .ZN(n399) );
  XNOR2_X1 U536 ( .A(n400), .B(n531), .ZN(n536) );
  XNOR2_X1 U537 ( .A(n534), .B(n401), .ZN(n400) );
  XNOR2_X1 U538 ( .A(n529), .B(n402), .ZN(n401) );
  NAND2_X1 U539 ( .A1(n405), .A2(n404), .ZN(n656) );
  XNOR2_X2 U540 ( .A(n406), .B(G472), .ZN(n565) );
  INV_X1 U541 ( .A(KEYINPUT78), .ZN(n408) );
  NAND2_X1 U542 ( .A1(n682), .A2(G469), .ZN(n414) );
  OR2_X1 U543 ( .A1(n682), .A2(n410), .ZN(n409) );
  NOR2_X1 U544 ( .A1(n758), .A2(KEYINPUT34), .ZN(n415) );
  XNOR2_X1 U545 ( .A(n419), .B(n369), .ZN(n632) );
  XNOR2_X1 U546 ( .A(n512), .B(n421), .ZN(n420) );
  INV_X2 U547 ( .A(G122), .ZN(n425) );
  NAND2_X1 U548 ( .A1(n422), .A2(n739), .ZN(n571) );
  INV_X1 U549 ( .A(n731), .ZN(n424) );
  XNOR2_X2 U550 ( .A(KEYINPUT72), .B(KEYINPUT4), .ZN(n456) );
  XNOR2_X2 U551 ( .A(n477), .B(G134), .ZN(n535) );
  INV_X1 U552 ( .A(n363), .ZN(n428) );
  NAND2_X1 U553 ( .A1(n434), .A2(n432), .ZN(n578) );
  NAND2_X1 U554 ( .A1(n437), .A2(n436), .ZN(n435) );
  NAND2_X1 U555 ( .A1(n441), .A2(n372), .ZN(n440) );
  NAND2_X1 U556 ( .A1(n562), .A2(n574), .ZN(n441) );
  AND2_X2 U557 ( .A1(n442), .A2(n446), .ZN(n445) );
  NAND2_X1 U558 ( .A1(n750), .A2(n370), .ZN(n442) );
  BUF_X1 U559 ( .A(n769), .Z(n772) );
  XOR2_X1 U560 ( .A(KEYINPUT113), .B(KEYINPUT30), .Z(n452) );
  XOR2_X1 U561 ( .A(n559), .B(n558), .Z(n453) );
  INV_X1 U562 ( .A(KEYINPUT35), .ZN(n542) );
  INV_X1 U563 ( .A(KEYINPUT60), .ZN(n652) );
  XNOR2_X2 U564 ( .A(KEYINPUT64), .B(G143), .ZN(n455) );
  XNOR2_X1 U565 ( .A(KEYINPUT82), .B(KEYINPUT18), .ZN(n458) );
  NAND2_X1 U566 ( .A1(n780), .A2(G224), .ZN(n457) );
  XNOR2_X1 U567 ( .A(n458), .B(n457), .ZN(n460) );
  XNOR2_X1 U568 ( .A(n460), .B(n459), .ZN(n461) );
  INV_X1 U569 ( .A(n641), .ZN(n462) );
  INV_X1 U570 ( .A(G902), .ZN(n537) );
  NAND2_X1 U571 ( .A1(n537), .A2(n463), .ZN(n466) );
  NAND2_X1 U572 ( .A1(n466), .A2(G210), .ZN(n465) );
  INV_X1 U573 ( .A(KEYINPUT93), .ZN(n464) );
  AND2_X1 U574 ( .A1(n466), .A2(G214), .ZN(n600) );
  XOR2_X1 U575 ( .A(KEYINPUT77), .B(KEYINPUT14), .Z(n469) );
  XNOR2_X1 U576 ( .A(n469), .B(n468), .ZN(n472) );
  NAND2_X1 U577 ( .A1(n472), .A2(G952), .ZN(n470) );
  XNOR2_X1 U578 ( .A(n470), .B(KEYINPUT94), .ZN(n749) );
  INV_X1 U579 ( .A(n749), .ZN(n471) );
  NAND2_X1 U580 ( .A1(n471), .A2(n780), .ZN(n583) );
  NAND2_X1 U581 ( .A1(G902), .A2(n472), .ZN(n580) );
  XNOR2_X1 U582 ( .A(G898), .B(KEYINPUT95), .ZN(n766) );
  NAND2_X1 U583 ( .A1(G953), .A2(n766), .ZN(n774) );
  OR2_X1 U584 ( .A1(n580), .A2(n774), .ZN(n473) );
  AND2_X1 U585 ( .A1(n583), .A2(n473), .ZN(n474) );
  NOR2_X2 U586 ( .A1(n609), .A2(n474), .ZN(n476) );
  INV_X1 U587 ( .A(KEYINPUT70), .ZN(n475) );
  XNOR2_X1 U588 ( .A(n479), .B(n478), .ZN(n480) );
  NAND2_X1 U589 ( .A1(G227), .A2(n780), .ZN(n481) );
  XNOR2_X1 U590 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U591 ( .A(n484), .B(n483), .ZN(n485) );
  INV_X1 U592 ( .A(KEYINPUT69), .ZN(n486) );
  XNOR2_X1 U593 ( .A(n486), .B(KEYINPUT1), .ZN(n487) );
  NAND2_X1 U594 ( .A1(G234), .A2(n780), .ZN(n489) );
  XOR2_X1 U595 ( .A(KEYINPUT8), .B(n489), .Z(n530) );
  NAND2_X1 U596 ( .A1(G221), .A2(n530), .ZN(n495) );
  XNOR2_X1 U597 ( .A(n365), .B(n492), .ZN(n493) );
  XNOR2_X1 U598 ( .A(n518), .B(n496), .ZN(n672) );
  NAND2_X1 U599 ( .A1(n672), .A2(n537), .ZN(n501) );
  NAND2_X1 U600 ( .A1(G234), .A2(n641), .ZN(n497) );
  XNOR2_X1 U601 ( .A(KEYINPUT20), .B(n497), .ZN(n502) );
  NAND2_X1 U602 ( .A1(G217), .A2(n502), .ZN(n499) );
  INV_X1 U603 ( .A(KEYINPUT25), .ZN(n498) );
  XNOR2_X1 U604 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X2 U605 ( .A(n501), .B(n500), .ZN(n723) );
  XOR2_X1 U606 ( .A(KEYINPUT100), .B(KEYINPUT21), .Z(n504) );
  NAND2_X1 U607 ( .A1(G221), .A2(n502), .ZN(n503) );
  XNOR2_X1 U608 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U609 ( .A(KEYINPUT99), .B(n505), .ZN(n547) );
  INV_X1 U610 ( .A(n547), .ZN(n724) );
  XNOR2_X1 U611 ( .A(n507), .B(n506), .ZN(n510) );
  XNOR2_X1 U612 ( .A(KEYINPUT80), .B(n508), .ZN(n522) );
  NAND2_X1 U613 ( .A1(n522), .A2(G210), .ZN(n509) );
  XNOR2_X1 U614 ( .A(n510), .B(n509), .ZN(n512) );
  INV_X1 U615 ( .A(KEYINPUT34), .ZN(n514) );
  XOR2_X1 U616 ( .A(KEYINPUT11), .B(n663), .Z(n516) );
  XNOR2_X1 U617 ( .A(G113), .B(n654), .ZN(n515) );
  XNOR2_X1 U618 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U619 ( .A(n518), .B(n517), .ZN(n526) );
  XNOR2_X1 U620 ( .A(n520), .B(n519), .ZN(n521) );
  XOR2_X1 U621 ( .A(n521), .B(KEYINPUT12), .Z(n524) );
  AND2_X1 U622 ( .A1(n522), .A2(G214), .ZN(n523) );
  NAND2_X1 U623 ( .A1(n647), .A2(n537), .ZN(n528) );
  XOR2_X1 U624 ( .A(KEYINPUT13), .B(G475), .Z(n527) );
  NAND2_X1 U625 ( .A1(G217), .A2(n530), .ZN(n531) );
  XOR2_X1 U626 ( .A(KEYINPUT104), .B(KEYINPUT9), .Z(n533) );
  XNOR2_X1 U627 ( .A(n704), .B(KEYINPUT7), .ZN(n532) );
  XNOR2_X1 U628 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U629 ( .A(n536), .B(n535), .ZN(n677) );
  NAND2_X1 U630 ( .A1(n677), .A2(n537), .ZN(n539) );
  XNOR2_X1 U631 ( .A(KEYINPUT106), .B(G478), .ZN(n538) );
  XNOR2_X1 U632 ( .A(n539), .B(n538), .ZN(n566) );
  NAND2_X1 U633 ( .A1(n568), .A2(n566), .ZN(n541) );
  INV_X1 U634 ( .A(KEYINPUT110), .ZN(n540) );
  XNOR2_X1 U635 ( .A(n541), .B(n540), .ZN(n612) );
  INV_X1 U636 ( .A(n661), .ZN(n544) );
  INV_X1 U637 ( .A(KEYINPUT44), .ZN(n572) );
  NOR2_X1 U638 ( .A1(n572), .A2(KEYINPUT90), .ZN(n543) );
  NAND2_X1 U639 ( .A1(n544), .A2(n543), .ZN(n546) );
  NAND2_X1 U640 ( .A1(n661), .A2(KEYINPUT90), .ZN(n545) );
  NAND2_X1 U641 ( .A1(n546), .A2(n545), .ZN(n562) );
  XNOR2_X1 U642 ( .A(n548), .B(KEYINPUT108), .ZN(n550) );
  NAND2_X1 U643 ( .A1(n549), .A2(n550), .ZN(n553) );
  INV_X1 U644 ( .A(KEYINPUT68), .ZN(n551) );
  XNOR2_X1 U645 ( .A(n551), .B(KEYINPUT22), .ZN(n552) );
  INV_X1 U646 ( .A(n719), .ZN(n555) );
  INV_X1 U647 ( .A(KEYINPUT67), .ZN(n556) );
  NOR2_X1 U648 ( .A1(n622), .A2(n723), .ZN(n557) );
  NAND2_X1 U649 ( .A1(n557), .A2(n719), .ZN(n559) );
  INV_X1 U650 ( .A(KEYINPUT83), .ZN(n558) );
  XNOR2_X1 U651 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n560) );
  XNOR2_X1 U652 ( .A(n561), .B(n560), .ZN(n658) );
  NAND2_X1 U653 ( .A1(n572), .A2(KEYINPUT90), .ZN(n563) );
  XNOR2_X1 U654 ( .A(n364), .B(KEYINPUT101), .ZN(n731) );
  INV_X1 U655 ( .A(KEYINPUT31), .ZN(n564) );
  NAND2_X1 U656 ( .A1(n720), .A2(n588), .ZN(n597) );
  INV_X1 U657 ( .A(n566), .ZN(n567) );
  NAND2_X1 U658 ( .A1(n568), .A2(n567), .ZN(n619) );
  OR2_X1 U659 ( .A1(n568), .A2(n567), .ZN(n715) );
  NAND2_X1 U660 ( .A1(n619), .A2(n715), .ZN(n739) );
  INV_X1 U661 ( .A(n723), .ZN(n586) );
  NOR2_X1 U662 ( .A1(n622), .A2(n586), .ZN(n569) );
  NAND2_X1 U663 ( .A1(n570), .A2(n569), .ZN(n698) );
  NAND2_X1 U664 ( .A1(n661), .A2(n572), .ZN(n573) );
  XNOR2_X1 U665 ( .A(n573), .B(KEYINPUT71), .ZN(n575) );
  NAND2_X1 U666 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U667 ( .A(n576), .B(KEYINPUT76), .ZN(n577) );
  INV_X1 U668 ( .A(KEYINPUT45), .ZN(n579) );
  NOR2_X1 U669 ( .A1(G900), .A2(n580), .ZN(n581) );
  NAND2_X1 U670 ( .A1(n581), .A2(G953), .ZN(n582) );
  NAND2_X1 U671 ( .A1(n583), .A2(n582), .ZN(n598) );
  NAND2_X1 U672 ( .A1(n724), .A2(n598), .ZN(n584) );
  XNOR2_X1 U673 ( .A(KEYINPUT73), .B(n584), .ZN(n585) );
  NAND2_X1 U674 ( .A1(n586), .A2(n585), .ZN(n620) );
  XNOR2_X1 U675 ( .A(n587), .B(KEYINPUT28), .ZN(n589) );
  NAND2_X1 U676 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U677 ( .A(n590), .B(KEYINPUT114), .ZN(n611) );
  INV_X1 U678 ( .A(n600), .ZN(n735) );
  NAND2_X1 U679 ( .A1(n736), .A2(n735), .ZN(n740) );
  NOR2_X1 U680 ( .A1(n738), .A2(n740), .ZN(n593) );
  NOR2_X1 U681 ( .A1(n611), .A2(n757), .ZN(n595) );
  XNOR2_X1 U682 ( .A(KEYINPUT116), .B(KEYINPUT42), .ZN(n594) );
  XNOR2_X1 U683 ( .A(n595), .B(n594), .ZN(n788) );
  INV_X1 U684 ( .A(KEYINPUT112), .ZN(n596) );
  XNOR2_X1 U685 ( .A(n597), .B(n596), .ZN(n599) );
  AND2_X1 U686 ( .A1(n599), .A2(n598), .ZN(n604) );
  XNOR2_X1 U687 ( .A(n602), .B(n452), .ZN(n603) );
  AND2_X1 U688 ( .A1(n604), .A2(n603), .ZN(n614) );
  NAND2_X1 U689 ( .A1(n614), .A2(n736), .ZN(n605) );
  INV_X1 U690 ( .A(KEYINPUT40), .ZN(n606) );
  INV_X1 U691 ( .A(KEYINPUT88), .ZN(n608) );
  BUF_X1 U692 ( .A(n609), .Z(n610) );
  NOR2_X1 U693 ( .A1(n611), .A2(n610), .ZN(n709) );
  NAND2_X1 U694 ( .A1(n709), .A2(n739), .ZN(n617) );
  NAND2_X1 U695 ( .A1(n617), .A2(KEYINPUT47), .ZN(n615) );
  AND2_X1 U696 ( .A1(n612), .A2(n428), .ZN(n613) );
  NAND2_X1 U697 ( .A1(n614), .A2(n613), .ZN(n655) );
  NAND2_X1 U698 ( .A1(n615), .A2(n655), .ZN(n616) );
  XNOR2_X1 U699 ( .A(n616), .B(KEYINPUT85), .ZN(n630) );
  OR2_X1 U700 ( .A1(n617), .A2(KEYINPUT47), .ZN(n628) );
  INV_X1 U701 ( .A(KEYINPUT111), .ZN(n618) );
  XNOR2_X1 U702 ( .A(n619), .B(n618), .ZN(n712) );
  NOR2_X1 U703 ( .A1(n620), .A2(n712), .ZN(n621) );
  NAND2_X1 U704 ( .A1(n622), .A2(n621), .ZN(n635) );
  OR2_X1 U705 ( .A1(n623), .A2(n635), .ZN(n625) );
  INV_X1 U706 ( .A(KEYINPUT36), .ZN(n624) );
  XNOR2_X1 U707 ( .A(n625), .B(n624), .ZN(n626) );
  AND2_X1 U708 ( .A1(n626), .A2(n719), .ZN(n717) );
  INV_X1 U709 ( .A(n717), .ZN(n627) );
  AND2_X1 U710 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U711 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U712 ( .A1(n632), .A2(n631), .ZN(n634) );
  INV_X1 U713 ( .A(KEYINPUT48), .ZN(n633) );
  XNOR2_X1 U714 ( .A(n634), .B(n633), .ZN(n640) );
  NOR2_X1 U715 ( .A1(n719), .A2(n635), .ZN(n636) );
  NAND2_X1 U716 ( .A1(n735), .A2(n636), .ZN(n637) );
  XNOR2_X1 U717 ( .A(n637), .B(KEYINPUT43), .ZN(n638) );
  NAND2_X1 U718 ( .A1(n592), .A2(n638), .ZN(n660) );
  AND2_X1 U719 ( .A1(n656), .A2(n660), .ZN(n639) );
  NAND2_X1 U720 ( .A1(n640), .A2(n639), .ZN(n779) );
  NOR2_X2 U721 ( .A1(n642), .A2(n779), .ZN(n750) );
  BUF_X1 U722 ( .A(n642), .Z(n643) );
  INV_X1 U723 ( .A(n779), .ZN(n644) );
  NAND2_X1 U724 ( .A1(n644), .A2(KEYINPUT2), .ZN(n645) );
  NAND2_X1 U725 ( .A1(n376), .A2(G475), .ZN(n649) );
  XNOR2_X1 U726 ( .A(n649), .B(n648), .ZN(n651) );
  INV_X1 U727 ( .A(G952), .ZN(n650) );
  NAND2_X1 U728 ( .A1(n650), .A2(G953), .ZN(n693) );
  NAND2_X1 U729 ( .A1(n651), .A2(n693), .ZN(n653) );
  XNOR2_X1 U730 ( .A(n653), .B(n652), .ZN(G60) );
  XNOR2_X1 U731 ( .A(n655), .B(n654), .ZN(G45) );
  XNOR2_X1 U732 ( .A(n656), .B(G134), .ZN(G36) );
  XOR2_X1 U733 ( .A(G131), .B(n657), .Z(G33) );
  XNOR2_X1 U734 ( .A(n658), .B(G119), .ZN(G21) );
  XNOR2_X1 U735 ( .A(n659), .B(G110), .ZN(G12) );
  XNOR2_X1 U736 ( .A(n660), .B(G140), .ZN(G42) );
  BUF_X1 U737 ( .A(n661), .Z(n662) );
  INV_X1 U738 ( .A(n662), .ZN(n665) );
  INV_X1 U739 ( .A(n663), .ZN(n664) );
  XNOR2_X1 U740 ( .A(n665), .B(n664), .ZN(G24) );
  NAND2_X1 U741 ( .A1(n687), .A2(G472), .ZN(n668) );
  XNOR2_X1 U742 ( .A(n668), .B(n667), .ZN(n669) );
  NAND2_X1 U743 ( .A1(n669), .A2(n693), .ZN(n671) );
  XNOR2_X1 U744 ( .A(KEYINPUT92), .B(KEYINPUT63), .ZN(n670) );
  XNOR2_X1 U745 ( .A(n671), .B(n670), .ZN(G57) );
  BUF_X1 U746 ( .A(n687), .Z(n679) );
  NAND2_X1 U747 ( .A1(n679), .A2(G217), .ZN(n674) );
  XOR2_X1 U748 ( .A(KEYINPUT124), .B(n672), .Z(n673) );
  XNOR2_X1 U749 ( .A(n674), .B(n673), .ZN(n675) );
  INV_X1 U750 ( .A(n693), .ZN(n685) );
  NOR2_X1 U751 ( .A1(n675), .A2(n685), .ZN(G66) );
  NAND2_X1 U752 ( .A1(n376), .A2(G478), .ZN(n676) );
  XOR2_X1 U753 ( .A(n677), .B(n676), .Z(n678) );
  NOR2_X1 U754 ( .A1(n678), .A2(n685), .ZN(G63) );
  NAND2_X1 U755 ( .A1(n679), .A2(G469), .ZN(n684) );
  XNOR2_X1 U756 ( .A(KEYINPUT123), .B(KEYINPUT57), .ZN(n680) );
  XNOR2_X1 U757 ( .A(n680), .B(KEYINPUT58), .ZN(n681) );
  XNOR2_X1 U758 ( .A(n682), .B(n681), .ZN(n683) );
  XNOR2_X1 U759 ( .A(n684), .B(n683), .ZN(n686) );
  NOR2_X1 U760 ( .A1(n686), .A2(n685), .ZN(G54) );
  NAND2_X1 U761 ( .A1(n377), .A2(G210), .ZN(n692) );
  BUF_X1 U762 ( .A(n688), .Z(n689) );
  XNOR2_X1 U763 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n690) );
  XNOR2_X1 U764 ( .A(n692), .B(n691), .ZN(n694) );
  NAND2_X1 U765 ( .A1(n694), .A2(n693), .ZN(n696) );
  XNOR2_X1 U766 ( .A(KEYINPUT87), .B(KEYINPUT56), .ZN(n695) );
  XNOR2_X1 U767 ( .A(n696), .B(n695), .ZN(G51) );
  XOR2_X1 U768 ( .A(G101), .B(KEYINPUT117), .Z(n697) );
  XNOR2_X1 U769 ( .A(n698), .B(n697), .ZN(G3) );
  NOR2_X1 U770 ( .A1(n700), .A2(n712), .ZN(n699) );
  XOR2_X1 U771 ( .A(G104), .B(n699), .Z(G6) );
  NOR2_X1 U772 ( .A1(n700), .A2(n715), .ZN(n702) );
  XNOR2_X1 U773 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n701) );
  XNOR2_X1 U774 ( .A(n702), .B(n701), .ZN(n703) );
  XNOR2_X1 U775 ( .A(n704), .B(n703), .ZN(G9) );
  XOR2_X1 U776 ( .A(KEYINPUT118), .B(KEYINPUT29), .Z(n706) );
  NAND2_X1 U777 ( .A1(n709), .A2(n404), .ZN(n705) );
  XNOR2_X1 U778 ( .A(n706), .B(n705), .ZN(n707) );
  XNOR2_X1 U779 ( .A(G128), .B(n707), .ZN(G30) );
  XOR2_X1 U780 ( .A(G146), .B(KEYINPUT119), .Z(n711) );
  INV_X1 U781 ( .A(n712), .ZN(n708) );
  NAND2_X1 U782 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U783 ( .A(n711), .B(n710), .ZN(G48) );
  NOR2_X1 U784 ( .A1(n714), .A2(n712), .ZN(n713) );
  XOR2_X1 U785 ( .A(G113), .B(n713), .Z(G15) );
  NOR2_X1 U786 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U787 ( .A(G116), .B(n716), .Z(G18) );
  XNOR2_X1 U788 ( .A(G125), .B(n717), .ZN(n718) );
  XNOR2_X1 U789 ( .A(n718), .B(KEYINPUT37), .ZN(G27) );
  NOR2_X1 U790 ( .A1(n720), .A2(n719), .ZN(n722) );
  XNOR2_X1 U791 ( .A(KEYINPUT50), .B(KEYINPUT120), .ZN(n721) );
  XNOR2_X1 U792 ( .A(n722), .B(n721), .ZN(n729) );
  NOR2_X1 U793 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U794 ( .A(KEYINPUT49), .B(n725), .ZN(n727) );
  NAND2_X1 U795 ( .A1(n727), .A2(n726), .ZN(n728) );
  OR2_X1 U796 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U797 ( .A1(n731), .A2(n730), .ZN(n733) );
  XOR2_X1 U798 ( .A(KEYINPUT51), .B(KEYINPUT121), .Z(n732) );
  XNOR2_X1 U799 ( .A(n733), .B(n732), .ZN(n734) );
  NOR2_X1 U800 ( .A1(n734), .A2(n757), .ZN(n746) );
  NOR2_X1 U801 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X1 U802 ( .A1(n738), .A2(n737), .ZN(n743) );
  INV_X1 U803 ( .A(n739), .ZN(n741) );
  NOR2_X1 U804 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U805 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U806 ( .A1(n744), .A2(n758), .ZN(n745) );
  NOR2_X1 U807 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U808 ( .A(n747), .B(KEYINPUT52), .ZN(n748) );
  NOR2_X1 U809 ( .A1(n749), .A2(n748), .ZN(n756) );
  BUF_X1 U810 ( .A(n750), .Z(n752) );
  XNOR2_X1 U811 ( .A(KEYINPUT84), .B(KEYINPUT2), .ZN(n751) );
  NOR2_X1 U812 ( .A1(n752), .A2(n751), .ZN(n754) );
  NOR2_X1 U813 ( .A1(n754), .A2(n753), .ZN(n755) );
  NOR2_X1 U814 ( .A1(n756), .A2(n755), .ZN(n761) );
  NOR2_X1 U815 ( .A1(n758), .A2(n757), .ZN(n759) );
  XOR2_X1 U816 ( .A(KEYINPUT122), .B(n759), .Z(n760) );
  NAND2_X1 U817 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U818 ( .A(n763), .B(KEYINPUT53), .ZN(G75) );
  NOR2_X1 U819 ( .A1(n643), .A2(G953), .ZN(n768) );
  NAND2_X1 U820 ( .A1(G953), .A2(G224), .ZN(n764) );
  XOR2_X1 U821 ( .A(KEYINPUT61), .B(n764), .Z(n765) );
  NOR2_X1 U822 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U823 ( .A1(n768), .A2(n767), .ZN(n776) );
  XOR2_X1 U824 ( .A(KEYINPUT125), .B(n362), .Z(n771) );
  XNOR2_X1 U825 ( .A(n772), .B(n771), .ZN(n773) );
  NAND2_X1 U826 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U827 ( .A(n776), .B(n775), .ZN(n777) );
  XNOR2_X1 U828 ( .A(KEYINPUT126), .B(n777), .ZN(G69) );
  XNOR2_X1 U829 ( .A(n779), .B(n782), .ZN(n781) );
  NAND2_X1 U830 ( .A1(n781), .A2(n780), .ZN(n786) );
  XNOR2_X1 U831 ( .A(n782), .B(G227), .ZN(n783) );
  NAND2_X1 U832 ( .A1(n783), .A2(G900), .ZN(n784) );
  NAND2_X1 U833 ( .A1(n784), .A2(G953), .ZN(n785) );
  NAND2_X1 U834 ( .A1(n786), .A2(n785), .ZN(n787) );
  XOR2_X1 U835 ( .A(KEYINPUT127), .B(n787), .Z(G72) );
  XOR2_X1 U836 ( .A(n788), .B(G137), .Z(G39) );
endmodule

