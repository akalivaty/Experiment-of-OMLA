//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 1 1 0 1 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 0 0 0 0 1 1 0 0 0 1 0 0 0 1 1 0 1 0 0 1 1 0 0 0 1 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1272, new_n1273,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT64), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G68), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n217));
  INV_X1    g0017(.A(G77), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  INV_X1    g0019(.A(G107), .ZN(new_n220));
  INV_X1    g0020(.A(G264), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n206), .B1(new_n216), .B2(new_n222), .ZN(new_n223));
  OR2_X1    g0023(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT65), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(new_n204), .ZN(new_n227));
  OAI21_X1  g0027(.A(G50), .B1(G58), .B2(G68), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI22_X1  g0029(.A1(new_n223), .A2(KEYINPUT1), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  AND3_X1   g0030(.A1(new_n210), .A2(new_n225), .A3(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n234), .B(new_n235), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  NAND3_X1  g0047(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n226), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT8), .B(G58), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n203), .A2(G20), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OAI22_X1  g0057(.A1(new_n253), .A2(new_n257), .B1(new_n255), .B2(new_n248), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(G1), .A2(G13), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G41), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G223), .A2(G1698), .ZN(new_n263));
  INV_X1    g0063(.A(G226), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n263), .B1(new_n264), .B2(G1698), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT3), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n265), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G87), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n262), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT79), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G274), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n276), .B1(new_n260), .B2(new_n261), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n262), .A2(G232), .A3(new_n278), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(G190), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n265), .A2(new_n270), .B1(G33), .B2(G87), .ZN(new_n284));
  OAI21_X1  g0084(.A(KEYINPUT79), .B1(new_n284), .B2(new_n262), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n275), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G200), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n287), .B1(new_n273), .B2(new_n282), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  AND2_X1   g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  NOR2_X1   g0090(.A1(KEYINPUT3), .A2(G33), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n293));
  OAI21_X1  g0093(.A(KEYINPUT66), .B1(new_n290), .B2(new_n291), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT66), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n268), .A2(new_n295), .A3(new_n269), .ZN(new_n296));
  AOI21_X1  g0096(.A(G20), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n293), .B1(new_n297), .B2(KEYINPUT7), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G68), .ZN(new_n299));
  NAND2_X1  g0099(.A1(G58), .A2(G68), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT78), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT78), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n302), .A2(G58), .A3(G68), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n301), .B(new_n303), .C1(G58), .C2(G68), .ZN(new_n304));
  NOR2_X1   g0104(.A1(G20), .A2(G33), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n304), .A2(G20), .B1(G159), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(KEYINPUT16), .B1(new_n299), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT7), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n308), .B1(new_n270), .B2(G20), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n293), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G68), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n311), .A2(KEYINPUT16), .A3(new_n306), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n251), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n259), .B(new_n289), .C1(new_n307), .C2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT17), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n304), .A2(G20), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n305), .A2(G159), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n319), .B1(new_n298), .B2(G68), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n251), .B(new_n312), .C1(new_n320), .C2(KEYINPUT16), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n321), .A2(KEYINPUT17), .A3(new_n259), .A4(new_n289), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n316), .A2(KEYINPUT80), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NOR3_X1   g0124(.A1(new_n270), .A2(new_n308), .A3(G20), .ZN(new_n325));
  NOR3_X1   g0125(.A1(new_n290), .A2(new_n291), .A3(KEYINPUT66), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n295), .B1(new_n268), .B2(new_n269), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n204), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n325), .B1(new_n328), .B2(new_n308), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n306), .B1(new_n329), .B2(new_n212), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT16), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n251), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n319), .B1(G68), .B2(new_n310), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n333), .B1(new_n334), .B2(KEYINPUT16), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n258), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  XOR2_X1   g0136(.A(KEYINPUT68), .B(G179), .Z(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n282), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n275), .A2(new_n339), .A3(new_n285), .ZN(new_n340));
  INV_X1    g0140(.A(G169), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(new_n273), .B2(new_n282), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(KEYINPUT18), .B1(new_n336), .B2(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n343), .B1(new_n321), .B2(new_n259), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT18), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(KEYINPUT80), .B1(new_n316), .B2(new_n322), .ZN(new_n349));
  NOR3_X1   g0149(.A1(new_n324), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n262), .A2(new_n278), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n280), .B1(new_n351), .B2(new_n213), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT13), .ZN(new_n354));
  NOR2_X1   g0154(.A1(G226), .A2(G1698), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n355), .B1(new_n233), .B2(G1698), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n294), .A2(new_n356), .A3(new_n296), .ZN(new_n357));
  NAND2_X1  g0157(.A1(G33), .A2(G97), .ZN(new_n358));
  AND2_X1   g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n353), .B(new_n354), .C1(new_n359), .C2(new_n262), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n262), .B1(new_n357), .B2(new_n358), .ZN(new_n361));
  OAI21_X1  g0161(.A(KEYINPUT13), .B1(new_n361), .B2(new_n352), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G179), .ZN(new_n364));
  OAI21_X1  g0164(.A(KEYINPUT77), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n341), .B1(new_n360), .B2(new_n362), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT14), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n366), .A2(KEYINPUT77), .A3(new_n367), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT76), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT14), .B1(new_n366), .B2(new_n371), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n366), .A2(new_n371), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n369), .B(new_n370), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n267), .A2(G20), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G77), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n212), .A2(G20), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n305), .A2(G50), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n251), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT11), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT11), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n379), .A2(new_n382), .A3(new_n251), .ZN(new_n383));
  INV_X1    g0183(.A(G13), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n384), .A2(G1), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT71), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(new_n386), .A3(G20), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n248), .A2(KEYINPUT71), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT12), .B1(new_n389), .B2(G68), .ZN(new_n390));
  OR4_X1    g0190(.A1(KEYINPUT12), .A2(new_n377), .A3(G1), .A4(new_n384), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n381), .A2(new_n383), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT72), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(new_n389), .B2(new_n333), .ZN(new_n394));
  AOI211_X1 g0194(.A(KEYINPUT72), .B(new_n251), .C1(new_n387), .C2(new_n388), .ZN(new_n395));
  OAI211_X1 g0195(.A(G68), .B(new_n256), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  AND2_X1   g0196(.A1(new_n392), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n374), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G190), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n397), .B1(new_n400), .B2(new_n363), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n287), .B1(new_n360), .B2(new_n362), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n350), .A2(new_n399), .A3(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n280), .B1(new_n351), .B2(new_n264), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n294), .A2(new_n296), .ZN(new_n407));
  MUX2_X1   g0207(.A(G222), .B(G223), .S(G1698), .Z(new_n408));
  OR2_X1    g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n262), .B1(new_n407), .B2(new_n218), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n406), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(G190), .ZN(new_n412));
  INV_X1    g0212(.A(G50), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n413), .B1(new_n203), .B2(G20), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n252), .A2(new_n414), .B1(new_n413), .B2(new_n249), .ZN(new_n415));
  NOR2_X1   g0215(.A1(G58), .A2(G68), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n204), .B1(new_n416), .B2(new_n413), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT67), .ZN(new_n418));
  XNOR2_X1  g0218(.A(new_n417), .B(new_n418), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n255), .A2(new_n375), .B1(G150), .B2(new_n305), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n415), .B1(new_n421), .B2(new_n333), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT9), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n412), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n415), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n419), .A2(new_n420), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n425), .B1(new_n426), .B2(new_n251), .ZN(new_n427));
  OAI22_X1  g0227(.A1(new_n427), .A2(KEYINPUT9), .B1(new_n287), .B2(new_n411), .ZN(new_n428));
  OAI21_X1  g0228(.A(KEYINPUT10), .B1(new_n424), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n409), .A2(new_n410), .ZN(new_n430));
  INV_X1    g0230(.A(new_n406), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n422), .A2(new_n423), .B1(new_n432), .B2(G200), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n427), .A2(KEYINPUT9), .B1(G190), .B2(new_n411), .ZN(new_n434));
  XNOR2_X1  g0234(.A(KEYINPUT73), .B(KEYINPUT10), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n429), .A2(new_n436), .A3(KEYINPUT74), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n262), .B1(new_n407), .B2(new_n220), .ZN(new_n438));
  NOR2_X1   g0238(.A1(G232), .A2(G1698), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n439), .B1(new_n213), .B2(G1698), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n438), .B1(new_n407), .B2(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n351), .A2(new_n219), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n443));
  NOR3_X1   g0243(.A1(new_n443), .A2(new_n276), .A3(new_n278), .ZN(new_n444));
  OR3_X1    g0244(.A1(new_n442), .A2(new_n444), .A3(KEYINPUT69), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT69), .B1(new_n442), .B2(new_n444), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n441), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(G200), .ZN(new_n448));
  OAI211_X1 g0248(.A(G77), .B(new_n256), .C1(new_n394), .C2(new_n395), .ZN(new_n449));
  XNOR2_X1  g0249(.A(KEYINPUT15), .B(G87), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n451), .A2(new_n375), .B1(G20), .B2(G77), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n255), .B1(KEYINPUT70), .B2(new_n305), .ZN(new_n453));
  AND2_X1   g0253(.A1(new_n305), .A2(KEYINPUT70), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n389), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n455), .A2(new_n251), .B1(new_n218), .B2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n441), .A2(new_n445), .A3(G190), .A4(new_n446), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n448), .A2(new_n449), .A3(new_n457), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n447), .A2(new_n341), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n457), .A2(new_n449), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n441), .A2(new_n445), .A3(new_n337), .A4(new_n446), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT74), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n433), .A2(new_n465), .A3(new_n434), .A4(new_n435), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n411), .A2(new_n337), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n422), .B(new_n467), .C1(G169), .C2(new_n411), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n437), .A2(new_n464), .A3(new_n466), .A4(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT75), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OR2_X1    g0271(.A1(new_n469), .A2(new_n470), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n405), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n221), .A2(G1698), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n270), .B(new_n474), .C1(G257), .C2(G1698), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G303), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n477), .B1(new_n294), .B2(new_n296), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n443), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(G41), .ZN(new_n480));
  AND2_X1   g0280(.A1(KEYINPUT84), .A2(KEYINPUT5), .ZN(new_n481));
  NOR2_X1   g0281(.A1(KEYINPUT84), .A2(KEYINPUT5), .ZN(new_n482));
  OAI211_X1 g0282(.A(KEYINPUT85), .B(new_n480), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n203), .B(G45), .C1(new_n480), .C2(KEYINPUT5), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  AND3_X1   g0285(.A1(new_n483), .A2(new_n277), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT84), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT5), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(KEYINPUT84), .A2(KEYINPUT5), .ZN(new_n490));
  AOI21_X1  g0290(.A(G41), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OR2_X1    g0291(.A1(new_n491), .A2(KEYINPUT85), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n486), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n485), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n495), .A2(G270), .A3(new_n262), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n496), .A2(KEYINPUT88), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT88), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n443), .B1(new_n485), .B2(new_n494), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n498), .B1(new_n499), .B2(G270), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n479), .B(new_n493), .C1(new_n497), .C2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G33), .A2(G283), .ZN(new_n502));
  INV_X1    g0302(.A(G97), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n502), .B(new_n204), .C1(G33), .C2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(G116), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G20), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(new_n251), .A3(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT20), .ZN(new_n508));
  OR2_X1    g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n508), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n509), .A2(new_n510), .B1(new_n505), .B2(new_n456), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n505), .B1(new_n203), .B2(G33), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n512), .B1(new_n394), .B2(new_n395), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n501), .A2(new_n514), .A3(G169), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT21), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g0317(.A(new_n496), .B(KEYINPUT88), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n518), .A2(G190), .A3(new_n493), .A4(new_n479), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n501), .A2(G200), .ZN(new_n520));
  INV_X1    g0320(.A(new_n514), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n501), .A2(new_n364), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n514), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n501), .A2(new_n514), .A3(KEYINPUT21), .A4(G169), .ZN(new_n525));
  AND4_X1   g0325(.A1(new_n517), .A2(new_n522), .A3(new_n524), .A4(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(G1698), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n215), .A2(new_n527), .ZN(new_n528));
  OAI221_X1 g0328(.A(new_n528), .B1(G257), .B2(new_n527), .C1(new_n290), .C2(new_n291), .ZN(new_n529));
  NAND2_X1  g0329(.A1(G33), .A2(G294), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n262), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(G264), .B(new_n262), .C1(new_n491), .C2(new_n484), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT90), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n495), .A2(KEYINPUT90), .A3(G264), .A4(new_n262), .ZN(new_n535));
  AOI221_X4 g0335(.A(new_n531), .B1(new_n486), .B2(new_n492), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n364), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n531), .B1(new_n534), .B2(new_n535), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n493), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n341), .ZN(new_n540));
  NOR3_X1   g0340(.A1(new_n214), .A2(KEYINPUT22), .A3(G20), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n294), .A2(new_n296), .A3(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n204), .B(G87), .C1(new_n290), .C2(new_n291), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT89), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n543), .A2(new_n544), .A3(KEYINPUT22), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n544), .B1(new_n543), .B2(KEYINPUT22), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n542), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT23), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n204), .B2(G107), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n220), .A2(KEYINPUT23), .A3(G20), .ZN(new_n550));
  NAND2_X1  g0350(.A1(G33), .A2(G116), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n549), .A2(new_n550), .B1(new_n552), .B2(new_n204), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n547), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(KEYINPUT24), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT24), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n547), .A2(new_n556), .A3(new_n553), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n333), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n252), .B1(G1), .B2(new_n267), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n559), .A2(new_n220), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n249), .A2(new_n220), .ZN(new_n561));
  XNOR2_X1  g0361(.A(new_n561), .B(KEYINPUT25), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n537), .B(new_n540), .C1(new_n558), .C2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n538), .A2(new_n400), .A3(new_n493), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n536), .B2(G200), .ZN(new_n567));
  AND3_X1   g0367(.A1(new_n547), .A2(new_n556), .A3(new_n553), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n556), .B1(new_n547), .B2(new_n553), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n251), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n567), .A2(new_n570), .A3(new_n563), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n565), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n559), .A2(new_n503), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n249), .A2(new_n503), .ZN(new_n574));
  XNOR2_X1  g0374(.A(new_n574), .B(KEYINPUT82), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT6), .ZN(new_n577));
  AND2_X1   g0377(.A1(G97), .A2(G107), .ZN(new_n578));
  NOR2_X1   g0378(.A1(G97), .A2(G107), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n220), .A2(KEYINPUT81), .A3(KEYINPUT6), .A4(G97), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT81), .ZN(new_n582));
  NAND2_X1  g0382(.A1(KEYINPUT6), .A2(G97), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n582), .B1(new_n583), .B2(G107), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n580), .A2(new_n581), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(G20), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n305), .A2(G77), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n588), .B1(G107), .B2(new_n298), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n576), .B1(new_n589), .B2(new_n333), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT83), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n527), .A2(G244), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n592), .B1(new_n268), .B2(new_n269), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n591), .B1(new_n593), .B2(KEYINPUT4), .ZN(new_n594));
  OAI211_X1 g0394(.A(G244), .B(new_n527), .C1(new_n290), .C2(new_n291), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT4), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n595), .A2(KEYINPUT83), .A3(new_n596), .ZN(new_n597));
  OAI22_X1  g0397(.A1(new_n592), .A2(new_n596), .B1(new_n215), .B2(new_n527), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n598), .A2(new_n294), .A3(new_n296), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n594), .A2(new_n502), .A3(new_n597), .A4(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n443), .ZN(new_n601));
  OAI211_X1 g0401(.A(G257), .B(new_n262), .C1(new_n491), .C2(new_n484), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n483), .A2(new_n485), .A3(new_n277), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n491), .A2(KEYINPUT85), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n601), .A2(new_n337), .A3(new_n606), .ZN(new_n607));
  NOR3_X1   g0407(.A1(new_n593), .A2(new_n591), .A3(KEYINPUT4), .ZN(new_n608));
  AOI21_X1  g0408(.A(KEYINPUT83), .B1(new_n595), .B2(new_n596), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n599), .A2(new_n502), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n262), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n341), .B1(new_n612), .B2(new_n605), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n590), .A2(new_n607), .A3(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT82), .ZN(new_n615));
  XNOR2_X1  g0415(.A(new_n574), .B(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n616), .B1(new_n503), .B2(new_n559), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n585), .A2(G20), .B1(G77), .B2(new_n305), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n618), .B1(new_n329), .B2(new_n220), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n617), .B1(new_n619), .B2(new_n251), .ZN(new_n620));
  OAI21_X1  g0420(.A(G200), .B1(new_n612), .B2(new_n605), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n605), .B1(new_n443), .B2(new_n600), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(G190), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n620), .A2(new_n621), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n203), .A2(new_n276), .A3(G45), .ZN(new_n625));
  INV_X1    g0425(.A(G45), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n215), .B1(new_n626), .B2(G1), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n262), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n213), .A2(new_n527), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n219), .A2(G1698), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n629), .B(new_n630), .C1(new_n290), .C2(new_n291), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n631), .A2(new_n551), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n337), .B(new_n628), .C1(new_n632), .C2(new_n262), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n262), .B1(new_n631), .B2(new_n551), .ZN(new_n634));
  INV_X1    g0434(.A(new_n628), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n341), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n389), .A2(new_n451), .ZN(new_n639));
  AOI21_X1  g0439(.A(G20), .B1(new_n268), .B2(new_n269), .ZN(new_n640));
  XNOR2_X1  g0440(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n204), .A2(G33), .A3(G97), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n640), .A2(G68), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n579), .A2(new_n214), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT19), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(KEYINPUT86), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT86), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(KEYINPUT19), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n358), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n644), .B1(new_n649), .B2(G20), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n643), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n639), .B1(new_n651), .B2(new_n251), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n559), .A2(new_n450), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n638), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n644), .ZN(new_n656));
  INV_X1    g0456(.A(new_n358), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n647), .A2(KEYINPUT19), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n645), .A2(KEYINPUT86), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n657), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n656), .B1(new_n660), .B2(new_n204), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n641), .A2(new_n642), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n204), .B(G68), .C1(new_n290), .C2(new_n291), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n251), .B1(new_n661), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(G200), .B1(new_n634), .B2(new_n635), .ZN(new_n666));
  INV_X1    g0466(.A(new_n639), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n252), .B(G87), .C1(G1), .C2(new_n267), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n665), .A2(new_n666), .A3(new_n667), .A4(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT87), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n652), .A2(KEYINPUT87), .A3(new_n666), .A4(new_n668), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n634), .A2(new_n635), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(G190), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n671), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  AND4_X1   g0475(.A1(new_n614), .A2(new_n624), .A3(new_n655), .A4(new_n675), .ZN(new_n676));
  AND4_X1   g0476(.A1(new_n473), .A2(new_n526), .A3(new_n572), .A4(new_n676), .ZN(G372));
  INV_X1    g0477(.A(new_n468), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n344), .A2(new_n347), .ZN(new_n679));
  INV_X1    g0479(.A(new_n463), .ZN(new_n680));
  AOI22_X1  g0480(.A1(new_n374), .A2(new_n398), .B1(new_n404), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n316), .A2(new_n322), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT80), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n323), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n679), .B1(new_n681), .B2(new_n685), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n686), .A2(KEYINPUT94), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n437), .A2(new_n466), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n688), .B1(new_n686), .B2(KEYINPUT94), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n678), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n614), .A2(new_n624), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT91), .ZN(new_n692));
  AND4_X1   g0492(.A1(new_n665), .A2(new_n666), .A3(new_n667), .A4(new_n668), .ZN(new_n693));
  AOI22_X1  g0493(.A1(new_n693), .A2(new_n674), .B1(new_n638), .B2(new_n654), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n691), .A2(new_n692), .A3(new_n571), .A4(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n614), .A2(new_n624), .A3(new_n694), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n567), .A2(new_n570), .A3(new_n563), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT91), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n524), .A2(new_n525), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n699), .A2(new_n517), .A3(new_n565), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n695), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT93), .ZN(new_n702));
  AND3_X1   g0502(.A1(new_n601), .A2(new_n337), .A3(new_n606), .ZN(new_n703));
  AOI21_X1  g0503(.A(G169), .B1(new_n601), .B2(new_n606), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n705), .A2(new_n675), .A3(new_n590), .A4(new_n655), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT26), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n702), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n652), .A2(new_n653), .ZN(new_n709));
  INV_X1    g0509(.A(new_n674), .ZN(new_n710));
  OAI22_X1  g0510(.A1(new_n709), .A2(new_n637), .B1(new_n669), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n707), .B1(new_n614), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(KEYINPUT92), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n637), .B1(new_n652), .B2(new_n653), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n710), .B1(new_n693), .B2(KEYINPUT87), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n714), .B1(new_n715), .B2(new_n671), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n607), .B1(G169), .B2(new_n622), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(new_n620), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n716), .A2(KEYINPUT93), .A3(KEYINPUT26), .A4(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT92), .ZN(new_n720));
  OAI211_X1 g0520(.A(new_n720), .B(new_n707), .C1(new_n614), .C2(new_n711), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n708), .A2(new_n713), .A3(new_n719), .A4(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n701), .A2(new_n722), .A3(new_n655), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n473), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n690), .A2(new_n724), .ZN(G369));
  NAND2_X1  g0525(.A1(new_n699), .A2(new_n517), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n385), .A2(new_n204), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT95), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT27), .ZN(new_n729));
  OR2_X1    g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n728), .A2(new_n729), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n730), .A2(new_n731), .A3(G213), .ZN(new_n732));
  INV_X1    g0532(.A(G343), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n521), .ZN(new_n736));
  MUX2_X1   g0536(.A(new_n526), .B(new_n726), .S(new_n736), .Z(new_n737));
  AND2_X1   g0537(.A1(new_n737), .A2(G330), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n734), .B1(new_n558), .B2(new_n564), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n572), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(new_n565), .B2(new_n735), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n734), .B1(new_n699), .B2(new_n517), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n572), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n565), .A2(new_n734), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n742), .A2(new_n747), .ZN(G399));
  INV_X1    g0548(.A(new_n207), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G41), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n644), .A2(G116), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n751), .A2(G1), .A3(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(new_n228), .B2(new_n751), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n754), .B(KEYINPUT28), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n716), .A2(new_n707), .A3(new_n718), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n718), .A2(new_n694), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n714), .B1(new_n757), .B2(KEYINPUT26), .ZN(new_n758));
  AND3_X1   g0558(.A1(new_n699), .A2(new_n517), .A3(new_n565), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n691), .A2(new_n571), .A3(new_n694), .ZN(new_n760));
  OAI211_X1 g0560(.A(new_n756), .B(new_n758), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n761), .A2(KEYINPUT29), .A3(new_n735), .ZN(new_n762));
  AND2_X1   g0562(.A1(new_n723), .A2(new_n735), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n762), .B1(new_n763), .B2(KEYINPUT29), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n572), .A2(new_n526), .A3(new_n676), .A4(new_n735), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT30), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n518), .A2(G179), .A3(new_n493), .A4(new_n479), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n622), .A2(new_n538), .A3(new_n673), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n622), .A2(new_n338), .A3(new_n673), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(new_n501), .A3(new_n539), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  NOR3_X1   g0572(.A1(new_n767), .A2(new_n768), .A3(new_n766), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n734), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT31), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OAI211_X1 g0576(.A(KEYINPUT31), .B(new_n734), .C1(new_n772), .C2(new_n773), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n765), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G330), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n764), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(KEYINPUT96), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT96), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n764), .A2(new_n782), .A3(new_n779), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n755), .B1(new_n784), .B2(G1), .ZN(G364));
  NOR2_X1   g0585(.A1(new_n384), .A2(G20), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n203), .B1(new_n786), .B2(G45), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n750), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n738), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n790), .B1(G330), .B2(new_n737), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G13), .A2(G33), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(G20), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n226), .B1(G20), .B2(new_n341), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT97), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n749), .A2(new_n270), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(G45), .B2(new_n228), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n800), .B1(new_n246), .B2(G45), .ZN(new_n801));
  INV_X1    g0601(.A(new_n407), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n802), .A2(G355), .A3(new_n207), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(G116), .B2(new_n207), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n798), .B1(new_n801), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(new_n789), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n204), .A2(G190), .A3(G200), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n338), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(G311), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n337), .A2(new_n204), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n400), .A2(G200), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(G322), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n407), .B1(new_n808), .B2(new_n809), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  NOR3_X1   g0614(.A1(new_n400), .A2(G179), .A3(G200), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(new_n204), .ZN(new_n816));
  INV_X1    g0616(.A(G294), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n204), .A2(G179), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n818), .A2(G190), .A3(G200), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n816), .A2(new_n817), .B1(new_n819), .B2(new_n477), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n807), .A2(new_n364), .ZN(new_n821));
  INV_X1    g0621(.A(G329), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n818), .A2(new_n400), .A3(G200), .ZN(new_n823));
  INV_X1    g0623(.A(G283), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n821), .A2(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NOR3_X1   g0625(.A1(new_n814), .A2(new_n820), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n810), .A2(G200), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(G190), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(G326), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n828), .A2(new_n400), .ZN(new_n832));
  XOR2_X1   g0632(.A(KEYINPUT33), .B(G317), .Z(new_n833));
  OAI211_X1 g0633(.A(new_n826), .B(new_n831), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n832), .A2(new_n212), .B1(new_n503), .B2(new_n816), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT98), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(G58), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT32), .ZN(new_n839));
  INV_X1    g0639(.A(G159), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n821), .A2(new_n840), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n812), .A2(new_n838), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(new_n839), .B2(new_n841), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n830), .A2(G50), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n808), .A2(new_n218), .B1(new_n220), .B2(new_n823), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n819), .A2(new_n214), .ZN(new_n846));
  NOR3_X1   g0646(.A1(new_n845), .A2(new_n407), .A3(new_n846), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n837), .A2(new_n843), .A3(new_n844), .A4(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n835), .A2(new_n836), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n834), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n806), .B1(new_n850), .B2(new_n795), .ZN(new_n851));
  INV_X1    g0651(.A(new_n794), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n851), .B1(new_n737), .B2(new_n852), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n791), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(G396));
  INV_X1    g0655(.A(KEYINPUT100), .ZN(new_n856));
  INV_X1    g0656(.A(new_n459), .ZN(new_n857));
  NOR3_X1   g0657(.A1(new_n857), .A2(new_n680), .A3(new_n734), .ZN(new_n858));
  AND3_X1   g0658(.A1(new_n723), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n856), .B1(new_n723), .B2(new_n858), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n734), .A2(new_n461), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n463), .B1(new_n857), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n680), .A2(new_n735), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI22_X1  g0664(.A1(new_n859), .A2(new_n860), .B1(new_n763), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n789), .B1(new_n865), .B2(new_n779), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n779), .B2(new_n865), .ZN(new_n867));
  INV_X1    g0667(.A(new_n789), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n795), .A2(new_n792), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n868), .B1(new_n218), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n270), .B1(new_n823), .B2(new_n212), .ZN(new_n871));
  INV_X1    g0671(.A(new_n816), .ZN(new_n872));
  INV_X1    g0672(.A(new_n821), .ZN(new_n873));
  AOI22_X1  g0673(.A1(G58), .A2(new_n872), .B1(new_n873), .B2(G132), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n413), .B2(new_n819), .ZN(new_n875));
  INV_X1    g0675(.A(new_n812), .ZN(new_n876));
  INV_X1    g0676(.A(new_n808), .ZN(new_n877));
  AOI22_X1  g0677(.A1(new_n876), .A2(G143), .B1(new_n877), .B2(G159), .ZN(new_n878));
  INV_X1    g0678(.A(G137), .ZN(new_n879));
  INV_X1    g0679(.A(G150), .ZN(new_n880));
  OAI221_X1 g0680(.A(new_n878), .B1(new_n829), .B2(new_n879), .C1(new_n880), .C2(new_n832), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT34), .ZN(new_n882));
  AOI211_X1 g0682(.A(new_n871), .B(new_n875), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n882), .B2(new_n881), .ZN(new_n884));
  OAI221_X1 g0684(.A(new_n407), .B1(new_n503), .B2(new_n816), .C1(new_n812), .C2(new_n817), .ZN(new_n885));
  OAI22_X1  g0685(.A1(new_n821), .A2(new_n809), .B1(new_n819), .B2(new_n220), .ZN(new_n886));
  OAI22_X1  g0686(.A1(new_n808), .A2(new_n505), .B1(new_n214), .B2(new_n823), .ZN(new_n887));
  NOR3_X1   g0687(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  OAI221_X1 g0688(.A(new_n888), .B1(new_n824), .B2(new_n832), .C1(new_n477), .C2(new_n829), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n884), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n891), .A2(KEYINPUT99), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n795), .B1(new_n891), .B2(KEYINPUT99), .ZN(new_n893));
  OAI221_X1 g0693(.A(new_n870), .B1(new_n793), .B2(new_n864), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n867), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(G384));
  NOR2_X1   g0696(.A1(new_n786), .A2(new_n203), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT101), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n723), .A2(new_n858), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT100), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n723), .A2(new_n856), .A3(new_n858), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n900), .A2(new_n901), .B1(new_n680), .B2(new_n735), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n398), .A2(new_n734), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n399), .A2(new_n404), .A3(new_n903), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n398), .B(new_n734), .C1(new_n374), .C2(new_n403), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n898), .B1(new_n902), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n863), .B1(new_n859), .B2(new_n860), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(KEYINPUT101), .A3(new_n906), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n345), .B1(new_n336), .B2(new_n289), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT37), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n321), .A2(new_n259), .ZN(new_n913));
  INV_X1    g0713(.A(new_n732), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT102), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n913), .A2(KEYINPUT102), .A3(new_n914), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n911), .B(new_n912), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n334), .A2(KEYINPUT16), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n259), .B1(new_n918), .B2(new_n313), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n914), .ZN(new_n920));
  INV_X1    g0720(.A(new_n919), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n920), .B(new_n314), .C1(new_n921), .C2(new_n343), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(KEYINPUT37), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n917), .A2(new_n923), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n924), .B(KEYINPUT38), .C1(new_n350), .C2(new_n920), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n679), .A2(new_n684), .A3(new_n323), .ZN(new_n927));
  INV_X1    g0727(.A(new_n920), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT38), .B1(new_n929), .B2(new_n924), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n908), .A2(new_n910), .A3(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n916), .A2(new_n915), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n314), .B1(new_n336), .B2(new_n343), .ZN(new_n935));
  OAI21_X1  g0735(.A(KEYINPUT37), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n344), .A2(new_n347), .A3(new_n316), .A4(new_n322), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n936), .A2(new_n917), .B1(new_n937), .B2(new_n934), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n925), .B1(KEYINPUT38), .B2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT39), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n929), .A2(new_n924), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT38), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n944), .A2(KEYINPUT39), .A3(new_n925), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n399), .A2(new_n734), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n946), .A2(new_n947), .B1(new_n348), .B2(new_n732), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n933), .A2(new_n948), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n473), .B(new_n762), .C1(new_n763), .C2(KEYINPUT29), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n690), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n949), .B(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n906), .A2(new_n778), .A3(new_n864), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n936), .A2(new_n917), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n937), .A2(new_n934), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n943), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n953), .B1(new_n956), .B2(new_n925), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT40), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n906), .A2(new_n778), .A3(new_n958), .A4(new_n864), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n957), .A2(new_n958), .B1(new_n931), .B2(new_n959), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n473), .A2(new_n778), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n960), .A2(new_n961), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n962), .A2(G330), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n897), .B1(new_n952), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n952), .B2(new_n964), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n585), .A2(KEYINPUT35), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n585), .A2(KEYINPUT35), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n967), .A2(G116), .A3(new_n227), .A4(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT36), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n229), .A2(G77), .A3(new_n303), .A4(new_n301), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(G50), .B2(new_n212), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n972), .A2(G1), .A3(new_n384), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n966), .A2(new_n970), .A3(new_n973), .ZN(G367));
  NAND2_X1  g0774(.A1(new_n652), .A2(new_n668), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n734), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT103), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n977), .A2(new_n711), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(new_n714), .B2(new_n977), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n794), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n797), .B1(new_n749), .B2(new_n451), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n799), .A2(new_n239), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n868), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(G317), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n808), .A2(new_n824), .B1(new_n821), .B2(new_n984), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n292), .B1(new_n220), .B2(new_n816), .C1(new_n812), .C2(new_n477), .ZN(new_n986));
  INV_X1    g0786(.A(new_n823), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n985), .B(new_n986), .C1(G97), .C2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n819), .ZN(new_n989));
  AOI21_X1  g0789(.A(KEYINPUT107), .B1(new_n989), .B2(G116), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT46), .ZN(new_n991));
  INV_X1    g0791(.A(new_n832), .ZN(new_n992));
  AOI22_X1  g0792(.A1(G294), .A2(new_n992), .B1(new_n830), .B2(G311), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n988), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT108), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n802), .B1(new_n879), .B2(new_n821), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n816), .A2(new_n212), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(G77), .B2(new_n987), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n998), .B1(new_n413), .B2(new_n808), .C1(new_n838), .C2(new_n819), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n996), .B(new_n999), .C1(G150), .C2(new_n876), .ZN(new_n1000));
  INV_X1    g0800(.A(G143), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1000), .B1(new_n1001), .B2(new_n829), .C1(new_n840), .C2(new_n832), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n995), .A2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT47), .Z(new_n1004));
  INV_X1    g0804(.A(new_n795), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n980), .B(new_n983), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n734), .A2(new_n590), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n691), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1007), .A2(new_n717), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT104), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT105), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1015), .A2(KEYINPUT44), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n746), .A2(new_n1014), .A3(new_n1017), .ZN(new_n1018));
  AND2_X1   g0818(.A1(new_n1015), .A2(KEYINPUT44), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1014), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n747), .A2(KEYINPUT45), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT45), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n746), .B2(new_n1014), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n742), .B1(new_n1022), .B2(new_n1027), .ZN(new_n1028));
  AND4_X1   g0828(.A1(new_n742), .A2(new_n1027), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n744), .B1(new_n741), .B2(new_n743), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(new_n738), .Z(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(new_n781), .B2(new_n783), .ZN(new_n1033));
  AND3_X1   g0833(.A1(new_n1030), .A2(new_n1033), .A3(KEYINPUT106), .ZN(new_n1034));
  AOI21_X1  g0834(.A(KEYINPUT106), .B1(new_n1030), .B2(new_n1033), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n784), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n750), .B(KEYINPUT41), .Z(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n788), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1014), .A2(new_n744), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT42), .Z(new_n1041));
  OR2_X1    g0841(.A1(new_n1014), .A2(new_n565), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n734), .B1(new_n1042), .B2(new_n614), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT43), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n1041), .A2(new_n1043), .B1(new_n1044), .B2(new_n979), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n979), .A2(new_n1044), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1045), .B(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n742), .A2(new_n1014), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1047), .B(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1006), .B1(new_n1039), .B2(new_n1049), .ZN(G387));
  NOR2_X1   g0850(.A1(new_n1033), .A2(new_n751), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1032), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1051), .B1(new_n784), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n292), .B1(new_n823), .B2(new_n505), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n809), .A2(new_n832), .B1(new_n829), .B2(new_n813), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT112), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n876), .A2(G317), .B1(new_n877), .B2(G303), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT48), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n872), .A2(G283), .B1(new_n989), .B2(G294), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT49), .Z(new_n1066));
  AOI211_X1 g0866(.A(new_n1054), .B(new_n1066), .C1(G326), .C2(new_n873), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n832), .A2(new_n254), .B1(new_n212), .B2(new_n808), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT111), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n829), .A2(new_n840), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n816), .A2(new_n450), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1072), .B1(new_n218), .B2(new_n819), .C1(new_n880), .C2(new_n821), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n270), .B1(new_n503), .B2(new_n823), .C1(new_n812), .C2(new_n413), .ZN(new_n1074));
  NOR4_X1   g0874(.A1(new_n1069), .A2(new_n1070), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n795), .B1(new_n1067), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n799), .B1(new_n236), .B2(new_n626), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n752), .ZN(new_n1078));
  AOI211_X1 g0878(.A(G45), .B(new_n1078), .C1(G68), .C2(G77), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT109), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OR3_X1    g0881(.A1(new_n254), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1082));
  OAI21_X1  g0882(.A(KEYINPUT50), .B1(new_n254), .B2(G50), .ZN(new_n1083));
  AND3_X1   g0883(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1077), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n802), .A2(new_n207), .A3(new_n1078), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(G107), .B2(new_n207), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n1086), .A2(KEYINPUT110), .A3(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1089), .A2(new_n797), .ZN(new_n1090));
  OAI21_X1  g0890(.A(KEYINPUT110), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n868), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1076), .B(new_n1092), .C1(new_n741), .C2(new_n852), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1053), .B(new_n1093), .C1(new_n787), .C2(new_n1032), .ZN(G393));
  OAI221_X1 g0894(.A(new_n750), .B1(new_n1033), .B2(new_n1030), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1030), .A2(new_n788), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n798), .B1(new_n503), .B2(new_n207), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n799), .A2(new_n243), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n789), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n992), .A2(G50), .B1(new_n255), .B2(new_n877), .ZN(new_n1100));
  OR2_X1    g0900(.A1(new_n1100), .A2(KEYINPUT113), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(KEYINPUT113), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n270), .B1(new_n823), .B2(new_n214), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n816), .A2(new_n218), .B1(new_n819), .B2(new_n212), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n1103), .B(new_n1104), .C1(G143), .C2(new_n873), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1101), .A2(new_n1102), .A3(new_n1105), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n829), .A2(new_n880), .B1(new_n840), .B2(new_n812), .ZN(new_n1107));
  XOR2_X1   g0907(.A(new_n1107), .B(KEYINPUT51), .Z(new_n1108));
  OAI22_X1  g0908(.A1(new_n829), .A2(new_n984), .B1(new_n809), .B2(new_n812), .ZN(new_n1109));
  XOR2_X1   g0909(.A(new_n1109), .B(KEYINPUT52), .Z(new_n1110));
  OAI22_X1  g0910(.A1(new_n808), .A2(new_n817), .B1(new_n816), .B2(new_n505), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n407), .B1(new_n220), .B2(new_n823), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n821), .A2(new_n813), .B1(new_n819), .B2(new_n824), .ZN(new_n1113));
  NOR3_X1   g0913(.A1(new_n1111), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n477), .B2(new_n832), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n1106), .A2(new_n1108), .B1(new_n1110), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1099), .B1(new_n1116), .B2(new_n795), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n1023), .B2(new_n852), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1095), .A2(new_n1096), .A3(new_n1118), .ZN(G390));
  INV_X1    g0919(.A(new_n947), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT114), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n906), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(KEYINPUT114), .B1(new_n904), .B2(new_n905), .ZN(new_n1123));
  OR2_X1    g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n761), .A2(new_n735), .A3(new_n862), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n863), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1120), .B(new_n939), .C1(new_n1124), .C2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n947), .B1(new_n909), .B2(new_n906), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1128), .B1(new_n1129), .B2(new_n946), .ZN(new_n1130));
  AND3_X1   g0930(.A1(new_n778), .A2(G330), .A3(new_n864), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n906), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1130), .A2(new_n1133), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1132), .B(new_n1128), .C1(new_n1129), .C2(new_n946), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n778), .A2(G330), .A3(new_n864), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n907), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1132), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1126), .B1(new_n906), .B2(new_n1131), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1136), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n909), .A2(new_n1138), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n473), .A2(G330), .A3(new_n778), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n950), .A2(new_n690), .A3(new_n1142), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1134), .A2(new_n1135), .A3(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1144), .B(KEYINPUT115), .ZN(new_n1146));
  AND2_X1   g0946(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n750), .B(new_n1145), .C1(new_n1146), .C2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT117), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1134), .A2(new_n788), .A3(new_n1135), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n869), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n789), .B1(new_n255), .B2(new_n1151), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(G107), .A2(new_n992), .B1(new_n830), .B2(G283), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n872), .A2(G77), .B1(new_n987), .B2(G68), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n877), .A2(G97), .B1(new_n873), .B2(G294), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n802), .B(new_n846), .C1(new_n876), .C2(G116), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .A4(new_n1156), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n830), .A2(G128), .B1(G132), .B2(new_n876), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT116), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n992), .A2(G137), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT53), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n989), .A2(new_n1161), .A3(G150), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1161), .B1(new_n989), .B2(G150), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n407), .B(new_n1163), .C1(G159), .C2(new_n872), .ZN(new_n1164));
  INV_X1    g0964(.A(G125), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n821), .A2(new_n1165), .B1(new_n823), .B2(new_n413), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(KEYINPUT54), .B(G143), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1166), .B1(new_n877), .B2(new_n1168), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1160), .A2(new_n1162), .A3(new_n1164), .A4(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1157), .B1(new_n1159), .B2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1152), .B1(new_n1171), .B2(new_n795), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n946), .B2(new_n793), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1149), .B1(new_n1150), .B2(new_n1173), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n1150), .A2(new_n1149), .A3(new_n1173), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1148), .B1(new_n1174), .B2(new_n1175), .ZN(G378));
  INV_X1    g0976(.A(new_n1143), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1145), .A2(new_n1177), .ZN(new_n1178));
  AND3_X1   g0978(.A1(new_n906), .A2(new_n778), .A3(new_n864), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n958), .B1(new_n939), .B2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n959), .B1(new_n925), .B2(new_n944), .ZN(new_n1181));
  OAI21_X1  g0981(.A(G330), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n437), .A2(new_n466), .A3(new_n468), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n732), .A2(new_n427), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1183), .B(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1185), .B(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1182), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1187), .ZN(new_n1189));
  OAI211_X1 g0989(.A(G330), .B(new_n1189), .C1(new_n1180), .C2(new_n1181), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n949), .A2(new_n1191), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n933), .A2(new_n948), .A3(new_n1188), .A4(new_n1190), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1178), .A2(new_n1194), .A3(KEYINPUT57), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT119), .ZN(new_n1196));
  AND3_X1   g0996(.A1(new_n1188), .A2(new_n1196), .A3(new_n1190), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1196), .B1(new_n1188), .B2(new_n1190), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n949), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n1199), .A2(new_n1193), .B1(new_n1177), .B2(new_n1145), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n750), .B(new_n1195), .C1(new_n1200), .C2(KEYINPUT57), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(G97), .A2(new_n992), .B1(new_n830), .B2(G116), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n823), .A2(new_n838), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n821), .A2(new_n824), .B1(new_n819), .B2(new_n218), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1203), .B(new_n1204), .C1(new_n877), .C2(new_n451), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n292), .A2(new_n480), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n997), .B(new_n1206), .C1(new_n876), .C2(G107), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1202), .A2(new_n1205), .A3(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT58), .ZN(new_n1209));
  AOI21_X1  g1009(.A(G50), .B1(new_n267), .B2(new_n480), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1208), .A2(new_n1209), .B1(new_n1206), .B2(new_n1210), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(G125), .A2(new_n830), .B1(new_n992), .B2(G132), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n819), .A2(new_n1167), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n1214), .A2(KEYINPUT118), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n877), .A2(G137), .B1(G150), .B2(new_n872), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n876), .A2(G128), .B1(KEYINPUT118), .B2(new_n1214), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1212), .A2(new_n1215), .A3(new_n1216), .A4(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(KEYINPUT59), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n267), .B(new_n480), .C1(new_n823), .C2(new_n840), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(G124), .B2(new_n873), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1219), .A2(new_n1221), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1218), .A2(KEYINPUT59), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1211), .B1(new_n1209), .B2(new_n1208), .C1(new_n1222), .C2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n795), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n868), .B1(new_n413), .B2(new_n869), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1225), .B(new_n1226), .C1(new_n1189), .C2(new_n793), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1199), .A2(new_n1193), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1228), .B1(new_n1229), .B2(new_n788), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1201), .A2(new_n1230), .ZN(G375));
  NAND2_X1  g1031(.A1(new_n1124), .A2(new_n792), .ZN(new_n1232));
  XOR2_X1   g1032(.A(new_n1232), .B(KEYINPUT121), .Z(new_n1233));
  OAI21_X1  g1033(.A(new_n1072), .B1(new_n812), .B2(new_n824), .ZN(new_n1234));
  XOR2_X1   g1034(.A(new_n1234), .B(KEYINPUT122), .Z(new_n1235));
  OAI21_X1  g1035(.A(new_n407), .B1(new_n218), .B2(new_n823), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n877), .A2(G107), .B1(G97), .B2(new_n989), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n477), .B2(new_n821), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n505), .A2(new_n832), .B1(new_n829), .B2(new_n817), .ZN(new_n1239));
  NOR4_X1   g1039(.A1(new_n1235), .A2(new_n1236), .A3(new_n1238), .A4(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n830), .A2(G132), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT123), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1241), .B(new_n1242), .ZN(new_n1243));
  OAI221_X1 g1043(.A(new_n1243), .B1(new_n879), .B2(new_n812), .C1(new_n832), .C2(new_n1167), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1244), .A2(KEYINPUT124), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n808), .A2(new_n880), .B1(new_n816), .B2(new_n413), .ZN(new_n1247));
  INV_X1    g1047(.A(G128), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n821), .A2(new_n1248), .B1(new_n819), .B2(new_n840), .ZN(new_n1249));
  NOR4_X1   g1049(.A1(new_n1247), .A2(new_n1249), .A3(new_n292), .A4(new_n1203), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n1244), .B2(KEYINPUT124), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1240), .B1(new_n1246), .B2(new_n1252), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n789), .B1(G68), .B2(new_n1151), .C1(new_n1253), .C2(new_n1005), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1138), .A2(new_n909), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  XOR2_X1   g1058(.A(new_n787), .B(KEYINPUT120), .Z(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n1233), .A2(new_n1255), .B1(new_n1258), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n1038), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1261), .B1(new_n1146), .B2(new_n1263), .ZN(G381));
  NOR4_X1   g1064(.A1(G393), .A2(G381), .A3(G396), .A4(G384), .ZN(new_n1265));
  INV_X1    g1065(.A(G390), .ZN(new_n1266));
  AND2_X1   g1066(.A1(new_n1150), .A2(new_n1173), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1148), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1265), .A2(new_n1266), .A3(new_n1269), .ZN(new_n1270));
  OR3_X1    g1070(.A1(new_n1270), .A2(G387), .A3(G375), .ZN(G407));
  NAND2_X1  g1071(.A1(new_n733), .A2(G213), .ZN(new_n1272));
  OR3_X1    g1072(.A1(G375), .A2(new_n1268), .A3(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(G407), .A2(G213), .A3(new_n1273), .ZN(G409));
  AND3_X1   g1074(.A1(new_n1201), .A2(G378), .A3(new_n1230), .ZN(new_n1275));
  AND4_X1   g1075(.A1(new_n933), .A2(new_n948), .A3(new_n1188), .A4(new_n1190), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(new_n933), .A2(new_n948), .B1(new_n1188), .B2(new_n1190), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1260), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n1227), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n941), .A2(new_n945), .ZN(new_n1280));
  OAI22_X1  g1080(.A1(new_n1280), .A2(new_n1120), .B1(new_n679), .B2(new_n914), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n909), .A2(new_n906), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n931), .B1(new_n1282), .B2(new_n898), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1281), .B1(new_n1283), .B2(new_n910), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1189), .B1(new_n960), .B2(G330), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1190), .ZN(new_n1286));
  OAI21_X1  g1086(.A(KEYINPUT119), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1188), .A2(new_n1196), .A3(new_n1190), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1284), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1178), .B(new_n1038), .C1(new_n1276), .C2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT125), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1279), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1229), .A2(KEYINPUT125), .A3(new_n1038), .A4(new_n1178), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1268), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1272), .B1(new_n1275), .B2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT126), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT60), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1297), .B1(new_n1258), .B2(new_n1177), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1258), .A2(new_n1177), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n750), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(KEYINPUT60), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1301), .A2(new_n1262), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1296), .B1(new_n1300), .B2(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n751), .B1(new_n1301), .B2(new_n1262), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1304), .A2(KEYINPUT126), .A3(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1303), .A2(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(G384), .B1(new_n1307), .B2(new_n1261), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1261), .ZN(new_n1309));
  AOI211_X1 g1109(.A(new_n895), .B(new_n1309), .C1(new_n1303), .C2(new_n1306), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n733), .A2(G213), .A3(G2897), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1311), .ZN(new_n1312));
  NOR3_X1   g1112(.A1(new_n1308), .A2(new_n1310), .A3(new_n1312), .ZN(new_n1313));
  NOR3_X1   g1113(.A1(new_n1300), .A2(new_n1302), .A3(new_n1296), .ZN(new_n1314));
  AOI21_X1  g1114(.A(KEYINPUT126), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1261), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n895), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1307), .A2(G384), .A3(new_n1261), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1311), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1313), .A2(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(KEYINPUT61), .B1(new_n1295), .B2(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1201), .A2(G378), .A3(new_n1230), .ZN(new_n1322));
  AND2_X1   g1122(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1322), .B1(new_n1323), .B2(new_n1268), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT62), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1308), .A2(new_n1310), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1324), .A2(new_n1325), .A3(new_n1272), .A4(new_n1326), .ZN(new_n1327));
  OAI211_X1 g1127(.A(new_n1272), .B(new_n1326), .C1(new_n1275), .C2(new_n1294), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1328), .A2(KEYINPUT62), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1321), .A2(new_n1327), .A3(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT127), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(G387), .A2(new_n1266), .ZN(new_n1332));
  OAI211_X1 g1132(.A(G390), .B(new_n1006), .C1(new_n1039), .C2(new_n1049), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1331), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1334));
  XNOR2_X1  g1134(.A(G393), .B(new_n854), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1335), .ZN(new_n1336));
  XNOR2_X1  g1136(.A(new_n1334), .B(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1330), .A2(new_n1337), .ZN(new_n1338));
  XNOR2_X1  g1138(.A(new_n1334), .B(new_n1335), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT63), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1328), .A2(new_n1340), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1324), .A2(KEYINPUT63), .A3(new_n1272), .A4(new_n1326), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1339), .A2(new_n1341), .A3(new_n1321), .A4(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1338), .A2(new_n1343), .ZN(G405));
  NAND2_X1  g1144(.A1(G375), .A2(new_n1269), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1345), .A2(new_n1322), .ZN(new_n1346));
  AND2_X1   g1146(.A1(new_n1346), .A2(new_n1326), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1346), .A2(new_n1326), .ZN(new_n1348));
  NOR2_X1   g1148(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1349), .A2(new_n1339), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n1337), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1350), .A2(new_n1351), .ZN(G402));
endmodule


