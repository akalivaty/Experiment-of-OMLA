//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 0 1 1 0 1 0 0 0 0 0 0 1 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 0 0 1 0 0 1 1 0 0 0 1 0 1 1 0 1 0 1 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966;
  INV_X1    g000(.A(KEYINPUT25), .ZN(new_n187));
  XNOR2_X1  g001(.A(G125), .B(G140), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT16), .ZN(new_n189));
  INV_X1    g003(.A(G125), .ZN(new_n190));
  OR3_X1    g004(.A1(new_n190), .A2(KEYINPUT16), .A3(G140), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n189), .A2(G146), .A3(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n188), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G128), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(KEYINPUT23), .A3(G119), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(G119), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n196), .B(new_n198), .C1(new_n200), .C2(KEYINPUT23), .ZN(new_n201));
  OR2_X1    g015(.A1(new_n201), .A2(G110), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT24), .B(G110), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n196), .A2(new_n199), .ZN(new_n204));
  AND2_X1   g018(.A1(new_n204), .A2(KEYINPUT75), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n204), .A2(KEYINPUT75), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n203), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n202), .A2(new_n207), .A3(KEYINPUT76), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(KEYINPUT76), .B1(new_n202), .B2(new_n207), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n192), .B(new_n194), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n201), .A2(G110), .ZN(new_n212));
  OR2_X1    g026(.A1(new_n205), .A2(new_n206), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n212), .B1(new_n213), .B2(new_n203), .ZN(new_n214));
  INV_X1    g028(.A(new_n192), .ZN(new_n215));
  AOI21_X1  g029(.A(G146), .B1(new_n189), .B2(new_n191), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n211), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT22), .B(G137), .ZN(new_n221));
  INV_X1    g035(.A(G953), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n222), .A2(G221), .A3(G234), .ZN(new_n223));
  XNOR2_X1  g037(.A(new_n221), .B(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n211), .A2(new_n219), .A3(new_n224), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n187), .B1(new_n228), .B2(G902), .ZN(new_n229));
  INV_X1    g043(.A(G902), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n226), .A2(new_n227), .A3(KEYINPUT25), .A4(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G217), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n233), .B1(G234), .B2(new_n230), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n234), .A2(G902), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n235), .B1(new_n228), .B2(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(G472), .A2(G902), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT66), .ZN(new_n240));
  INV_X1    g054(.A(G131), .ZN(new_n241));
  INV_X1    g055(.A(G137), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G134), .ZN(new_n243));
  INV_X1    g057(.A(G134), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G137), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n241), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n246), .A2(KEYINPUT65), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT65), .ZN(new_n248));
  AOI211_X1 g062(.A(new_n248), .B(new_n241), .C1(new_n243), .C2(new_n245), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G143), .ZN(new_n251));
  OAI21_X1  g065(.A(KEYINPUT1), .B1(new_n251), .B2(G146), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(G146), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n193), .A2(G143), .ZN(new_n254));
  OAI211_X1 g068(.A(G128), .B(new_n252), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n193), .A2(G143), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n251), .A2(G146), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n256), .B(new_n257), .C1(KEYINPUT1), .C2(new_n197), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT11), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n259), .B1(new_n244), .B2(G137), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n242), .A2(KEYINPUT11), .A3(G134), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n260), .A2(new_n261), .A3(new_n241), .A4(new_n245), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n255), .A2(new_n258), .A3(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n240), .B1(new_n250), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n260), .A2(new_n261), .A3(new_n245), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(KEYINPUT64), .A3(G131), .ZN(new_n266));
  NAND2_X1  g080(.A1(KEYINPUT64), .A2(G131), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n260), .A2(new_n261), .A3(new_n267), .A4(new_n245), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n256), .A2(new_n257), .A3(KEYINPUT0), .A4(G128), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n253), .A2(new_n254), .ZN(new_n271));
  XNOR2_X1  g085(.A(KEYINPUT0), .B(G128), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n255), .A2(new_n258), .A3(new_n262), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n246), .A2(KEYINPUT65), .ZN(new_n277));
  XNOR2_X1  g091(.A(G134), .B(G137), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n248), .B1(new_n278), .B2(new_n241), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n276), .A2(KEYINPUT66), .A3(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n264), .A2(new_n275), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT30), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AND2_X1   g098(.A1(KEYINPUT2), .A2(G113), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT2), .ZN(new_n286));
  INV_X1    g100(.A(G113), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n287), .A3(KEYINPUT67), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT67), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n289), .B1(KEYINPUT2), .B2(G113), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n285), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  XNOR2_X1  g105(.A(G116), .B(G119), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n195), .A2(G116), .ZN(new_n294));
  INV_X1    g108(.A(G116), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G119), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT69), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT69), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n292), .A2(new_n299), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n298), .B(new_n300), .C1(new_n291), .C2(KEYINPUT68), .ZN(new_n301));
  AND2_X1   g115(.A1(new_n291), .A2(KEYINPUT68), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n293), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  AOI22_X1  g117(.A1(new_n274), .A2(new_n269), .B1(new_n276), .B2(new_n280), .ZN(new_n304));
  AOI21_X1  g118(.A(KEYINPUT70), .B1(new_n304), .B2(KEYINPUT30), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n276), .A2(new_n280), .ZN(new_n306));
  AND4_X1   g120(.A1(KEYINPUT70), .A2(new_n306), .A3(new_n275), .A4(KEYINPUT30), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n284), .B(new_n303), .C1(new_n305), .C2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n275), .ZN(new_n309));
  OR2_X1    g123(.A1(new_n309), .A2(new_n303), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n311));
  INV_X1    g125(.A(G210), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n312), .A2(G237), .A3(G953), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n311), .B(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT26), .B(G101), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n314), .B(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n308), .A2(new_n310), .A3(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT72), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n308), .A2(KEYINPUT72), .A3(new_n310), .A4(new_n316), .ZN(new_n320));
  AND3_X1   g134(.A1(new_n319), .A2(KEYINPUT31), .A3(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT28), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n310), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n282), .A2(new_n303), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT73), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n282), .A2(KEYINPUT73), .A3(new_n303), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(new_n310), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n324), .B1(new_n329), .B2(KEYINPUT28), .ZN(new_n330));
  OAI22_X1  g144(.A1(new_n330), .A2(new_n316), .B1(KEYINPUT31), .B2(new_n317), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n239), .B1(new_n321), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT74), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT32), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n328), .A2(new_n310), .ZN(new_n335));
  AOI21_X1  g149(.A(KEYINPUT73), .B1(new_n282), .B2(new_n303), .ZN(new_n336));
  OAI21_X1  g150(.A(KEYINPUT28), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n316), .B1(new_n337), .B2(new_n323), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n317), .A2(KEYINPUT31), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n319), .A2(KEYINPUT31), .A3(new_n320), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT74), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n342), .A2(new_n343), .A3(new_n239), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n333), .A2(new_n334), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G472), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n330), .A2(new_n316), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT29), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n308), .A2(new_n310), .ZN(new_n349));
  INV_X1    g163(.A(new_n316), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n347), .A2(new_n348), .A3(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n309), .B(new_n303), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT28), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n354), .A2(KEYINPUT29), .A3(new_n316), .A4(new_n323), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n355), .A2(new_n230), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n346), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n239), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n358), .B1(new_n340), .B2(new_n341), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n357), .B1(KEYINPUT32), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n238), .B1(new_n345), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(G214), .B1(G237), .B2(G902), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n363), .B(KEYINPUT84), .ZN(new_n364));
  XNOR2_X1  g178(.A(KEYINPUT81), .B(G101), .ZN(new_n365));
  INV_X1    g179(.A(G104), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G107), .ZN(new_n367));
  INV_X1    g181(.A(G107), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G104), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT79), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n367), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT80), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(new_n368), .A3(G104), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT3), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n374), .A2(new_n370), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n375), .B1(new_n374), .B2(new_n370), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n365), .B(new_n372), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  NOR3_X1   g192(.A1(new_n366), .A2(KEYINPUT80), .A3(G107), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT3), .B1(new_n379), .B2(KEYINPUT79), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n374), .A2(new_n370), .A3(new_n375), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n371), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G101), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n378), .B(KEYINPUT4), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n372), .B1(new_n376), .B2(new_n377), .ZN(new_n385));
  XOR2_X1   g199(.A(KEYINPUT82), .B(KEYINPUT4), .Z(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(G101), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n384), .A2(new_n303), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT85), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT5), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n391), .B1(new_n298), .B2(new_n300), .ZN(new_n392));
  OAI21_X1  g206(.A(G113), .B1(new_n294), .B2(KEYINPUT5), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n293), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n383), .B1(new_n369), .B2(new_n367), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n378), .A2(new_n396), .ZN(new_n397));
  OR2_X1    g211(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n384), .A2(KEYINPUT85), .A3(new_n303), .A4(new_n387), .ZN(new_n399));
  XNOR2_X1  g213(.A(G110), .B(G122), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n390), .A2(new_n398), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT87), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n399), .A2(new_n398), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT87), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n403), .A2(new_n404), .A3(new_n390), .A4(new_n400), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n255), .A2(new_n258), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n190), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT88), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n408), .B(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n273), .A2(G125), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G224), .ZN(new_n413));
  OAI21_X1  g227(.A(KEYINPUT7), .B1(new_n413), .B2(G953), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n395), .B1(new_n382), .B2(new_n365), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n394), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n400), .B(KEYINPUT8), .ZN(new_n417));
  AOI21_X1  g231(.A(KEYINPUT89), .B1(new_n292), .B2(KEYINPUT5), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n418), .A2(new_n393), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n292), .A2(KEYINPUT89), .A3(KEYINPUT5), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n419), .A2(new_n420), .B1(new_n291), .B2(new_n292), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n417), .B1(new_n421), .B2(new_n397), .ZN(new_n422));
  OAI22_X1  g236(.A1(new_n412), .A2(new_n414), .B1(new_n416), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT90), .ZN(new_n424));
  OR2_X1    g238(.A1(new_n410), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n410), .A2(new_n424), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n426), .A3(new_n411), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n423), .B1(new_n427), .B2(new_n414), .ZN(new_n428));
  AOI21_X1  g242(.A(G902), .B1(new_n406), .B2(new_n428), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n303), .A2(new_n387), .ZN(new_n430));
  AOI21_X1  g244(.A(KEYINPUT85), .B1(new_n430), .B2(new_n384), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n399), .A2(new_n398), .ZN(new_n432));
  OAI21_X1  g246(.A(KEYINPUT86), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT86), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n390), .A2(new_n434), .A3(new_n398), .A4(new_n399), .ZN(new_n435));
  INV_X1    g249(.A(new_n400), .ZN(new_n436));
  AND4_X1   g250(.A1(KEYINPUT6), .A2(new_n433), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n406), .A2(KEYINPUT6), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n390), .A2(new_n398), .A3(new_n399), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n400), .B1(new_n439), .B2(KEYINPUT86), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n435), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n437), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n413), .A2(G953), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n412), .B(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n429), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(G210), .B1(G237), .B2(G902), .ZN(new_n447));
  XOR2_X1   g261(.A(new_n447), .B(KEYINPUT91), .Z(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n429), .B(new_n447), .C1(new_n442), .C2(new_n445), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n364), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G237), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(new_n222), .A3(G214), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(G143), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT18), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n454), .B1(new_n455), .B2(new_n241), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n453), .B(new_n251), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(KEYINPUT18), .A3(G131), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n188), .B(new_n193), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n456), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(G113), .B(G122), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(G104), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT92), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n464), .B1(new_n457), .B2(G131), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n454), .A2(KEYINPUT92), .A3(new_n241), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n457), .A2(G131), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  XOR2_X1   g282(.A(KEYINPUT93), .B(KEYINPUT19), .Z(new_n469));
  NOR2_X1   g283(.A1(new_n469), .A2(new_n188), .ZN(new_n470));
  NAND2_X1  g284(.A1(KEYINPUT93), .A2(KEYINPUT19), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n470), .B1(new_n188), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n215), .B1(new_n472), .B2(new_n193), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n463), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT94), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT17), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n475), .B1(new_n467), .B2(new_n476), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n457), .A2(KEYINPUT94), .A3(KEYINPUT17), .A4(G131), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n465), .A2(new_n466), .A3(new_n476), .A4(new_n467), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n479), .A2(new_n217), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n460), .ZN(new_n482));
  INV_X1    g296(.A(new_n462), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n474), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(G475), .A2(G902), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(KEYINPUT20), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT20), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n484), .A2(new_n489), .A3(new_n486), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n483), .A2(KEYINPUT95), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n230), .B1(new_n482), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n492), .B1(new_n481), .B2(new_n460), .ZN(new_n495));
  OAI21_X1  g309(.A(G475), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT96), .ZN(new_n499));
  INV_X1    g313(.A(G122), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n499), .B1(new_n500), .B2(G116), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n295), .A2(KEYINPUT96), .A3(G122), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n500), .A2(G116), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(G107), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n503), .A2(new_n368), .A3(new_n504), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n251), .A2(G128), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n197), .A2(G143), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n511), .A3(new_n244), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT13), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n511), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n510), .A2(new_n513), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT97), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT97), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n510), .A2(new_n517), .A3(new_n513), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n514), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n512), .B1(new_n519), .B2(new_n244), .ZN(new_n520));
  OR2_X1    g334(.A1(new_n503), .A2(KEYINPUT14), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n503), .A2(KEYINPUT14), .B1(G116), .B2(new_n500), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n368), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n510), .A2(new_n511), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(G134), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n512), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n507), .ZN(new_n527));
  OAI22_X1  g341(.A1(new_n509), .A2(new_n520), .B1(new_n523), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT9), .B(G234), .ZN(new_n529));
  NOR3_X1   g343(.A1(new_n529), .A2(new_n233), .A3(G953), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  OR2_X1    g346(.A1(new_n523), .A2(new_n527), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n508), .B(new_n512), .C1(new_n244), .C2(new_n519), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n530), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n230), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT98), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n528), .A2(new_n531), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n533), .A2(new_n534), .A3(new_n530), .ZN(new_n539));
  AOI21_X1  g353(.A(G902), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT98), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT15), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(G478), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT99), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n545), .B1(new_n540), .B2(new_n541), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n537), .A2(new_n542), .B1(new_n544), .B2(G478), .ZN(new_n551));
  OAI21_X1  g365(.A(KEYINPUT99), .B1(new_n551), .B2(new_n548), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(G952), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n554), .A2(G953), .ZN(new_n555));
  NAND2_X1  g369(.A1(G234), .A2(G237), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT21), .B(G898), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n556), .A2(G902), .A3(G953), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n557), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n498), .A2(new_n553), .A3(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(G469), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n384), .A2(new_n274), .A3(new_n387), .ZN(new_n565));
  INV_X1    g379(.A(new_n269), .ZN(new_n566));
  INV_X1    g380(.A(new_n407), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(new_n378), .A3(new_n396), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT10), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n415), .A2(KEYINPUT10), .A3(new_n567), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n565), .A2(new_n566), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(G110), .B(G140), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n222), .A2(G227), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n573), .B(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT12), .ZN(new_n578));
  OAI21_X1  g392(.A(KEYINPUT83), .B1(new_n415), .B2(new_n567), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT83), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n397), .A2(new_n580), .A3(new_n407), .ZN(new_n581));
  AOI22_X1  g395(.A1(new_n579), .A2(new_n581), .B1(new_n567), .B2(new_n415), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n578), .B1(new_n582), .B2(new_n566), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n415), .A2(KEYINPUT83), .A3(new_n567), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n580), .B1(new_n397), .B2(new_n407), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n568), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n586), .A2(KEYINPUT12), .A3(new_n269), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n577), .B1(new_n583), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n565), .A2(new_n570), .A3(new_n571), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n269), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n576), .B1(new_n590), .B2(new_n572), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n564), .B(new_n230), .C1(new_n588), .C2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n590), .A2(new_n576), .A3(new_n572), .ZN(new_n593));
  INV_X1    g407(.A(new_n572), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n594), .B1(new_n583), .B2(new_n587), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n575), .B(KEYINPUT78), .ZN(new_n596));
  OAI211_X1 g410(.A(G469), .B(new_n593), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(G469), .A2(G902), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n592), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(G221), .B1(new_n529), .B2(G902), .ZN(new_n600));
  XOR2_X1   g414(.A(new_n600), .B(KEYINPUT77), .Z(new_n601));
  NAND2_X1  g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n451), .A2(new_n563), .A3(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n362), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(new_n365), .ZN(G3));
  INV_X1    g420(.A(new_n447), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n446), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n364), .B1(new_n608), .B2(new_n450), .ZN(new_n609));
  OR2_X1    g423(.A1(new_n532), .A2(KEYINPUT101), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n532), .A2(KEYINPUT101), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n610), .A2(KEYINPUT33), .A3(new_n538), .A4(new_n611), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT100), .B(KEYINPUT33), .Z(new_n613));
  OAI21_X1  g427(.A(new_n613), .B1(new_n532), .B2(new_n535), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n230), .A2(G478), .ZN(new_n616));
  OAI22_X1  g430(.A1(new_n615), .A2(new_n616), .B1(G478), .B2(new_n540), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n497), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  AND3_X1   g433(.A1(new_n609), .A2(new_n561), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n342), .A2(new_n230), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(G472), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n622), .A2(new_n333), .A3(new_n344), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n238), .A2(new_n602), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n620), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT34), .B(G104), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G6));
  NOR2_X1   g442(.A1(new_n553), .A2(new_n497), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n609), .A2(new_n561), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n630), .A2(new_n624), .A3(new_n625), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT35), .B(G107), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G9));
  NAND2_X1  g447(.A1(new_n220), .A2(KEYINPUT102), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n225), .A2(KEYINPUT36), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT102), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n211), .A2(new_n219), .A3(new_n636), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n634), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n635), .B1(new_n634), .B2(new_n637), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n236), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n235), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n562), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n624), .A2(new_n451), .A3(new_n603), .A4(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT37), .B(G110), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G12));
  AOI21_X1  g459(.A(new_n641), .B1(new_n345), .B2(new_n360), .ZN(new_n646));
  AOI211_X1 g460(.A(new_n364), .B(new_n602), .C1(new_n608), .C2(new_n450), .ZN(new_n647));
  XOR2_X1   g461(.A(new_n557), .B(KEYINPUT103), .Z(new_n648));
  OAI21_X1  g462(.A(new_n648), .B1(G900), .B2(new_n560), .ZN(new_n649));
  XOR2_X1   g463(.A(new_n649), .B(KEYINPUT104), .Z(new_n650));
  NOR3_X1   g464(.A1(new_n553), .A2(new_n497), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n646), .A2(new_n647), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT105), .B(G128), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G30));
  INV_X1    g468(.A(KEYINPUT108), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n449), .A2(new_n450), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n656), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n235), .A2(new_n640), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n660), .A2(new_n364), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n319), .A2(new_n320), .ZN(new_n663));
  AND2_X1   g477(.A1(new_n353), .A2(new_n350), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n230), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  AOI22_X1  g479(.A1(new_n359), .A2(KEYINPUT32), .B1(G472), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n345), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n497), .A2(new_n552), .A3(new_n550), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n662), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n650), .B(KEYINPUT39), .Z(new_n672));
  NAND2_X1  g486(.A1(new_n603), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT107), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT40), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n655), .B1(new_n671), .B2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n675), .B(KEYINPUT40), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n679), .A2(new_n662), .A3(KEYINPUT108), .A4(new_n670), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(new_n251), .ZN(G45));
  NOR2_X1   g496(.A1(new_n618), .A2(new_n650), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n646), .A2(new_n647), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G146), .ZN(G48));
  INV_X1    g499(.A(new_n561), .ZN(new_n686));
  AOI211_X1 g500(.A(new_n686), .B(new_n364), .C1(new_n608), .C2(new_n450), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n230), .B1(new_n588), .B2(new_n591), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(G469), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n689), .A2(new_n592), .A3(new_n600), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT109), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n689), .A2(KEYINPUT109), .A3(new_n592), .A4(new_n600), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n361), .A2(new_n687), .A3(new_n619), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT41), .B(G113), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G15));
  NAND4_X1  g512(.A1(new_n361), .A2(new_n687), .A3(new_n629), .A4(new_n695), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G116), .ZN(G18));
  AOI211_X1 g514(.A(new_n364), .B(new_n690), .C1(new_n608), .C2(new_n450), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n646), .A2(new_n701), .A3(new_n563), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G119), .ZN(G21));
  AOI21_X1  g517(.A(new_n316), .B1(new_n354), .B2(new_n323), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n339), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n358), .B1(new_n705), .B2(new_n341), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n621), .A2(KEYINPUT110), .A3(G472), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT110), .ZN(new_n708));
  AOI21_X1  g522(.A(G902), .B1(new_n340), .B2(new_n341), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n708), .B1(new_n709), .B2(new_n346), .ZN(new_n710));
  AOI211_X1 g524(.A(new_n238), .B(new_n706), .C1(new_n707), .C2(new_n710), .ZN(new_n711));
  AOI211_X1 g525(.A(new_n364), .B(new_n669), .C1(new_n608), .C2(new_n450), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n692), .A2(new_n561), .A3(new_n693), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n711), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G122), .ZN(G24));
  AOI211_X1 g530(.A(new_n706), .B(new_n641), .C1(new_n707), .C2(new_n710), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n683), .A3(new_n701), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G125), .ZN(G27));
  NAND2_X1  g533(.A1(new_n599), .A2(new_n600), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT111), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n599), .A2(KEYINPUT111), .A3(new_n600), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n364), .ZN(new_n725));
  INV_X1    g539(.A(new_n429), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n440), .A2(KEYINPUT6), .A3(new_n435), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n440), .A2(new_n435), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT6), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n729), .B1(new_n402), .B2(new_n405), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n727), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n726), .B1(new_n731), .B2(new_n444), .ZN(new_n732));
  INV_X1    g546(.A(new_n448), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n450), .B(new_n725), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n724), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n332), .A2(new_n334), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n238), .B1(new_n360), .B2(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n735), .A2(new_n737), .A3(KEYINPUT42), .A4(new_n683), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n361), .A2(new_n735), .A3(new_n683), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT112), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT42), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n739), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n740), .B1(new_n739), .B2(new_n741), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n738), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G131), .ZN(G33));
  NAND3_X1  g559(.A1(new_n361), .A2(new_n735), .A3(new_n651), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G134), .ZN(G36));
  NAND2_X1  g561(.A1(new_n498), .A2(new_n617), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(KEYINPUT43), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n749), .A2(new_n624), .A3(new_n641), .ZN(new_n750));
  OR2_X1    g564(.A1(new_n750), .A2(KEYINPUT44), .ZN(new_n751));
  INV_X1    g565(.A(new_n734), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n593), .B1(new_n595), .B2(new_n596), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n754));
  OR2_X1    g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n564), .B1(new_n753), .B2(new_n754), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n598), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT46), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n592), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n758), .A2(new_n759), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n600), .B(new_n672), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n750), .A2(KEYINPUT44), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n751), .A2(new_n752), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  XOR2_X1   g580(.A(KEYINPUT113), .B(G137), .Z(new_n767));
  XNOR2_X1  g581(.A(new_n766), .B(new_n767), .ZN(G39));
  OAI21_X1  g582(.A(new_n600), .B1(new_n761), .B2(new_n762), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(KEYINPUT47), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n345), .A2(new_n360), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n772), .A2(new_n238), .A3(new_n683), .A4(new_n752), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G140), .ZN(G42));
  NAND2_X1  g589(.A1(new_n554), .A2(new_n222), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n646), .B(new_n647), .C1(new_n651), .C2(new_n683), .ZN(new_n777));
  INV_X1    g591(.A(new_n669), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n660), .A2(new_n720), .A3(new_n650), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n667), .A2(new_n609), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n777), .A2(new_n718), .A3(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT52), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n696), .A2(new_n699), .A3(new_n715), .A4(new_n702), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(KEYINPUT114), .ZN(new_n784));
  AOI211_X1 g598(.A(new_n641), .B(new_n562), .C1(new_n345), .C2(new_n360), .ZN(new_n785));
  INV_X1    g599(.A(new_n450), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n731), .A2(new_n444), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n447), .B1(new_n787), .B2(new_n429), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n725), .B(new_n778), .C1(new_n786), .C2(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(new_n713), .ZN(new_n790));
  AOI22_X1  g604(.A1(new_n785), .A2(new_n701), .B1(new_n790), .B2(new_n711), .ZN(new_n791));
  AOI211_X1 g605(.A(new_n238), .B(new_n694), .C1(new_n345), .C2(new_n360), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n792), .B1(new_n620), .B2(new_n630), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT114), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n791), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n546), .A2(new_n549), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n498), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n686), .B1(new_n797), .B2(new_n618), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n624), .A2(new_n451), .A3(new_n625), .A4(new_n798), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n643), .B(new_n799), .C1(new_n362), .C2(new_n604), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n717), .A2(new_n683), .A3(new_n735), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n497), .A2(new_n796), .A3(new_n650), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n603), .A2(new_n802), .A3(new_n660), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n771), .A2(new_n752), .A3(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n801), .A2(new_n746), .A3(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n800), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n744), .A2(new_n784), .A3(new_n795), .A4(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n782), .B1(new_n807), .B2(KEYINPUT115), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n784), .A2(new_n795), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT115), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n809), .A2(new_n810), .A3(new_n744), .A4(new_n806), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT116), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n808), .A2(KEYINPUT53), .A3(new_n811), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n808), .A2(new_n811), .A3(KEYINPUT116), .A4(KEYINPUT53), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n817), .A2(KEYINPUT54), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT53), .B1(new_n808), .B2(new_n811), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n813), .B1(new_n783), .B2(KEYINPUT117), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n791), .A2(new_n793), .A3(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n821), .A2(new_n744), .A3(new_n806), .A4(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(KEYINPUT118), .B1(new_n824), .B2(new_n782), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n744), .A2(new_n806), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n696), .A2(new_n699), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n715), .A2(new_n702), .ZN(new_n828));
  OAI21_X1  g642(.A(KEYINPUT117), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n829), .A2(KEYINPUT53), .A3(new_n823), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT52), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n781), .B(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n826), .A2(new_n830), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n825), .A2(new_n834), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n820), .A2(new_n835), .A3(KEYINPUT54), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n819), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n749), .A2(new_n648), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n711), .ZN(new_n840));
  NOR4_X1   g654(.A1(new_n840), .A2(new_n725), .A3(new_n659), .A4(new_n690), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(KEYINPUT50), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n689), .A2(new_n592), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n770), .B1(new_n601), .B2(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n844), .A2(new_n711), .A3(new_n752), .A4(new_n839), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n734), .A2(new_n690), .ZN(new_n846));
  NOR4_X1   g660(.A1(new_n846), .A2(new_n667), .A3(new_n238), .A4(new_n557), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n497), .A2(new_n617), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n846), .A2(new_n749), .A3(new_n648), .ZN(new_n849));
  AOI22_X1  g663(.A1(new_n847), .A2(new_n848), .B1(new_n849), .B2(new_n717), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n842), .A2(new_n845), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT51), .ZN(new_n852));
  OR2_X1    g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n851), .A2(new_n852), .ZN(new_n854));
  INV_X1    g668(.A(new_n701), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n555), .B1(new_n840), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n849), .A2(new_n737), .ZN(new_n857));
  XOR2_X1   g671(.A(new_n857), .B(KEYINPUT48), .Z(new_n858));
  AOI211_X1 g672(.A(new_n856), .B(new_n858), .C1(new_n619), .C2(new_n847), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n853), .A2(new_n854), .A3(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n776), .B1(new_n838), .B2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n238), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n862), .A2(new_n725), .A3(new_n601), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n843), .A2(KEYINPUT49), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n863), .A2(new_n748), .A3(new_n864), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n865), .B(new_n668), .C1(KEYINPUT49), .C2(new_n843), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n866), .A2(new_n659), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n861), .A2(new_n867), .ZN(G75));
  OAI21_X1  g682(.A(G902), .B1(new_n820), .B2(new_n835), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(KEYINPUT119), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n871), .B(G902), .C1(new_n820), .C2(new_n835), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n870), .A2(new_n448), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n442), .A2(new_n445), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n787), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT55), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n876), .A2(KEYINPUT56), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n222), .A2(G952), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT56), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n880), .B1(new_n869), .B2(new_n312), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n879), .B1(new_n881), .B2(new_n876), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n878), .A2(new_n882), .ZN(G51));
  XOR2_X1   g697(.A(new_n598), .B(KEYINPUT57), .Z(new_n884));
  INV_X1    g698(.A(KEYINPUT54), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n825), .A2(new_n834), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n885), .B1(new_n814), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n884), .B1(new_n887), .B2(new_n836), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n888), .B1(new_n591), .B2(new_n588), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n870), .A2(new_n755), .A3(new_n756), .A4(new_n872), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n879), .B1(new_n889), .B2(new_n890), .ZN(G54));
  AND2_X1   g705(.A1(KEYINPUT58), .A2(G475), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n870), .A2(new_n872), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n485), .ZN(new_n894));
  INV_X1    g708(.A(new_n879), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n870), .A2(new_n484), .A3(new_n872), .A4(new_n892), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(G60));
  INV_X1    g711(.A(new_n615), .ZN(new_n898));
  NAND2_X1  g712(.A1(G478), .A2(G902), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT59), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n898), .B(new_n900), .C1(new_n887), .C2(new_n836), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n895), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n838), .A2(new_n900), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n902), .B1(new_n903), .B2(new_n615), .ZN(G63));
  NAND2_X1  g718(.A1(G217), .A2(G902), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT120), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT60), .ZN(new_n907));
  OAI221_X1 g721(.A(new_n907), .B1(new_n638), .B2(new_n639), .C1(new_n820), .C2(new_n835), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n895), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n228), .B(KEYINPUT121), .Z(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n814), .A2(new_n886), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n911), .B1(new_n912), .B2(new_n907), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT61), .ZN(new_n914));
  OR3_X1    g728(.A1(new_n909), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n914), .B1(new_n909), .B2(new_n913), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(G66));
  INV_X1    g731(.A(new_n809), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n918), .A2(new_n800), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n919), .A2(G953), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT122), .ZN(new_n921));
  OAI21_X1  g735(.A(G953), .B1(new_n558), .B2(new_n413), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n442), .B1(G898), .B2(new_n222), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n923), .B(new_n924), .ZN(G69));
  OAI21_X1  g739(.A(new_n284), .B1(new_n305), .B2(new_n307), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(new_n472), .Z(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT123), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n777), .A2(new_n718), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n678), .A2(new_n680), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(KEYINPUT62), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n774), .A2(new_n766), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT62), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n678), .A2(new_n680), .A3(new_n933), .A4(new_n929), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n734), .B1(new_n618), .B2(new_n797), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n675), .A2(new_n361), .A3(new_n935), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n931), .A2(new_n932), .A3(new_n934), .A4(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n928), .B1(new_n937), .B2(new_n222), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n764), .A2(new_n712), .A3(new_n737), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n939), .A2(new_n746), .A3(new_n929), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n932), .A2(new_n744), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n222), .ZN(new_n942));
  INV_X1    g756(.A(new_n927), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(G900), .B2(G953), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n938), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n222), .B1(G227), .B2(G900), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n945), .B(new_n946), .Z(G72));
  XNOR2_X1  g761(.A(KEYINPUT124), .B(KEYINPUT63), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n346), .A2(new_n230), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n948), .B(new_n949), .Z(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n951), .B1(new_n941), .B2(new_n919), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n349), .B(KEYINPUT126), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n350), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT127), .Z(new_n955));
  OAI21_X1  g769(.A(new_n895), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n919), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n950), .B1(new_n937), .B2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT125), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI211_X1 g774(.A(KEYINPUT125), .B(new_n950), .C1(new_n937), .C2(new_n957), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n953), .A2(new_n350), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n956), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n319), .A2(new_n320), .A3(new_n351), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n817), .A2(new_n818), .A3(new_n950), .A4(new_n965), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n964), .A2(new_n966), .ZN(G57));
endmodule


