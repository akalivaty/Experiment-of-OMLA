

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591;

  XNOR2_X1 U322 ( .A(n459), .B(KEYINPUT38), .ZN(n511) );
  XOR2_X1 U323 ( .A(n480), .B(KEYINPUT28), .Z(n537) );
  NAND2_X1 U324 ( .A1(n543), .A2(n484), .ZN(n290) );
  AND2_X1 U325 ( .A1(G226GAT), .A2(G233GAT), .ZN(n291) );
  XOR2_X1 U326 ( .A(G64GAT), .B(G92GAT), .Z(n292) );
  NAND2_X1 U327 ( .A1(n588), .A2(n587), .ZN(n293) );
  INV_X1 U328 ( .A(KEYINPUT25), .ZN(n391) );
  XNOR2_X1 U329 ( .A(n391), .B(KEYINPUT102), .ZN(n392) );
  XNOR2_X1 U330 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n441) );
  XNOR2_X1 U331 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U332 ( .A(n442), .B(n441), .ZN(n446) );
  XNOR2_X1 U333 ( .A(n379), .B(n291), .ZN(n380) );
  NOR2_X1 U334 ( .A1(n477), .A2(n476), .ZN(n478) );
  XNOR2_X1 U335 ( .A(n442), .B(n380), .ZN(n381) );
  NOR2_X1 U336 ( .A1(n589), .A2(n421), .ZN(n422) );
  XNOR2_X1 U337 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U338 ( .A(n386), .B(n385), .ZN(n388) );
  INV_X1 U339 ( .A(G43GAT), .ZN(n460) );
  XNOR2_X1 U340 ( .A(KEYINPUT96), .B(n414), .ZN(n584) );
  XNOR2_X1 U341 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U342 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U343 ( .A(n488), .B(n487), .ZN(G1349GAT) );
  XNOR2_X1 U344 ( .A(n463), .B(n462), .ZN(G1330GAT) );
  XOR2_X1 U345 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n294) );
  XNOR2_X1 U346 ( .A(KEYINPUT37), .B(n294), .ZN(n423) );
  XNOR2_X1 U347 ( .A(KEYINPUT36), .B(KEYINPUT106), .ZN(n313) );
  XOR2_X1 U348 ( .A(KEYINPUT11), .B(KEYINPUT70), .Z(n296) );
  XNOR2_X1 U349 ( .A(G92GAT), .B(KEYINPUT71), .ZN(n295) );
  XNOR2_X1 U350 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U351 ( .A(n297), .B(G106GAT), .Z(n299) );
  XOR2_X1 U352 ( .A(G50GAT), .B(KEYINPUT69), .Z(n332) );
  XNOR2_X1 U353 ( .A(G218GAT), .B(n332), .ZN(n298) );
  XNOR2_X1 U354 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U355 ( .A(G99GAT), .B(G85GAT), .Z(n451) );
  XOR2_X1 U356 ( .A(n300), .B(n451), .Z(n303) );
  XNOR2_X1 U357 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n301) );
  XNOR2_X1 U358 ( .A(n301), .B(KEYINPUT7), .ZN(n430) );
  XOR2_X1 U359 ( .A(G29GAT), .B(G134GAT), .Z(n402) );
  XNOR2_X1 U360 ( .A(n430), .B(n402), .ZN(n302) );
  XNOR2_X1 U361 ( .A(n303), .B(n302), .ZN(n312) );
  XOR2_X1 U362 ( .A(KEYINPUT65), .B(KEYINPUT10), .Z(n305) );
  XNOR2_X1 U363 ( .A(KEYINPUT9), .B(KEYINPUT72), .ZN(n304) );
  XNOR2_X1 U364 ( .A(n305), .B(n304), .ZN(n310) );
  XNOR2_X1 U365 ( .A(G36GAT), .B(G190GAT), .ZN(n306) );
  XNOR2_X1 U366 ( .A(n306), .B(KEYINPUT73), .ZN(n382) );
  XOR2_X1 U367 ( .A(n382), .B(G162GAT), .Z(n308) );
  NAND2_X1 U368 ( .A1(G232GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U369 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U370 ( .A(n310), .B(n309), .Z(n311) );
  XOR2_X1 U371 ( .A(n312), .B(n311), .Z(n469) );
  XOR2_X1 U372 ( .A(n313), .B(n469), .Z(n589) );
  XOR2_X1 U373 ( .A(G64GAT), .B(G57GAT), .Z(n315) );
  XNOR2_X1 U374 ( .A(G211GAT), .B(G155GAT), .ZN(n314) );
  XNOR2_X1 U375 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U376 ( .A(G71GAT), .B(KEYINPUT13), .Z(n443) );
  XOR2_X1 U377 ( .A(n316), .B(n443), .Z(n318) );
  XNOR2_X1 U378 ( .A(G127GAT), .B(G78GAT), .ZN(n317) );
  XNOR2_X1 U379 ( .A(n318), .B(n317), .ZN(n323) );
  XOR2_X1 U380 ( .A(G8GAT), .B(G183GAT), .Z(n379) );
  XNOR2_X1 U381 ( .A(G15GAT), .B(G22GAT), .ZN(n319) );
  XNOR2_X1 U382 ( .A(n319), .B(G1GAT), .ZN(n434) );
  XOR2_X1 U383 ( .A(n379), .B(n434), .Z(n321) );
  NAND2_X1 U384 ( .A1(G231GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U385 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U386 ( .A(n323), .B(n322), .Z(n331) );
  XOR2_X1 U387 ( .A(KEYINPUT12), .B(KEYINPUT74), .Z(n325) );
  XNOR2_X1 U388 ( .A(KEYINPUT14), .B(KEYINPUT78), .ZN(n324) );
  XNOR2_X1 U389 ( .A(n325), .B(n324), .ZN(n329) );
  XOR2_X1 U390 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n327) );
  XNOR2_X1 U391 ( .A(KEYINPUT75), .B(KEYINPUT15), .ZN(n326) );
  XNOR2_X1 U392 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U393 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U394 ( .A(n331), .B(n330), .Z(n582) );
  INV_X1 U395 ( .A(n582), .ZN(n561) );
  XOR2_X1 U396 ( .A(KEYINPUT101), .B(KEYINPUT26), .Z(n377) );
  XOR2_X1 U397 ( .A(KEYINPUT22), .B(KEYINPUT85), .Z(n334) );
  XOR2_X1 U398 ( .A(G106GAT), .B(G78GAT), .Z(n448) );
  XNOR2_X1 U399 ( .A(n332), .B(n448), .ZN(n333) );
  XNOR2_X1 U400 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U401 ( .A(n335), .B(KEYINPUT24), .Z(n342) );
  XOR2_X1 U402 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n337) );
  XNOR2_X1 U403 ( .A(G218GAT), .B(KEYINPUT21), .ZN(n336) );
  XNOR2_X1 U404 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U405 ( .A(n338), .B(KEYINPUT89), .Z(n340) );
  XNOR2_X1 U406 ( .A(G197GAT), .B(G211GAT), .ZN(n339) );
  XNOR2_X1 U407 ( .A(n340), .B(n339), .ZN(n384) );
  XNOR2_X1 U408 ( .A(G22GAT), .B(n384), .ZN(n341) );
  XNOR2_X1 U409 ( .A(n342), .B(n341), .ZN(n346) );
  XOR2_X1 U410 ( .A(KEYINPUT23), .B(KEYINPUT86), .Z(n344) );
  NAND2_X1 U411 ( .A1(G228GAT), .A2(G233GAT), .ZN(n343) );
  XNOR2_X1 U412 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U413 ( .A(n346), .B(n345), .Z(n354) );
  XOR2_X1 U414 ( .A(G148GAT), .B(G155GAT), .Z(n348) );
  XNOR2_X1 U415 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n347) );
  XNOR2_X1 U416 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U417 ( .A(KEYINPUT2), .B(KEYINPUT90), .Z(n350) );
  XNOR2_X1 U418 ( .A(G162GAT), .B(KEYINPUT91), .ZN(n349) );
  XNOR2_X1 U419 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U420 ( .A(n352), .B(n351), .Z(n410) );
  XNOR2_X1 U421 ( .A(n410), .B(G204GAT), .ZN(n353) );
  XNOR2_X1 U422 ( .A(n354), .B(n353), .ZN(n480) );
  XOR2_X1 U423 ( .A(G127GAT), .B(KEYINPUT0), .Z(n356) );
  XNOR2_X1 U424 ( .A(G113GAT), .B(KEYINPUT79), .ZN(n355) );
  XNOR2_X1 U425 ( .A(n356), .B(n355), .ZN(n401) );
  XOR2_X1 U426 ( .A(n401), .B(G99GAT), .Z(n358) );
  NAND2_X1 U427 ( .A1(G227GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U428 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U429 ( .A(n359), .B(G190GAT), .Z(n367) );
  XOR2_X1 U430 ( .A(KEYINPUT82), .B(KEYINPUT17), .Z(n361) );
  XNOR2_X1 U431 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n360) );
  XNOR2_X1 U432 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U433 ( .A(G169GAT), .B(n362), .ZN(n387) );
  XOR2_X1 U434 ( .A(G71GAT), .B(G176GAT), .Z(n364) );
  XNOR2_X1 U435 ( .A(G15GAT), .B(G183GAT), .ZN(n363) );
  XNOR2_X1 U436 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U437 ( .A(n387), .B(n365), .Z(n366) );
  XNOR2_X1 U438 ( .A(n367), .B(n366), .ZN(n375) );
  XOR2_X1 U439 ( .A(KEYINPUT83), .B(KEYINPUT84), .Z(n369) );
  XNOR2_X1 U440 ( .A(KEYINPUT20), .B(KEYINPUT81), .ZN(n368) );
  XNOR2_X1 U441 ( .A(n369), .B(n368), .ZN(n373) );
  XOR2_X1 U442 ( .A(KEYINPUT80), .B(G120GAT), .Z(n371) );
  XNOR2_X1 U443 ( .A(G43GAT), .B(G134GAT), .ZN(n370) );
  XNOR2_X1 U444 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U445 ( .A(n373), .B(n372), .Z(n374) );
  XNOR2_X1 U446 ( .A(n375), .B(n374), .ZN(n567) );
  NAND2_X1 U447 ( .A1(n480), .A2(n567), .ZN(n376) );
  XNOR2_X1 U448 ( .A(n377), .B(n376), .ZN(n586) );
  XNOR2_X1 U449 ( .A(KEYINPUT27), .B(KEYINPUT99), .ZN(n389) );
  XNOR2_X1 U450 ( .A(G176GAT), .B(G204GAT), .ZN(n378) );
  XNOR2_X1 U451 ( .A(n292), .B(n378), .ZN(n442) );
  XOR2_X1 U452 ( .A(n381), .B(KEYINPUT97), .Z(n386) );
  XNOR2_X1 U453 ( .A(n382), .B(KEYINPUT98), .ZN(n383) );
  XNOR2_X1 U454 ( .A(n388), .B(n387), .ZN(n529) );
  XOR2_X1 U455 ( .A(n389), .B(n529), .Z(n415) );
  NOR2_X1 U456 ( .A1(n586), .A2(n415), .ZN(n553) );
  NOR2_X1 U457 ( .A1(n567), .A2(n529), .ZN(n390) );
  NOR2_X1 U458 ( .A1(n480), .A2(n390), .ZN(n393) );
  NOR2_X1 U459 ( .A1(n553), .A2(n394), .ZN(n395) );
  XNOR2_X1 U460 ( .A(KEYINPUT103), .B(n395), .ZN(n413) );
  XOR2_X1 U461 ( .A(KEYINPUT5), .B(KEYINPUT94), .Z(n397) );
  XNOR2_X1 U462 ( .A(KEYINPUT95), .B(KEYINPUT93), .ZN(n396) );
  XNOR2_X1 U463 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U464 ( .A(n398), .B(G85GAT), .Z(n400) );
  XOR2_X1 U465 ( .A(G120GAT), .B(G57GAT), .Z(n447) );
  XNOR2_X1 U466 ( .A(G1GAT), .B(n447), .ZN(n399) );
  XNOR2_X1 U467 ( .A(n400), .B(n399), .ZN(n406) );
  XOR2_X1 U468 ( .A(n402), .B(n401), .Z(n404) );
  NAND2_X1 U469 ( .A1(G225GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U470 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U471 ( .A(n406), .B(n405), .Z(n412) );
  XOR2_X1 U472 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n408) );
  XNOR2_X1 U473 ( .A(KEYINPUT92), .B(KEYINPUT6), .ZN(n407) );
  XNOR2_X1 U474 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U475 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U476 ( .A(n412), .B(n411), .ZN(n414) );
  NAND2_X1 U477 ( .A1(n413), .A2(n414), .ZN(n420) );
  INV_X1 U478 ( .A(n415), .ZN(n416) );
  NAND2_X1 U479 ( .A1(n537), .A2(n416), .ZN(n417) );
  NOR2_X1 U480 ( .A1(n584), .A2(n417), .ZN(n541) );
  XNOR2_X1 U481 ( .A(KEYINPUT100), .B(n541), .ZN(n418) );
  NAND2_X1 U482 ( .A1(n418), .A2(n567), .ZN(n419) );
  NAND2_X1 U483 ( .A1(n420), .A2(n419), .ZN(n496) );
  NAND2_X1 U484 ( .A1(n561), .A2(n496), .ZN(n421) );
  XOR2_X1 U485 ( .A(n423), .B(n422), .Z(n526) );
  XOR2_X1 U486 ( .A(G8GAT), .B(G141GAT), .Z(n425) );
  XNOR2_X1 U487 ( .A(G169GAT), .B(G197GAT), .ZN(n424) );
  XNOR2_X1 U488 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U489 ( .A(KEYINPUT67), .B(KEYINPUT30), .Z(n427) );
  XNOR2_X1 U490 ( .A(KEYINPUT66), .B(KEYINPUT29), .ZN(n426) );
  XNOR2_X1 U491 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U492 ( .A(n429), .B(n428), .ZN(n440) );
  XOR2_X1 U493 ( .A(n430), .B(KEYINPUT68), .Z(n432) );
  NAND2_X1 U494 ( .A1(G229GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U495 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U496 ( .A(n433), .B(G50GAT), .ZN(n438) );
  XOR2_X1 U497 ( .A(G29GAT), .B(G36GAT), .Z(n436) );
  XNOR2_X1 U498 ( .A(G113GAT), .B(n434), .ZN(n435) );
  XNOR2_X1 U499 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U500 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U501 ( .A(n440), .B(n439), .Z(n554) );
  XNOR2_X1 U502 ( .A(G148GAT), .B(n443), .ZN(n444) );
  XNOR2_X1 U503 ( .A(n444), .B(KEYINPUT33), .ZN(n445) );
  XNOR2_X1 U504 ( .A(n446), .B(n445), .ZN(n450) );
  XNOR2_X1 U505 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U506 ( .A(n450), .B(n449), .ZN(n452) );
  NAND2_X1 U507 ( .A1(n452), .A2(n451), .ZN(n456) );
  INV_X1 U508 ( .A(n451), .ZN(n454) );
  INV_X1 U509 ( .A(n452), .ZN(n453) );
  NAND2_X1 U510 ( .A1(n454), .A2(n453), .ZN(n455) );
  NAND2_X1 U511 ( .A1(n456), .A2(n455), .ZN(n458) );
  NAND2_X1 U512 ( .A1(G230GAT), .A2(G233GAT), .ZN(n457) );
  XOR2_X2 U513 ( .A(n458), .B(n457), .Z(n577) );
  NOR2_X1 U514 ( .A1(n554), .A2(n577), .ZN(n497) );
  NAND2_X1 U515 ( .A1(n526), .A2(n497), .ZN(n459) );
  NOR2_X1 U516 ( .A1(n511), .A2(n567), .ZN(n463) );
  XNOR2_X1 U517 ( .A(KEYINPUT40), .B(KEYINPUT110), .ZN(n461) );
  INV_X1 U518 ( .A(n554), .ZN(n574) );
  NOR2_X1 U519 ( .A1(n561), .A2(n589), .ZN(n464) );
  XNOR2_X1 U520 ( .A(KEYINPUT45), .B(n464), .ZN(n466) );
  INV_X1 U521 ( .A(n577), .ZN(n465) );
  NAND2_X1 U522 ( .A1(n466), .A2(n465), .ZN(n467) );
  XOR2_X1 U523 ( .A(KEYINPUT121), .B(n467), .Z(n468) );
  NOR2_X1 U524 ( .A1(n574), .A2(n468), .ZN(n477) );
  INV_X1 U525 ( .A(n469), .ZN(n564) );
  NAND2_X1 U526 ( .A1(n561), .A2(n564), .ZN(n474) );
  XOR2_X1 U527 ( .A(KEYINPUT120), .B(KEYINPUT46), .Z(n472) );
  XNOR2_X1 U528 ( .A(n577), .B(KEYINPUT64), .ZN(n470) );
  XOR2_X1 U529 ( .A(n470), .B(KEYINPUT41), .Z(n543) );
  AND2_X1 U530 ( .A1(n543), .A2(n574), .ZN(n471) );
  XOR2_X1 U531 ( .A(n472), .B(n471), .Z(n473) );
  NOR2_X1 U532 ( .A1(n474), .A2(n473), .ZN(n475) );
  XOR2_X1 U533 ( .A(KEYINPUT47), .B(n475), .Z(n476) );
  XNOR2_X1 U534 ( .A(KEYINPUT48), .B(n478), .ZN(n551) );
  NOR2_X1 U535 ( .A1(n529), .A2(n551), .ZN(n479) );
  XNOR2_X1 U536 ( .A(n479), .B(KEYINPUT54), .ZN(n587) );
  INV_X1 U537 ( .A(n480), .ZN(n481) );
  AND2_X1 U538 ( .A1(n584), .A2(n481), .ZN(n482) );
  AND2_X1 U539 ( .A1(n587), .A2(n482), .ZN(n483) );
  XNOR2_X1 U540 ( .A(n483), .B(KEYINPUT55), .ZN(n566) );
  INV_X1 U541 ( .A(n567), .ZN(n484) );
  OR2_X1 U542 ( .A1(n566), .A2(n290), .ZN(n488) );
  XOR2_X1 U543 ( .A(G176GAT), .B(KEYINPUT57), .Z(n486) );
  XOR2_X1 U544 ( .A(KEYINPUT123), .B(KEYINPUT56), .Z(n485) );
  INV_X1 U545 ( .A(G190GAT), .ZN(n493) );
  XNOR2_X1 U546 ( .A(KEYINPUT124), .B(KEYINPUT58), .ZN(n491) );
  OR2_X1 U547 ( .A1(n567), .A2(n564), .ZN(n489) );
  NOR2_X1 U548 ( .A1(n566), .A2(n489), .ZN(n490) );
  XNOR2_X1 U549 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U550 ( .A(n493), .B(n492), .ZN(G1351GAT) );
  NAND2_X1 U551 ( .A1(n564), .A2(n582), .ZN(n494) );
  XOR2_X1 U552 ( .A(KEYINPUT16), .B(n494), .Z(n495) );
  AND2_X1 U553 ( .A1(n496), .A2(n495), .ZN(n514) );
  NAND2_X1 U554 ( .A1(n497), .A2(n514), .ZN(n498) );
  XNOR2_X1 U555 ( .A(KEYINPUT104), .B(n498), .ZN(n504) );
  NOR2_X1 U556 ( .A1(n504), .A2(n584), .ZN(n499) );
  XOR2_X1 U557 ( .A(G1GAT), .B(n499), .Z(n500) );
  XNOR2_X1 U558 ( .A(KEYINPUT34), .B(n500), .ZN(G1324GAT) );
  NOR2_X1 U559 ( .A1(n504), .A2(n529), .ZN(n501) );
  XOR2_X1 U560 ( .A(G8GAT), .B(n501), .Z(G1325GAT) );
  NOR2_X1 U561 ( .A1(n504), .A2(n567), .ZN(n503) );
  XNOR2_X1 U562 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n503), .B(n502), .ZN(G1326GAT) );
  XNOR2_X1 U564 ( .A(G22GAT), .B(KEYINPUT105), .ZN(n506) );
  NOR2_X1 U565 ( .A1(n537), .A2(n504), .ZN(n505) );
  XNOR2_X1 U566 ( .A(n506), .B(n505), .ZN(G1327GAT) );
  NOR2_X1 U567 ( .A1(n511), .A2(n584), .ZN(n509) );
  XOR2_X1 U568 ( .A(G29GAT), .B(KEYINPUT109), .Z(n507) );
  XNOR2_X1 U569 ( .A(KEYINPUT39), .B(n507), .ZN(n508) );
  XNOR2_X1 U570 ( .A(n509), .B(n508), .ZN(G1328GAT) );
  NOR2_X1 U571 ( .A1(n511), .A2(n529), .ZN(n510) );
  XOR2_X1 U572 ( .A(G36GAT), .B(n510), .Z(G1329GAT) );
  NOR2_X1 U573 ( .A1(n537), .A2(n511), .ZN(n512) );
  XOR2_X1 U574 ( .A(G50GAT), .B(n512), .Z(G1331GAT) );
  NAND2_X1 U575 ( .A1(n554), .A2(n543), .ZN(n513) );
  XNOR2_X1 U576 ( .A(n513), .B(KEYINPUT111), .ZN(n527) );
  NAND2_X1 U577 ( .A1(n527), .A2(n514), .ZN(n515) );
  XNOR2_X1 U578 ( .A(n515), .B(KEYINPUT112), .ZN(n523) );
  NOR2_X1 U579 ( .A1(n523), .A2(n584), .ZN(n517) );
  XNOR2_X1 U580 ( .A(KEYINPUT113), .B(KEYINPUT42), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U582 ( .A(G57GAT), .B(n518), .ZN(G1332GAT) );
  NOR2_X1 U583 ( .A1(n523), .A2(n529), .ZN(n519) );
  XOR2_X1 U584 ( .A(KEYINPUT114), .B(n519), .Z(n520) );
  XNOR2_X1 U585 ( .A(G64GAT), .B(n520), .ZN(G1333GAT) );
  NOR2_X1 U586 ( .A1(n523), .A2(n567), .ZN(n522) );
  XNOR2_X1 U587 ( .A(G71GAT), .B(KEYINPUT115), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n522), .B(n521), .ZN(G1334GAT) );
  XNOR2_X1 U589 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n525) );
  NOR2_X1 U590 ( .A1(n537), .A2(n523), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n525), .B(n524), .ZN(G1335GAT) );
  NAND2_X1 U592 ( .A1(n527), .A2(n526), .ZN(n536) );
  NOR2_X1 U593 ( .A1(n584), .A2(n536), .ZN(n528) );
  XOR2_X1 U594 ( .A(G85GAT), .B(n528), .Z(G1336GAT) );
  NOR2_X1 U595 ( .A1(n529), .A2(n536), .ZN(n530) );
  XOR2_X1 U596 ( .A(KEYINPUT116), .B(n530), .Z(n531) );
  XNOR2_X1 U597 ( .A(G92GAT), .B(n531), .ZN(G1337GAT) );
  NOR2_X1 U598 ( .A1(n567), .A2(n536), .ZN(n533) );
  XNOR2_X1 U599 ( .A(G99GAT), .B(KEYINPUT117), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n533), .B(n532), .ZN(G1338GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n535) );
  XNOR2_X1 U602 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n534) );
  XNOR2_X1 U603 ( .A(n535), .B(n534), .ZN(n539) );
  NOR2_X1 U604 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U605 ( .A(n539), .B(n538), .Z(G1339GAT) );
  NOR2_X1 U606 ( .A1(n567), .A2(n551), .ZN(n540) );
  NAND2_X1 U607 ( .A1(n541), .A2(n540), .ZN(n548) );
  NOR2_X1 U608 ( .A1(n554), .A2(n548), .ZN(n542) );
  XOR2_X1 U609 ( .A(G113GAT), .B(n542), .Z(G1340GAT) );
  INV_X1 U610 ( .A(n543), .ZN(n557) );
  NOR2_X1 U611 ( .A1(n557), .A2(n548), .ZN(n545) );
  XNOR2_X1 U612 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(G1341GAT) );
  NOR2_X1 U614 ( .A1(n561), .A2(n548), .ZN(n546) );
  XOR2_X1 U615 ( .A(KEYINPUT50), .B(n546), .Z(n547) );
  XNOR2_X1 U616 ( .A(G127GAT), .B(n547), .ZN(G1342GAT) );
  NOR2_X1 U617 ( .A1(n564), .A2(n548), .ZN(n550) );
  XNOR2_X1 U618 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n549) );
  XNOR2_X1 U619 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  NOR2_X1 U620 ( .A1(n584), .A2(n551), .ZN(n552) );
  NAND2_X1 U621 ( .A1(n553), .A2(n552), .ZN(n563) );
  NOR2_X1 U622 ( .A1(n554), .A2(n563), .ZN(n555) );
  XOR2_X1 U623 ( .A(KEYINPUT122), .B(n555), .Z(n556) );
  XNOR2_X1 U624 ( .A(G141GAT), .B(n556), .ZN(G1344GAT) );
  NOR2_X1 U625 ( .A1(n557), .A2(n563), .ZN(n559) );
  XNOR2_X1 U626 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U628 ( .A(G148GAT), .B(n560), .ZN(G1345GAT) );
  NOR2_X1 U629 ( .A1(n561), .A2(n563), .ZN(n562) );
  XOR2_X1 U630 ( .A(G155GAT), .B(n562), .Z(G1346GAT) );
  NOR2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U632 ( .A(G162GAT), .B(n565), .Z(G1347GAT) );
  NOR2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n569) );
  NAND2_X1 U634 ( .A1(n569), .A2(n574), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n568), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U636 ( .A1(n582), .A2(n569), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n570), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n572) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n571) );
  XNOR2_X1 U640 ( .A(n572), .B(n571), .ZN(n576) );
  NAND2_X1 U641 ( .A1(n587), .A2(n584), .ZN(n573) );
  NOR2_X1 U642 ( .A1(n586), .A2(n573), .ZN(n581) );
  NAND2_X1 U643 ( .A1(n581), .A2(n574), .ZN(n575) );
  XOR2_X1 U644 ( .A(n576), .B(n575), .Z(G1352GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n579) );
  NAND2_X1 U646 ( .A1(n577), .A2(n581), .ZN(n578) );
  XNOR2_X1 U647 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U648 ( .A(G204GAT), .B(n580), .ZN(G1353GAT) );
  NAND2_X1 U649 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n583), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U651 ( .A(n584), .ZN(n585) );
  NOR2_X1 U652 ( .A1(n586), .A2(n585), .ZN(n588) );
  NOR2_X1 U653 ( .A1(n589), .A2(n293), .ZN(n590) );
  XOR2_X1 U654 ( .A(KEYINPUT62), .B(n590), .Z(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

