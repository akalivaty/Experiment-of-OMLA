//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 1 1 1 0 0 0 1 0 0 1 1 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n970, new_n971, new_n972;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT90), .ZN(new_n203));
  NAND2_X1  g002(.A1(G71gat), .A2(G78gat), .ZN(new_n204));
  OR2_X1    g003(.A1(G71gat), .A2(G78gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT9), .ZN(new_n206));
  OR2_X1    g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n203), .B1(new_n204), .B2(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(new_n205), .B(KEYINPUT89), .Z(new_n209));
  INV_X1    g008(.A(KEYINPUT88), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n210), .B(new_n204), .C1(new_n202), .C2(new_n206), .ZN(new_n211));
  NAND4_X1  g010(.A1(new_n202), .A2(KEYINPUT88), .A3(G71gat), .A4(G78gat), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n209), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n208), .A2(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n214), .A2(KEYINPUT21), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n215), .B(G127gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(G231gat), .A2(G233gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n216), .B(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(G15gat), .B(G22gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT16), .ZN(new_n220));
  AOI21_X1  g019(.A(G1gat), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  XOR2_X1   g020(.A(new_n221), .B(G8gat), .Z(new_n222));
  NAND2_X1  g021(.A1(new_n219), .A2(KEYINPUT85), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n222), .B(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT21), .ZN(new_n225));
  INV_X1    g024(.A(new_n214), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  XOR2_X1   g026(.A(KEYINPUT91), .B(G155gat), .Z(new_n228));
  XNOR2_X1  g027(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n218), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n231));
  XNOR2_X1  g030(.A(G183gat), .B(G211gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n230), .B(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT14), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n235), .B1(G29gat), .B2(G36gat), .ZN(new_n236));
  NOR2_X1   g035(.A1(G29gat), .A2(G36gat), .ZN(new_n237));
  MUX2_X1   g036(.A(new_n236), .B(new_n235), .S(new_n237), .Z(new_n238));
  XNOR2_X1  g037(.A(G43gat), .B(G50gat), .ZN(new_n239));
  AOI22_X1  g038(.A1(new_n238), .A2(KEYINPUT84), .B1(KEYINPUT15), .B2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n238), .B1(KEYINPUT15), .B2(new_n239), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(KEYINPUT17), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT94), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT93), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT7), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(G85gat), .ZN(new_n248));
  INV_X1    g047(.A(G92gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n247), .B(new_n250), .C1(new_n244), .C2(new_n246), .ZN(new_n253));
  NAND2_X1  g052(.A1(G99gat), .A2(G106gat), .ZN(new_n254));
  AOI22_X1  g053(.A1(KEYINPUT8), .A2(new_n254), .B1(new_n248), .B2(new_n249), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT95), .ZN(new_n256));
  AND2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n255), .A2(new_n256), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n252), .B(new_n253), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G99gat), .B(G106gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n260), .B(KEYINPUT96), .ZN(new_n261));
  OAI21_X1  g060(.A(KEYINPUT97), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  OR2_X1    g061(.A1(new_n255), .A2(new_n256), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n255), .A2(new_n256), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n251), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n260), .B(KEYINPUT96), .Z(new_n266));
  INV_X1    g065(.A(KEYINPUT97), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n265), .A2(new_n266), .A3(new_n267), .A4(new_n253), .ZN(new_n268));
  AOI22_X1  g067(.A1(new_n262), .A2(new_n268), .B1(new_n261), .B2(new_n259), .ZN(new_n269));
  OR2_X1    g068(.A1(new_n243), .A2(new_n269), .ZN(new_n270));
  XOR2_X1   g069(.A(G190gat), .B(G218gat), .Z(new_n271));
  NAND3_X1  g070(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n262), .A2(new_n268), .ZN(new_n273));
  INV_X1    g072(.A(new_n259), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n273), .B1(new_n266), .B2(new_n274), .ZN(new_n275));
  OR2_X1    g074(.A1(new_n275), .A2(new_n242), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n270), .A2(new_n271), .A3(new_n272), .A4(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT98), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(KEYINPUT92), .ZN(new_n280));
  XNOR2_X1  g079(.A(G134gat), .B(G162gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n270), .A2(new_n272), .A3(new_n276), .ZN(new_n284));
  INV_X1    g083(.A(new_n271), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(new_n277), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n283), .B(new_n287), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n234), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n275), .A2(new_n226), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n259), .A2(KEYINPUT99), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n263), .A2(new_n264), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT99), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n292), .A2(new_n293), .A3(new_n252), .A4(new_n253), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n291), .A2(new_n294), .A3(new_n261), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n273), .A2(new_n295), .A3(new_n214), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n290), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(G230gat), .A2(G233gat), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT10), .ZN(new_n301));
  NOR3_X1   g100(.A1(new_n275), .A2(new_n301), .A3(new_n226), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n296), .B(new_n301), .C1(new_n269), .C2(new_n214), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT100), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n290), .A2(KEYINPUT100), .A3(new_n301), .A4(new_n296), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n302), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n300), .B1(new_n307), .B2(new_n299), .ZN(new_n308));
  XNOR2_X1  g107(.A(G120gat), .B(G148gat), .ZN(new_n309));
  INV_X1    g108(.A(G176gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n309), .B(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G204gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n308), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n313), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n300), .B(new_n315), .C1(new_n307), .C2(new_n299), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT101), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n314), .A2(KEYINPUT101), .A3(new_n316), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n289), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT87), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT36), .ZN(new_n326));
  INV_X1    g125(.A(G190gat), .ZN(new_n327));
  AND2_X1   g126(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G183gat), .A2(G190gat), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT67), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT24), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT24), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n331), .A2(new_n332), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n330), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT25), .ZN(new_n338));
  NAND2_X1  g137(.A1(G169gat), .A2(G176gat), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT66), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n339), .B(new_n340), .ZN(new_n341));
  NOR2_X1   g140(.A1(G169gat), .A2(G176gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT23), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT65), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n344), .B1(new_n342), .B2(KEYINPUT23), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT23), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n346), .B(KEYINPUT65), .C1(G169gat), .C2(G176gat), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n341), .A2(new_n343), .A3(new_n345), .A4(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(KEYINPUT69), .B1(new_n338), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT25), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n327), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n351));
  INV_X1    g150(.A(G183gat), .ZN(new_n352));
  OAI21_X1  g151(.A(G190gat), .B1(new_n335), .B2(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n351), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n350), .B1(new_n348), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n345), .A2(new_n347), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n339), .A2(new_n340), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n343), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT69), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n361), .A2(new_n362), .A3(KEYINPUT25), .A4(new_n337), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n349), .A2(new_n356), .A3(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT28), .ZN(new_n365));
  OR2_X1    g164(.A1(new_n328), .A2(new_n329), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT27), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n365), .B(new_n327), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT27), .B(G183gat), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n365), .B1(new_n371), .B2(new_n327), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n372), .B1(G183gat), .B2(G190gat), .ZN(new_n373));
  INV_X1    g172(.A(new_n341), .ZN(new_n374));
  XOR2_X1   g173(.A(new_n342), .B(KEYINPUT26), .Z(new_n375));
  OAI211_X1 g174(.A(new_n370), .B(new_n373), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n364), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G113gat), .B(G120gat), .ZN(new_n378));
  OAI21_X1  g177(.A(G127gat), .B1(new_n378), .B2(KEYINPUT1), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT1), .ZN(new_n380));
  INV_X1    g179(.A(G127gat), .ZN(new_n381));
  INV_X1    g180(.A(G113gat), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n382), .A2(G120gat), .ZN(new_n383));
  INV_X1    g182(.A(G120gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n384), .A2(G113gat), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n380), .B(new_n381), .C1(new_n383), .C2(new_n385), .ZN(new_n386));
  AND3_X1   g185(.A1(new_n379), .A2(G134gat), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(G134gat), .B1(new_n379), .B2(new_n386), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT70), .ZN(new_n389));
  NOR3_X1   g188(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(G134gat), .ZN(new_n391));
  NOR3_X1   g190(.A1(new_n378), .A2(KEYINPUT1), .A3(G127gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n384), .A2(G113gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n382), .A2(G120gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n381), .B1(new_n395), .B2(new_n380), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n391), .B1(new_n392), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n379), .A2(G134gat), .A3(new_n386), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT70), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n390), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(KEYINPUT71), .B1(new_n377), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n377), .A2(new_n400), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n389), .B1(new_n387), .B2(new_n388), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n397), .A2(KEYINPUT70), .A3(new_n398), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT71), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n405), .A2(new_n406), .A3(new_n364), .A4(new_n376), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n401), .A2(new_n402), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(G227gat), .A2(G233gat), .ZN(new_n409));
  XOR2_X1   g208(.A(new_n409), .B(KEYINPUT64), .Z(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(G15gat), .B(G43gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n412), .B(G71gat), .ZN(new_n413));
  XOR2_X1   g212(.A(new_n413), .B(G99gat), .Z(new_n414));
  XOR2_X1   g213(.A(KEYINPUT72), .B(KEYINPUT33), .Z(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT32), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT73), .B1(new_n411), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT73), .ZN(new_n420));
  AOI211_X1 g219(.A(new_n420), .B(new_n417), .C1(new_n408), .C2(new_n410), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n410), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n401), .A2(new_n423), .A3(new_n402), .A4(new_n407), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n424), .B(KEYINPUT34), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n415), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n411), .B1(KEYINPUT32), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n414), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n422), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n426), .B1(new_n422), .B2(new_n429), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n326), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT75), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n419), .ZN(new_n435));
  INV_X1    g234(.A(new_n421), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n429), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(new_n425), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n426), .A3(new_n429), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n440), .A2(KEYINPUT75), .A3(new_n326), .ZN(new_n441));
  AND2_X1   g240(.A1(new_n425), .A2(KEYINPUT74), .ZN(new_n442));
  OR2_X1    g241(.A1(new_n437), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n437), .A2(new_n442), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(KEYINPUT36), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n434), .A2(new_n441), .A3(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(G211gat), .B(G218gat), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT76), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n447), .B(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n450));
  INV_X1    g249(.A(G197gat), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n312), .ZN(new_n452));
  NAND2_X1  g251(.A1(G197gat), .A2(G204gat), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n450), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  XOR2_X1   g253(.A(new_n449), .B(new_n454), .Z(new_n455));
  NAND2_X1  g254(.A1(G155gat), .A2(G162gat), .ZN(new_n456));
  INV_X1    g255(.A(G155gat), .ZN(new_n457));
  INV_X1    g256(.A(G162gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(G141gat), .B(G148gat), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n456), .B(new_n459), .C1(new_n460), .C2(KEYINPUT2), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT3), .ZN(new_n462));
  INV_X1    g261(.A(G141gat), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(G148gat), .ZN(new_n464));
  INV_X1    g263(.A(G148gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(G141gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n459), .A2(new_n456), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n456), .A2(KEYINPUT2), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n461), .A2(new_n462), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT29), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n455), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n449), .B(new_n454), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT3), .B1(new_n475), .B2(new_n472), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n470), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n474), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(G228gat), .A2(G233gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n480), .B(G22gat), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  OR2_X1    g281(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT81), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n479), .A2(new_n482), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(KEYINPUT31), .B(G50gat), .ZN(new_n487));
  OR2_X1    g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(G78gat), .B(G106gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n486), .A2(new_n487), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n489), .B1(new_n488), .B2(new_n490), .ZN(new_n492));
  OR2_X1    g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  XOR2_X1   g292(.A(G8gat), .B(G36gat), .Z(new_n494));
  XNOR2_X1  g293(.A(new_n494), .B(G64gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(new_n249), .ZN(new_n496));
  INV_X1    g295(.A(G226gat), .ZN(new_n497));
  INV_X1    g296(.A(G233gat), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n499), .A2(KEYINPUT29), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT77), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n377), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n364), .A2(KEYINPUT77), .A3(new_n376), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n501), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n364), .A2(new_n499), .A3(new_n376), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n455), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n503), .A2(new_n499), .A3(new_n504), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n377), .A2(new_n500), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(new_n475), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n508), .A2(KEYINPUT37), .A3(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT83), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n508), .A2(new_n511), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT37), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AOI211_X1 g315(.A(KEYINPUT83), .B(KEYINPUT37), .C1(new_n508), .C2(new_n511), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n496), .B(new_n512), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT38), .ZN(new_n519));
  NOR3_X1   g318(.A1(new_n505), .A2(new_n455), .A3(new_n507), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n475), .B1(new_n509), .B2(new_n510), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT38), .B1(new_n522), .B2(KEYINPUT37), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n523), .B(new_n496), .C1(new_n516), .C2(new_n517), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT79), .ZN(new_n525));
  NOR3_X1   g324(.A1(new_n387), .A2(new_n388), .A3(new_n477), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT4), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n478), .A2(new_n397), .A3(new_n398), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n529), .A2(KEYINPUT79), .A3(KEYINPUT4), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  AOI211_X1 g330(.A(KEYINPUT4), .B(new_n477), .C1(new_n403), .C2(new_n404), .ZN(new_n532));
  OAI21_X1  g331(.A(KEYINPUT80), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n477), .A2(KEYINPUT3), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n534), .B(new_n471), .C1(new_n387), .C2(new_n388), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT78), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n535), .A2(new_n536), .ZN(new_n538));
  OR2_X1    g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n405), .A2(new_n527), .A3(new_n478), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT80), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n540), .A2(new_n541), .A3(new_n528), .A4(new_n530), .ZN(new_n542));
  NAND2_X1  g341(.A1(G225gat), .A2(G233gat), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n544), .A2(KEYINPUT5), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n533), .A2(new_n539), .A3(new_n542), .A4(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n477), .B1(new_n387), .B2(new_n388), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(new_n529), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(new_n544), .ZN(new_n549));
  OAI22_X1  g348(.A1(new_n537), .A2(new_n538), .B1(KEYINPUT4), .B2(new_n526), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n405), .A2(KEYINPUT4), .A3(new_n478), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(new_n543), .ZN(new_n552));
  OAI211_X1 g351(.A(KEYINPUT5), .B(new_n549), .C1(new_n550), .C2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n546), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G1gat), .B(G29gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT0), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(G57gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(new_n248), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT6), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n546), .A2(new_n553), .A3(new_n558), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n554), .A2(KEYINPUT6), .A3(new_n559), .ZN(new_n564));
  AND2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n496), .ZN(new_n566));
  AND3_X1   g365(.A1(new_n509), .A2(new_n475), .A3(new_n510), .ZN(new_n567));
  AND3_X1   g366(.A1(new_n364), .A2(KEYINPUT77), .A3(new_n376), .ZN(new_n568));
  AOI21_X1  g367(.A(KEYINPUT77), .B1(new_n364), .B2(new_n376), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n500), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n475), .B1(new_n570), .B2(new_n506), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n566), .B1(new_n567), .B2(new_n571), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n519), .A2(new_n524), .A3(new_n565), .A4(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT39), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n548), .A2(new_n544), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n533), .A2(new_n539), .A3(new_n542), .ZN(new_n576));
  AOI211_X1 g375(.A(new_n574), .B(new_n575), .C1(new_n576), .C2(new_n544), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n576), .A2(new_n574), .A3(new_n544), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(new_n558), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT40), .ZN(new_n580));
  NOR3_X1   g379(.A1(new_n577), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n508), .A2(new_n496), .A3(new_n511), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n572), .A2(KEYINPUT30), .A3(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT30), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n514), .A2(new_n584), .A3(new_n566), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n580), .B1(new_n577), .B2(new_n579), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT82), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI211_X1 g389(.A(KEYINPUT82), .B(new_n580), .C1(new_n577), .C2(new_n579), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n587), .A2(new_n560), .A3(new_n590), .A4(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n493), .B1(new_n573), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n491), .A2(new_n492), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n563), .A2(new_n564), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(new_n586), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n446), .B1(new_n593), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n596), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n599), .A2(new_n594), .A3(new_n443), .A4(new_n444), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT35), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n493), .A2(new_n440), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n596), .A2(KEYINPUT35), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n598), .A2(new_n605), .ZN(new_n606));
  OR2_X1    g405(.A1(new_n224), .A2(new_n242), .ZN(new_n607));
  NAND2_X1  g406(.A1(G229gat), .A2(G233gat), .ZN(new_n608));
  INV_X1    g407(.A(new_n224), .ZN(new_n609));
  OAI211_X1 g408(.A(new_n607), .B(new_n608), .C1(new_n243), .C2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT18), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n224), .B(new_n242), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n608), .B(KEYINPUT13), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n610), .A2(new_n611), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n612), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G113gat), .B(G141gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(G197gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT11), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(G169gat), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n622), .B(KEYINPUT12), .Z(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n618), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n612), .A2(new_n617), .A3(new_n623), .A4(new_n616), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT86), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n626), .A2(new_n627), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n625), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n325), .B1(new_n606), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n631), .ZN(new_n633));
  AOI211_X1 g432(.A(KEYINPUT87), .B(new_n633), .C1(new_n598), .C2(new_n605), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n324), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT102), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI22_X1  g436(.A1(new_n600), .A2(KEYINPUT35), .B1(new_n602), .B2(new_n603), .ZN(new_n638));
  INV_X1    g437(.A(new_n597), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n591), .A2(new_n560), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n576), .A2(new_n544), .ZN(new_n641));
  INV_X1    g440(.A(new_n575), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n641), .A2(KEYINPUT39), .A3(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n643), .A2(new_n558), .A3(new_n578), .ZN(new_n644));
  AOI21_X1  g443(.A(KEYINPUT82), .B1(new_n644), .B2(new_n580), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n640), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n514), .A2(new_n515), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(KEYINPUT83), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n514), .A2(new_n513), .A3(new_n515), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n566), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n595), .B1(new_n650), .B2(new_n523), .ZN(new_n651));
  INV_X1    g450(.A(new_n572), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n652), .B1(new_n518), .B2(KEYINPUT38), .ZN(new_n653));
  AOI22_X1  g452(.A1(new_n646), .A2(new_n587), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n639), .B1(new_n654), .B2(new_n493), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n638), .B1(new_n655), .B2(new_n446), .ZN(new_n656));
  OAI21_X1  g455(.A(KEYINPUT87), .B1(new_n656), .B2(new_n633), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n606), .A2(new_n325), .A3(new_n631), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n659), .A2(KEYINPUT102), .A3(new_n324), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n637), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(new_n565), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g462(.A(KEYINPUT42), .B(G8gat), .Z(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n586), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n661), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n665), .B1(new_n667), .B2(new_n220), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n661), .A2(KEYINPUT16), .A3(new_n666), .A4(new_n664), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT42), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n668), .A2(new_n669), .A3(new_n671), .ZN(G1325gat));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n446), .A2(KEYINPUT103), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT103), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n434), .A2(new_n441), .A3(new_n675), .A4(new_n445), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(KEYINPUT102), .B1(new_n659), .B2(new_n324), .ZN(new_n678));
  AOI211_X1 g477(.A(new_n636), .B(new_n323), .C1(new_n657), .C2(new_n658), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(G15gat), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n440), .A2(G15gat), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n682), .B1(new_n678), .B2(new_n679), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n673), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n674), .A2(new_n676), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n685), .B1(new_n637), .B2(new_n660), .ZN(new_n686));
  INV_X1    g485(.A(G15gat), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n683), .B(new_n673), .C1(new_n686), .C2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n684), .A2(new_n689), .ZN(G1326gat));
  NAND2_X1  g489(.A1(new_n661), .A2(new_n493), .ZN(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT43), .B(G22gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n638), .B1(new_n685), .B2(new_n655), .ZN(new_n695));
  INV_X1    g494(.A(new_n288), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n694), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n234), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n698), .A2(new_n321), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n700), .A2(new_n633), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n606), .A2(KEYINPUT44), .A3(new_n288), .ZN(new_n702));
  AND3_X1   g501(.A1(new_n697), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(new_n565), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(G29gat), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n659), .A2(new_n288), .A3(new_n699), .ZN(new_n706));
  OR3_X1    g505(.A1(new_n706), .A2(G29gat), .A3(new_n595), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n707), .A2(KEYINPUT45), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n707), .A2(KEYINPUT45), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n705), .B1(new_n708), .B2(new_n709), .ZN(G1328gat));
  NOR2_X1   g509(.A1(new_n586), .A2(G36gat), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  OR3_X1    g511(.A1(new_n706), .A2(KEYINPUT46), .A3(new_n712), .ZN(new_n713));
  AOI211_X1 g512(.A(new_n694), .B(new_n696), .C1(new_n598), .C2(new_n605), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n573), .A2(new_n592), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n597), .B1(new_n715), .B2(new_n594), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n716), .B1(new_n674), .B2(new_n676), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n288), .B1(new_n717), .B2(new_n638), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n714), .B1(new_n718), .B2(new_n694), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n719), .A2(KEYINPUT105), .A3(new_n666), .A4(new_n701), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n697), .A2(new_n666), .A3(new_n701), .A4(new_n702), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT105), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n720), .A2(new_n723), .A3(G36gat), .ZN(new_n724));
  OAI21_X1  g523(.A(KEYINPUT46), .B1(new_n706), .B2(new_n712), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n713), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(KEYINPUT106), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT106), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n713), .A2(new_n724), .A3(new_n728), .A4(new_n725), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(G1329gat));
  INV_X1    g529(.A(G43gat), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n731), .B1(new_n706), .B2(new_n440), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n703), .A2(G43gat), .A3(new_n677), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT107), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(KEYINPUT47), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n732), .A2(new_n733), .A3(new_n735), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n734), .A2(KEYINPUT47), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1330gat));
  NAND3_X1  g537(.A1(new_n703), .A2(G50gat), .A3(new_n493), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n706), .A2(new_n594), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(G50gat), .B2(new_n740), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g541(.A1(new_n695), .A2(new_n631), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n322), .A2(new_n234), .A3(new_n288), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n565), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g547(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n746), .A2(new_n666), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT108), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT108), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n746), .A2(new_n752), .A3(new_n666), .A4(new_n749), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(G1333gat));
  OAI21_X1  g555(.A(G71gat), .B1(new_n745), .B2(new_n685), .ZN(new_n757));
  OR2_X1    g556(.A1(new_n745), .A2(G71gat), .ZN(new_n758));
  XOR2_X1   g557(.A(new_n440), .B(KEYINPUT109), .Z(new_n759));
  OAI21_X1  g558(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n760), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n493), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(G78gat), .ZN(G1335gat));
  INV_X1    g562(.A(KEYINPUT112), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n565), .A2(new_n248), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT111), .B1(new_n695), .B2(new_n696), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT111), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n767), .B(new_n288), .C1(new_n717), .C2(new_n638), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n633), .A2(new_n234), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n766), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n766), .A2(new_n768), .A3(KEYINPUT51), .A4(new_n770), .ZN(new_n774));
  AOI211_X1 g573(.A(new_n322), .B(new_n765), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT110), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n769), .A2(new_n322), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n719), .A2(new_n776), .A3(new_n565), .A4(new_n777), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n697), .A2(new_n565), .A3(new_n702), .A4(new_n777), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(KEYINPUT110), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n778), .A2(new_n780), .A3(G85gat), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n764), .B1(new_n775), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n778), .A2(new_n780), .A3(G85gat), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n773), .A2(new_n774), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n321), .ZN(new_n785));
  OAI211_X1 g584(.A(KEYINPUT112), .B(new_n783), .C1(new_n785), .C2(new_n765), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n782), .A2(new_n786), .ZN(G1336gat));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n771), .A2(new_n788), .A3(new_n772), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n772), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n766), .A2(new_n768), .A3(new_n770), .A4(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n322), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n586), .A2(G92gat), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n719), .A2(new_n666), .A3(new_n777), .ZN(new_n794));
  AOI22_X1  g593(.A1(new_n792), .A2(new_n793), .B1(G92gat), .B2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n784), .A2(new_n321), .A3(new_n793), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n794), .A2(G92gat), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n796), .ZN(new_n799));
  OAI22_X1  g598(.A1(new_n795), .A2(new_n796), .B1(new_n797), .B2(new_n799), .ZN(G1337gat));
  AND2_X1   g599(.A1(new_n719), .A2(new_n777), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n801), .A2(KEYINPUT114), .A3(new_n677), .ZN(new_n802));
  XNOR2_X1  g601(.A(KEYINPUT115), .B(G99gat), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT114), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n719), .A2(new_n777), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n804), .B1(new_n805), .B2(new_n685), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n802), .A2(new_n803), .A3(new_n806), .ZN(new_n807));
  OR2_X1    g606(.A1(new_n440), .A2(new_n803), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n807), .B1(new_n785), .B2(new_n808), .ZN(G1338gat));
  INV_X1    g608(.A(G106gat), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n810), .B1(new_n801), .B2(new_n493), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n321), .A2(new_n810), .A3(new_n493), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n812), .B1(new_n789), .B2(new_n791), .ZN(new_n813));
  OAI21_X1  g612(.A(KEYINPUT53), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  OR2_X1    g613(.A1(new_n811), .A2(KEYINPUT53), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n812), .B1(new_n773), .B2(new_n774), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(G1339gat));
  NOR2_X1   g616(.A1(new_n666), .A2(new_n595), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n607), .B1(new_n243), .B2(new_n609), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n820), .A2(G229gat), .A3(G233gat), .ZN(new_n821));
  OR2_X1    g620(.A1(new_n613), .A2(new_n615), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n622), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OR2_X1    g622(.A1(new_n626), .A2(new_n627), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n823), .B1(new_n824), .B2(new_n628), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n288), .B1(new_n825), .B2(new_n321), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n827), .B1(new_n307), .B2(new_n299), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n305), .A2(new_n306), .ZN(new_n829));
  INV_X1    g628(.A(new_n302), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n298), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n828), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n299), .B1(new_n829), .B2(new_n830), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n315), .B1(new_n834), .B2(new_n827), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n833), .A2(new_n835), .A3(KEYINPUT55), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n833), .A2(new_n835), .A3(KEYINPUT116), .A4(KEYINPUT55), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(KEYINPUT55), .B1(new_n833), .B2(new_n835), .ZN(new_n841));
  INV_X1    g640(.A(new_n316), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n840), .A2(new_n631), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n826), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n840), .A2(new_n825), .A3(new_n843), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n288), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n847), .A3(new_n234), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n289), .A2(new_n633), .A3(new_n322), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n819), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n850), .A2(new_n602), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n382), .B1(new_n851), .B2(new_n631), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT117), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n594), .A2(new_n443), .A3(new_n444), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n856), .A2(new_n382), .A3(new_n631), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n853), .A2(new_n857), .ZN(G1340gat));
  INV_X1    g657(.A(new_n851), .ZN(new_n859));
  OAI21_X1  g658(.A(G120gat), .B1(new_n859), .B2(new_n322), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n856), .A2(new_n384), .A3(new_n321), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(G1341gat));
  AOI21_X1  g661(.A(G127gat), .B1(new_n856), .B2(new_n698), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n234), .A2(new_n381), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n863), .B1(new_n851), .B2(new_n864), .ZN(G1342gat));
  NAND3_X1  g664(.A1(new_n856), .A2(new_n391), .A3(new_n288), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n866), .A2(KEYINPUT56), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n867), .A2(KEYINPUT118), .ZN(new_n868));
  OR2_X1    g667(.A1(new_n866), .A2(KEYINPUT56), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(KEYINPUT118), .ZN(new_n870));
  OAI21_X1  g669(.A(G134gat), .B1(new_n859), .B2(new_n696), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n868), .A2(new_n869), .A3(new_n870), .A4(new_n871), .ZN(G1343gat));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n685), .A2(new_n818), .ZN(new_n874));
  OR2_X1    g673(.A1(new_n874), .A2(KEYINPUT119), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(KEYINPUT119), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n594), .B1(new_n848), .B2(new_n849), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(KEYINPUT57), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n878), .A2(KEYINPUT57), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n877), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(G141gat), .B1(new_n882), .B2(new_n633), .ZN(new_n883));
  AOI211_X1 g682(.A(new_n594), .B(new_n874), .C1(new_n849), .C2(new_n848), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n884), .A2(new_n463), .A3(new_n631), .ZN(new_n885));
  AOI211_X1 g684(.A(new_n873), .B(KEYINPUT58), .C1(new_n883), .C2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT58), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(KEYINPUT120), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT58), .ZN(new_n889));
  AND4_X1   g688(.A1(new_n888), .A2(new_n883), .A3(new_n889), .A4(new_n885), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n886), .A2(new_n890), .ZN(G1344gat));
  OAI21_X1  g690(.A(G148gat), .B1(new_n882), .B2(new_n322), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI211_X1 g693(.A(KEYINPUT121), .B(G148gat), .C1(new_n882), .C2(new_n322), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n894), .A2(KEYINPUT59), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n884), .A2(new_n465), .A3(new_n321), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n892), .A2(new_n893), .A3(new_n898), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n896), .A2(new_n897), .A3(new_n899), .ZN(G1345gat));
  AOI21_X1  g699(.A(G155gat), .B1(new_n884), .B2(new_n698), .ZN(new_n901));
  INV_X1    g700(.A(new_n882), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n234), .A2(new_n457), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(G1346gat));
  AOI21_X1  g703(.A(G162gat), .B1(new_n884), .B2(new_n288), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n696), .A2(new_n458), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n905), .B1(new_n902), .B2(new_n906), .ZN(G1347gat));
  NAND2_X1  g706(.A1(new_n848), .A2(new_n849), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n565), .A2(new_n586), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(new_n855), .A3(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(G169gat), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n911), .A2(new_n912), .A3(new_n631), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n759), .A2(new_n493), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n908), .A2(new_n909), .A3(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n908), .A2(KEYINPUT122), .A3(new_n909), .A4(new_n915), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(new_n631), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n914), .B1(new_n921), .B2(G169gat), .ZN(new_n922));
  AOI211_X1 g721(.A(KEYINPUT123), .B(new_n912), .C1(new_n920), .C2(new_n631), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n913), .B1(new_n922), .B2(new_n923), .ZN(G1348gat));
  NAND4_X1  g723(.A1(new_n918), .A2(G176gat), .A3(new_n321), .A4(new_n919), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT124), .ZN(new_n926));
  OR2_X1    g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n310), .B1(new_n910), .B2(new_n322), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n925), .A2(new_n926), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(KEYINPUT125), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT125), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n927), .A2(new_n932), .A3(new_n928), .A4(new_n929), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(G1349gat));
  NAND3_X1  g733(.A1(new_n918), .A2(new_n698), .A3(new_n919), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT126), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(new_n366), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n918), .A2(KEYINPUT126), .A3(new_n698), .A4(new_n919), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n911), .A2(new_n371), .A3(new_n698), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(KEYINPUT60), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT60), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n940), .A2(new_n944), .A3(new_n941), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(new_n945), .ZN(G1350gat));
  NAND3_X1  g745(.A1(new_n911), .A2(new_n327), .A3(new_n288), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT61), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n920), .A2(new_n288), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n948), .B1(new_n949), .B2(G190gat), .ZN(new_n950));
  AOI211_X1 g749(.A(KEYINPUT61), .B(new_n327), .C1(new_n920), .C2(new_n288), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n947), .B1(new_n950), .B2(new_n951), .ZN(G1351gat));
  INV_X1    g751(.A(new_n881), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(new_n879), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n685), .A2(new_n909), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g755(.A(G197gat), .B1(new_n956), .B2(new_n633), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n878), .A2(new_n955), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n631), .A2(new_n451), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(G1352gat));
  OAI21_X1  g759(.A(G204gat), .B1(new_n956), .B2(new_n322), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n958), .A2(G204gat), .A3(new_n322), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n962), .B(KEYINPUT62), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n961), .A2(new_n963), .ZN(G1353gat));
  OR3_X1    g763(.A1(new_n958), .A2(G211gat), .A3(new_n234), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n954), .A2(new_n698), .A3(new_n955), .ZN(new_n966));
  AND3_X1   g765(.A1(new_n966), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n967));
  AOI21_X1  g766(.A(KEYINPUT63), .B1(new_n966), .B2(G211gat), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n965), .B1(new_n967), .B2(new_n968), .ZN(G1354gat));
  NOR3_X1   g768(.A1(new_n958), .A2(G218gat), .A3(new_n696), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n954), .A2(new_n288), .A3(new_n955), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n970), .B1(new_n971), .B2(G218gat), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


