//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 1 1 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 0 1 0 1 0 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 1 1 0 0 0 1 1 0 0 1 0 0 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n776, new_n777, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  NAND3_X1  g001(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT79), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT22), .B(G137), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G128), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G119), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n193), .B(KEYINPUT74), .ZN(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G128), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT75), .ZN(new_n197));
  XNOR2_X1  g011(.A(new_n196), .B(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(KEYINPUT24), .B(G110), .ZN(new_n199));
  NOR3_X1   g013(.A1(new_n194), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT23), .B1(new_n192), .B2(G119), .ZN(new_n201));
  AOI21_X1  g015(.A(KEYINPUT76), .B1(new_n192), .B2(G119), .ZN(new_n202));
  XNOR2_X1  g016(.A(new_n201), .B(new_n202), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n200), .B1(G110), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G140), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G125), .ZN(new_n206));
  INV_X1    g020(.A(G125), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G140), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT77), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n206), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(KEYINPUT77), .A3(G140), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(KEYINPUT16), .A3(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT16), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n206), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n212), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT78), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT78), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n212), .A2(new_n218), .A3(new_n213), .A4(new_n215), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n212), .A2(new_n215), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G146), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n217), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n204), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n199), .B1(new_n194), .B2(new_n198), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n224), .B1(G110), .B2(new_n203), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n213), .B1(new_n212), .B2(new_n215), .ZN(new_n226));
  AND3_X1   g040(.A1(new_n206), .A2(new_n208), .A3(new_n213), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  AND3_X1   g043(.A1(new_n223), .A2(KEYINPUT80), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(KEYINPUT80), .B1(new_n223), .B2(new_n229), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n191), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n191), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n223), .A2(new_n229), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n233), .B1(new_n234), .B2(KEYINPUT80), .ZN(new_n235));
  INV_X1    g049(.A(G234), .ZN(new_n236));
  AOI21_X1  g050(.A(G902), .B1(new_n236), .B2(G217), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n232), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT81), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT81), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n232), .A2(new_n235), .A3(new_n240), .A4(new_n237), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G902), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n232), .A2(new_n243), .A3(new_n235), .ZN(new_n244));
  OR2_X1    g058(.A1(new_n244), .A2(KEYINPUT25), .ZN(new_n245));
  OAI21_X1  g059(.A(G217), .B1(new_n236), .B2(G902), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n246), .B1(new_n244), .B2(KEYINPUT25), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n242), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  XOR2_X1   g063(.A(KEYINPUT2), .B(G113), .Z(new_n250));
  NAND2_X1  g064(.A1(new_n195), .A2(G116), .ZN(new_n251));
  INV_X1    g065(.A(G116), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G119), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n250), .A2(new_n251), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n251), .A2(new_n253), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT2), .B(G113), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n192), .A2(KEYINPUT1), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n213), .A2(G143), .ZN(new_n261));
  INV_X1    g075(.A(G143), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G146), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n260), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n264), .A2(KEYINPUT66), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT66), .ZN(new_n266));
  XNOR2_X1  g080(.A(G143), .B(G146), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n266), .B1(new_n267), .B2(new_n260), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n262), .A2(G146), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT64), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n263), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n262), .A2(KEYINPUT64), .A3(G146), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n269), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n192), .B1(new_n261), .B2(KEYINPUT1), .ZN(new_n274));
  OAI22_X1  g088(.A1(new_n265), .A2(new_n268), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G137), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT65), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT65), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G137), .ZN(new_n279));
  AND2_X1   g093(.A1(KEYINPUT11), .A2(G134), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n277), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G131), .ZN(new_n282));
  NAND2_X1  g096(.A1(KEYINPUT11), .A2(G134), .ZN(new_n283));
  NOR2_X1   g097(.A1(KEYINPUT11), .A2(G134), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n283), .B1(new_n284), .B2(G137), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n281), .A2(new_n282), .A3(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G134), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n277), .A2(new_n279), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n282), .B1(G134), .B2(G137), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n275), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n281), .A2(new_n285), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G131), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n286), .ZN(new_n295));
  AND3_X1   g109(.A1(new_n262), .A2(KEYINPUT64), .A3(G146), .ZN(new_n296));
  AOI21_X1  g110(.A(KEYINPUT64), .B1(new_n262), .B2(G146), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n261), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  AND2_X1   g112(.A1(KEYINPUT0), .A2(G128), .ZN(new_n299));
  NOR2_X1   g113(.A1(KEYINPUT0), .A2(G128), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI22_X1  g115(.A1(new_n298), .A2(new_n301), .B1(new_n267), .B2(new_n299), .ZN(new_n302));
  AOI22_X1  g116(.A1(new_n292), .A2(KEYINPUT67), .B1(new_n295), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT67), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n275), .A2(new_n291), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n259), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n267), .A2(new_n266), .A3(new_n260), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n264), .A2(KEYINPUT66), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT1), .ZN(new_n309));
  OAI21_X1  g123(.A(G128), .B1(new_n269), .B2(new_n309), .ZN(new_n310));
  AOI22_X1  g124(.A1(new_n307), .A2(new_n308), .B1(new_n298), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n286), .A2(new_n290), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT69), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT69), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n275), .A2(new_n291), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n295), .A2(new_n302), .ZN(new_n316));
  AND4_X1   g130(.A1(new_n259), .A2(new_n313), .A3(new_n315), .A4(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT28), .B1(new_n306), .B2(new_n317), .ZN(new_n318));
  NOR2_X1   g132(.A1(G237), .A2(G953), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G210), .ZN(new_n320));
  XOR2_X1   g134(.A(new_n320), .B(KEYINPUT27), .Z(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT26), .B(G101), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n321), .B(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n316), .A2(new_n292), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT70), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT70), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n316), .A2(new_n292), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n326), .A2(new_n259), .A3(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT28), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n318), .A2(new_n324), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT29), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT67), .B1(new_n311), .B2(new_n312), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(new_n305), .A3(new_n316), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT30), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT68), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n292), .A2(KEYINPUT69), .B1(new_n295), .B2(new_n302), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(KEYINPUT30), .A3(new_n315), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT68), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n336), .A2(new_n342), .A3(new_n337), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n339), .A2(new_n258), .A3(new_n341), .A4(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n340), .A2(new_n259), .A3(new_n315), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n324), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n334), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n331), .A2(KEYINPUT72), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n259), .B1(new_n340), .B2(new_n315), .ZN(new_n349));
  OAI21_X1  g163(.A(KEYINPUT28), .B1(new_n349), .B2(new_n317), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT72), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n329), .A2(new_n351), .A3(new_n330), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n323), .A2(new_n333), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n348), .A2(new_n350), .A3(new_n352), .A4(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n243), .ZN(new_n355));
  OAI21_X1  g169(.A(G472), .B1(new_n347), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(G472), .A2(G902), .ZN(new_n357));
  XOR2_X1   g171(.A(new_n357), .B(KEYINPUT71), .Z(new_n358));
  INV_X1    g172(.A(KEYINPUT32), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n344), .A2(new_n324), .A3(new_n345), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n361), .A2(KEYINPUT31), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT31), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n344), .A2(new_n363), .A3(new_n324), .A4(new_n345), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n318), .A2(new_n331), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n323), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n360), .B1(new_n362), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n356), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n361), .A2(KEYINPUT31), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n370), .A2(new_n366), .A3(new_n364), .ZN(new_n371));
  INV_X1    g185(.A(new_n358), .ZN(new_n372));
  AOI21_X1  g186(.A(KEYINPUT32), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(KEYINPUT73), .B1(new_n369), .B2(new_n373), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n243), .B(new_n354), .C1(new_n334), .C2(new_n346), .ZN(new_n375));
  AOI22_X1  g189(.A1(new_n371), .A2(new_n360), .B1(new_n375), .B2(G472), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n372), .B1(new_n362), .B2(new_n367), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n359), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT73), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n376), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n249), .B1(new_n374), .B2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(G110), .B(G122), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G107), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n384), .A2(G104), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(KEYINPUT83), .A3(G104), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n385), .B1(KEYINPUT3), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT3), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n388), .A2(new_n384), .A3(KEYINPUT83), .A4(G104), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT4), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n391), .A3(G101), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n258), .ZN(new_n393));
  INV_X1    g207(.A(G101), .ZN(new_n394));
  AOI211_X1 g208(.A(KEYINPUT84), .B(new_n394), .C1(new_n387), .C2(new_n389), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n386), .A2(KEYINPUT3), .ZN(new_n396));
  INV_X1    g210(.A(G104), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G107), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n396), .A2(new_n394), .A3(new_n389), .A4(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(KEYINPUT4), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT84), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n402), .B1(new_n390), .B2(G101), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n393), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n251), .A2(new_n253), .A3(KEYINPUT5), .ZN(new_n406));
  OAI21_X1  g220(.A(G113), .B1(new_n251), .B2(KEYINPUT5), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n254), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n397), .A2(G107), .ZN(new_n409));
  OAI21_X1  g223(.A(G101), .B1(new_n409), .B2(new_n385), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n399), .A2(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n383), .B1(new_n405), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n412), .ZN(new_n414));
  NOR3_X1   g228(.A1(new_n403), .A2(new_n395), .A3(new_n400), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n382), .B(new_n414), .C1(new_n415), .C2(new_n393), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n413), .A2(KEYINPUT6), .A3(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT6), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n418), .B(new_n383), .C1(new_n405), .C2(new_n412), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n311), .A2(new_n207), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n298), .A2(new_n301), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n267), .A2(new_n299), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G125), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n187), .A2(G224), .ZN(new_n426));
  XOR2_X1   g240(.A(new_n425), .B(new_n426), .Z(new_n427));
  NAND3_X1  g241(.A1(new_n417), .A2(new_n419), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT88), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n408), .A2(new_n411), .A3(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n382), .B(KEYINPUT8), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n408), .A2(new_n411), .ZN(new_n432));
  OAI21_X1  g246(.A(KEYINPUT88), .B1(new_n408), .B2(new_n411), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n430), .B(new_n431), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n426), .A2(KEYINPUT7), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n425), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n420), .A2(new_n424), .A3(KEYINPUT7), .A4(new_n426), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n434), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(G902), .B1(new_n438), .B2(new_n416), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n428), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(G210), .B1(G237), .B2(G902), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n441), .B(KEYINPUT89), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n442), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n428), .A2(new_n439), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n443), .A2(KEYINPUT90), .A3(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(G214), .B1(G237), .B2(G902), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT90), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n440), .A2(new_n448), .A3(new_n442), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n446), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(G113), .B(G122), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n451), .B(new_n397), .ZN(new_n452));
  INV_X1    g266(.A(G237), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n453), .A2(new_n187), .A3(G214), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n262), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n319), .A2(G143), .A3(G214), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G131), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT17), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n455), .A2(new_n282), .A3(new_n456), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n457), .A2(KEYINPUT17), .A3(G131), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OR2_X1    g277(.A1(new_n222), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n211), .ZN(new_n465));
  XNOR2_X1  g279(.A(G125), .B(G140), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n465), .B1(new_n209), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n227), .B1(new_n467), .B2(G146), .ZN(new_n468));
  NAND2_X1  g282(.A1(KEYINPUT18), .A2(G131), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n454), .A2(new_n262), .ZN(new_n471));
  AOI21_X1  g285(.A(G143), .B1(new_n319), .B2(G214), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n455), .A2(new_n456), .A3(new_n469), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OR2_X1    g289(.A1(new_n468), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n452), .B1(new_n464), .B2(new_n476), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n452), .B(new_n476), .C1(new_n222), .C2(new_n463), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n243), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(G475), .ZN(new_n481));
  INV_X1    g295(.A(G952), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n482), .A2(G953), .ZN(new_n483));
  NAND2_X1  g297(.A1(G234), .A2(G237), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(KEYINPUT21), .B(G898), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n484), .A2(G902), .A3(G953), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n485), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n468), .A2(new_n475), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n210), .A2(KEYINPUT19), .A3(new_n211), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT19), .ZN(new_n492));
  AOI21_X1  g306(.A(KEYINPUT91), .B1(new_n466), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n210), .A2(KEYINPUT91), .A3(KEYINPUT19), .A4(new_n211), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n213), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n220), .A2(G146), .B1(new_n458), .B2(new_n460), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n490), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT92), .B1(new_n499), .B2(new_n452), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n458), .A2(new_n460), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n221), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(G146), .B1(new_n494), .B2(new_n495), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n476), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT92), .ZN(new_n505));
  INV_X1    g319(.A(new_n452), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n500), .A2(new_n507), .A3(new_n478), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT20), .ZN(new_n509));
  NOR2_X1   g323(.A1(G475), .A2(G902), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n509), .B1(new_n508), .B2(new_n510), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n481), .B(new_n489), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT9), .B(G234), .ZN(new_n515));
  INV_X1    g329(.A(G217), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n515), .A2(new_n516), .A3(G953), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT97), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT96), .ZN(new_n520));
  INV_X1    g334(.A(G122), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n520), .B(KEYINPUT14), .C1(new_n521), .C2(G116), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(G116), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n252), .A2(G122), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n520), .B1(new_n525), .B2(KEYINPUT14), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n519), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  OR2_X1    g341(.A1(new_n525), .A2(KEYINPUT14), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT14), .B1(new_n521), .B2(G116), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT96), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n530), .A2(KEYINPUT97), .A3(new_n523), .A4(new_n522), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n527), .A2(new_n528), .A3(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT98), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n532), .A2(new_n533), .A3(G107), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n533), .B1(new_n532), .B2(G107), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n523), .A2(new_n525), .A3(new_n384), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n262), .A2(G128), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n192), .A2(G143), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT95), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n537), .A2(new_n538), .A3(KEYINPUT95), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(G134), .A3(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(G134), .B1(new_n541), .B2(new_n542), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n536), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR3_X1   g360(.A1(new_n534), .A2(new_n535), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n545), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n523), .A2(new_n525), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(G107), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n536), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n192), .A2(G143), .ZN(new_n553));
  OAI21_X1  g367(.A(KEYINPUT93), .B1(new_n553), .B2(KEYINPUT13), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT93), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT13), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n537), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n554), .A2(new_n538), .A3(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT94), .ZN(new_n559));
  OR2_X1    g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n558), .A2(new_n559), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n553), .A2(KEYINPUT13), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n552), .B1(new_n563), .B2(G134), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n518), .B1(new_n547), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT99), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n532), .A2(G107), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(KEYINPUT98), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n532), .A2(new_n533), .A3(G107), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n548), .A2(new_n543), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n568), .A2(new_n536), .A3(new_n569), .A4(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n561), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n562), .B1(new_n558), .B2(new_n559), .ZN(new_n573));
  OAI21_X1  g387(.A(G134), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n574), .A2(new_n548), .A3(new_n551), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n571), .A2(new_n575), .A3(new_n517), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n565), .A2(new_n566), .A3(new_n576), .ZN(new_n577));
  OAI211_X1 g391(.A(KEYINPUT99), .B(new_n518), .C1(new_n547), .C2(new_n564), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(new_n243), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(G478), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(KEYINPUT15), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n581), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n577), .A2(new_n243), .A3(new_n578), .A4(new_n583), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n514), .A2(KEYINPUT100), .A3(new_n582), .A4(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT100), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n582), .A2(new_n584), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n586), .B1(new_n587), .B2(new_n513), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n450), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(G221), .B1(new_n515), .B2(G902), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(KEYINPUT82), .ZN(new_n591));
  INV_X1    g405(.A(G469), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n592), .A2(new_n243), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n392), .A2(new_n302), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n390), .A2(new_n402), .A3(G101), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n595), .A2(KEYINPUT4), .A3(new_n399), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n594), .B1(new_n596), .B2(new_n403), .ZN(new_n597));
  INV_X1    g411(.A(new_n295), .ZN(new_n598));
  OAI22_X1  g412(.A1(new_n265), .A2(new_n268), .B1(new_n267), .B2(new_n274), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n599), .A2(new_n399), .A3(new_n410), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT10), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n275), .A2(KEYINPUT10), .A3(new_n399), .A4(new_n410), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n597), .A2(new_n598), .A3(new_n602), .A4(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(G110), .B(G140), .ZN(new_n605));
  AND2_X1   g419(.A1(new_n187), .A2(G227), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n604), .A2(KEYINPUT87), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(KEYINPUT87), .B1(new_n604), .B2(new_n608), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n311), .A2(new_n411), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n600), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT12), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n598), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT85), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n308), .A2(new_n307), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n298), .A2(new_n310), .ZN(new_n619));
  AND3_X1   g433(.A1(new_n411), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n267), .ZN(new_n621));
  AOI22_X1  g435(.A1(new_n308), .A2(new_n307), .B1(new_n621), .B2(new_n310), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n622), .A2(new_n411), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n617), .B1(new_n620), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n600), .A2(new_n612), .A3(KEYINPUT85), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n624), .A2(new_n625), .A3(new_n295), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n626), .A2(KEYINPUT86), .A3(new_n614), .ZN(new_n627));
  AOI21_X1  g441(.A(KEYINPUT86), .B1(new_n626), .B2(new_n614), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n616), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n611), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n597), .A2(new_n602), .A3(new_n603), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n295), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n604), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n607), .ZN(new_n634));
  AOI21_X1  g448(.A(G902), .B1(new_n630), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n593), .B1(new_n635), .B2(new_n592), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n632), .A2(new_n608), .A3(new_n604), .ZN(new_n637));
  INV_X1    g451(.A(new_n604), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n626), .A2(new_n614), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT86), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n626), .A2(KEYINPUT86), .A3(new_n614), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n638), .B1(new_n643), .B2(new_n616), .ZN(new_n644));
  OAI211_X1 g458(.A(G469), .B(new_n637), .C1(new_n644), .C2(new_n608), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n591), .B1(new_n636), .B2(new_n645), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n589), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n381), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT101), .B(G101), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G3));
  NAND2_X1  g464(.A1(new_n371), .A2(new_n243), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n651), .A2(G472), .B1(new_n372), .B2(new_n371), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n641), .A2(new_n642), .B1(new_n613), .B2(new_n615), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n604), .A2(new_n608), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT87), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n604), .A2(KEYINPUT87), .A3(new_n608), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n634), .B1(new_n654), .B2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n660), .A2(new_n592), .A3(new_n243), .ZN(new_n661));
  INV_X1    g475(.A(new_n593), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n661), .A2(new_n645), .A3(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n591), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n653), .A2(new_n249), .A3(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n447), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n667), .B1(new_n443), .B2(new_n445), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n489), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT33), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n577), .A2(new_n670), .A3(new_n578), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n565), .A2(KEYINPUT33), .A3(new_n576), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n580), .A2(G902), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n579), .A2(new_n580), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n481), .B1(new_n511), .B2(new_n512), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n669), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n666), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT34), .B(G104), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G6));
  OAI211_X1 g496(.A(new_n587), .B(new_n481), .C1(new_n512), .C2(new_n511), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n683), .A2(new_n669), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n666), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT35), .B(G107), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G9));
  NAND2_X1  g501(.A1(new_n585), .A2(new_n588), .ZN(new_n688));
  INV_X1    g502(.A(new_n450), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n688), .A2(new_n652), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n245), .A2(new_n247), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n191), .A2(KEYINPUT36), .ZN(new_n692));
  XOR2_X1   g506(.A(new_n234), .B(new_n692), .Z(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n237), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n663), .A2(new_n664), .A3(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n690), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT37), .B(G110), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G12));
  NAND2_X1  g514(.A1(new_n374), .A2(new_n380), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n443), .A2(new_n445), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  XOR2_X1   g517(.A(new_n485), .B(KEYINPUT102), .Z(new_n704));
  OAI21_X1  g518(.A(new_n704), .B1(G900), .B2(new_n488), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NOR4_X1   g520(.A1(new_n683), .A2(new_n667), .A3(new_n703), .A4(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n701), .A2(new_n697), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G128), .ZN(G30));
  XNOR2_X1  g523(.A(new_n705), .B(KEYINPUT39), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n646), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g525(.A(new_n711), .B(KEYINPUT40), .Z(new_n712));
  AND2_X1   g526(.A1(new_n344), .A2(new_n345), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n713), .A2(new_n323), .ZN(new_n714));
  OR2_X1    g528(.A1(new_n349), .A2(new_n317), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n243), .B1(new_n715), .B2(new_n324), .ZN(new_n716));
  OAI21_X1  g530(.A(G472), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n378), .A2(new_n368), .A3(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n446), .A2(new_n449), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(KEYINPUT38), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n587), .A2(new_n677), .A3(new_n447), .ZN(new_n722));
  NOR4_X1   g536(.A1(new_n719), .A2(new_n721), .A3(new_n695), .A4(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n712), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G143), .ZN(G45));
  AOI21_X1  g539(.A(new_n696), .B1(new_n374), .B2(new_n380), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n676), .A2(new_n677), .A3(new_n705), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT103), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n676), .A2(KEYINPUT103), .A3(new_n677), .A4(new_n705), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n729), .A2(new_n668), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(KEYINPUT104), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT104), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n729), .A2(new_n733), .A3(new_n668), .A4(new_n730), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n726), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G146), .ZN(G48));
  AOI22_X1  g550(.A1(new_n611), .A2(new_n629), .B1(new_n607), .B2(new_n633), .ZN(new_n737));
  OAI21_X1  g551(.A(G469), .B1(new_n737), .B2(G902), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n248), .A2(new_n664), .A3(new_n661), .A4(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n739), .B1(new_n374), .B2(new_n380), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n679), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT105), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT105), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n740), .A2(new_n743), .A3(new_n679), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(KEYINPUT41), .B(G113), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(G15));
  INV_X1    g561(.A(new_n739), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n701), .A2(new_n684), .A3(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT106), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n740), .A2(KEYINPUT106), .A3(new_n684), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G116), .ZN(G18));
  NAND4_X1  g568(.A1(new_n738), .A2(new_n661), .A3(new_n664), .A4(new_n668), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n691), .A2(new_n694), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n757), .A2(new_n688), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n701), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G119), .ZN(G21));
  NAND2_X1  g574(.A1(new_n352), .A2(new_n350), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n351), .B1(new_n329), .B2(new_n330), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n323), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT107), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n370), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n364), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n764), .B1(new_n370), .B2(new_n763), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n372), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n651), .A2(G472), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n768), .A2(new_n248), .A3(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n738), .A2(new_n661), .A3(new_n664), .A4(new_n489), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n771), .A2(new_n703), .A3(new_n722), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G122), .ZN(G24));
  AND2_X1   g588(.A1(new_n768), .A2(new_n769), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n729), .A2(new_n730), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n776), .A3(new_n757), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G125), .ZN(G27));
  AOI21_X1  g592(.A(new_n667), .B1(new_n446), .B2(new_n449), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n663), .A2(new_n779), .A3(new_n664), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n701), .A2(new_n248), .A3(new_n776), .A4(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT42), .ZN(new_n782));
  INV_X1    g596(.A(new_n356), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n364), .A2(new_n366), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n358), .B1(new_n784), .B2(new_n370), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n368), .B1(new_n785), .B2(KEYINPUT32), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n783), .B1(new_n786), .B2(KEYINPUT108), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT108), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n378), .A2(new_n788), .A3(new_n368), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n249), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n729), .A2(new_n730), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n663), .A2(new_n779), .A3(KEYINPUT42), .A4(new_n664), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  AOI22_X1  g607(.A1(new_n781), .A2(new_n782), .B1(new_n790), .B2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(new_n282), .ZN(G33));
  NOR2_X1   g609(.A1(new_n683), .A2(new_n706), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n381), .A2(new_n796), .A3(new_n780), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(new_n287), .ZN(G36));
  OAI21_X1  g612(.A(new_n637), .B1(new_n644), .B2(new_n608), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT45), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n592), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n801), .B1(new_n800), .B2(new_n799), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT46), .B1(new_n802), .B2(new_n662), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n803), .B1(new_n592), .B2(new_n635), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n802), .A2(KEYINPUT46), .A3(new_n662), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n591), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(new_n710), .ZN(new_n807));
  INV_X1    g621(.A(new_n779), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n677), .B(KEYINPUT109), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n676), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n677), .A2(KEYINPUT43), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  AOI22_X1  g626(.A1(new_n810), .A2(KEYINPUT43), .B1(new_n676), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n813), .A2(new_n653), .A3(new_n695), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT44), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n808), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n816), .B1(new_n815), .B2(new_n814), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n807), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(new_n276), .ZN(G39));
  NAND2_X1  g633(.A1(new_n804), .A2(new_n805), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(new_n664), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT47), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n806), .A2(KEYINPUT47), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR4_X1   g639(.A1(new_n701), .A2(new_n248), .A3(new_n791), .A4(new_n808), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(G140), .ZN(G42));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT111), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n758), .A2(new_n701), .B1(new_n770), .B2(new_n772), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n740), .A2(new_n743), .A3(new_n679), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n743), .B1(new_n740), .B2(new_n679), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n740), .A2(KEYINPUT106), .A3(new_n684), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT106), .B1(new_n740), .B2(new_n684), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n830), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  AOI22_X1  g652(.A1(new_n381), .A2(new_n647), .B1(new_n690), .B2(new_n697), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n696), .A2(new_n808), .ZN(new_n840));
  OR3_X1    g654(.A1(new_n587), .A2(new_n677), .A3(new_n706), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n841), .B1(new_n374), .B2(new_n380), .ZN(new_n842));
  AND4_X1   g656(.A1(new_n769), .A2(new_n768), .A3(new_n729), .A4(new_n730), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n840), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n683), .A2(new_n678), .ZN(new_n845));
  MUX2_X1   g659(.A(new_n683), .B(new_n845), .S(KEYINPUT112), .Z(new_n846));
  AND2_X1   g660(.A1(new_n689), .A2(new_n489), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n666), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n839), .A2(new_n844), .A3(new_n848), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n849), .A2(new_n794), .A3(new_n797), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT52), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n722), .A2(new_n703), .A3(new_n706), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n646), .A2(new_n718), .A3(new_n756), .A4(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n708), .A2(new_n777), .A3(new_n853), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n726), .A2(new_n732), .A3(new_n734), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n851), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n726), .A2(new_n707), .B1(new_n843), .B2(new_n757), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n857), .A2(KEYINPUT52), .A3(new_n735), .A4(new_n853), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n745), .A2(new_n753), .A3(KEYINPUT111), .A4(new_n831), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n838), .A2(new_n850), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n838), .A2(new_n850), .A3(new_n860), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n856), .A2(new_n858), .A3(KEYINPUT113), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT113), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n866), .B(new_n851), .C1(new_n854), .C2(new_n855), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n862), .B1(new_n864), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n863), .B1(KEYINPUT114), .B2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT114), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n871), .B(new_n862), .C1(new_n864), .C2(new_n868), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n829), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n834), .A2(new_n837), .A3(new_n862), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n874), .A2(new_n865), .A3(new_n850), .A4(new_n867), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n861), .A2(KEYINPUT115), .A3(new_n862), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT115), .B1(new_n861), .B2(new_n862), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n829), .B(new_n875), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(KEYINPUT116), .B1(new_n873), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n869), .A2(KEYINPUT114), .ZN(new_n881));
  INV_X1    g695(.A(new_n863), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n881), .A2(new_n872), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(KEYINPUT54), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT116), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n884), .A2(new_n885), .A3(new_n878), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n738), .A2(new_n661), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n591), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n823), .A2(new_n824), .A3(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n704), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n813), .A2(new_n890), .A3(new_n770), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n779), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n738), .A2(new_n661), .A3(new_n664), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n895), .A2(new_n447), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n891), .A2(new_n721), .A3(new_n896), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT50), .Z(new_n898));
  NAND2_X1  g712(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT51), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n808), .A2(new_n895), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n249), .A2(new_n485), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n719), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  OR3_X1    g718(.A1(new_n904), .A2(new_n677), .A3(new_n676), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n813), .A2(new_n890), .A3(new_n902), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT117), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n775), .A2(new_n695), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n907), .A2(KEYINPUT118), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT118), .B1(new_n907), .B2(new_n909), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n905), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OR2_X1    g726(.A1(new_n912), .A2(KEYINPUT119), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(KEYINPUT119), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n901), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n900), .B1(new_n899), .B2(new_n912), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n907), .A2(new_n790), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT48), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n483), .B1(new_n904), .B2(new_n678), .ZN(new_n919));
  INV_X1    g733(.A(new_n755), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n919), .B1(new_n920), .B2(new_n891), .ZN(new_n921));
  AND4_X1   g735(.A1(new_n915), .A2(new_n916), .A3(new_n918), .A4(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n880), .A2(new_n886), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n482), .A2(new_n187), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR4_X1   g739(.A1(new_n810), .A2(new_n249), .A3(new_n591), .A4(new_n667), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT110), .Z(new_n927));
  XNOR2_X1  g741(.A(new_n887), .B(KEYINPUT49), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n927), .A2(new_n719), .A3(new_n721), .A4(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n925), .A2(new_n929), .ZN(G75));
  NAND2_X1  g744(.A1(new_n861), .A2(new_n862), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT115), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n861), .A2(KEYINPUT115), .A3(new_n862), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n243), .B1(new_n935), .B2(new_n875), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n442), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT56), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n417), .A2(new_n419), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(new_n427), .ZN(new_n940));
  XOR2_X1   g754(.A(KEYINPUT120), .B(KEYINPUT55), .Z(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n937), .A2(new_n938), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n942), .B1(new_n937), .B2(new_n938), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n187), .A2(G952), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(G51));
  XNOR2_X1  g760(.A(new_n593), .B(KEYINPUT57), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n829), .B1(new_n935), .B2(new_n875), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n947), .B1(new_n948), .B2(new_n879), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n660), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n802), .B(KEYINPUT121), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n936), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n945), .B1(new_n950), .B2(new_n952), .ZN(G54));
  NAND3_X1  g767(.A1(new_n936), .A2(KEYINPUT58), .A3(G475), .ZN(new_n954));
  INV_X1    g768(.A(new_n508), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n954), .A2(new_n955), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n956), .A2(new_n957), .A3(new_n945), .ZN(G60));
  NAND2_X1  g772(.A1(new_n671), .A2(new_n672), .ZN(new_n959));
  NAND2_X1  g773(.A1(G478), .A2(G902), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT59), .Z(new_n961));
  NOR2_X1   g775(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n962), .B1(new_n948), .B2(new_n879), .ZN(new_n963));
  INV_X1    g777(.A(new_n945), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n961), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n884), .A2(new_n885), .A3(new_n878), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n885), .B1(new_n884), .B2(new_n878), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n965), .B1(new_n969), .B2(new_n959), .ZN(G63));
  NAND2_X1  g784(.A1(new_n935), .A2(new_n875), .ZN(new_n971));
  NAND2_X1  g785(.A1(G217), .A2(G902), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT122), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT60), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n232), .A2(new_n235), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n693), .B(KEYINPUT123), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n971), .A2(new_n974), .A3(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n977), .A2(new_n964), .A3(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT61), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n977), .A2(KEYINPUT61), .A3(new_n964), .A4(new_n979), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(G66));
  AOI21_X1  g798(.A(new_n187), .B1(new_n487), .B2(G224), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n838), .A2(new_n860), .A3(new_n848), .A4(new_n839), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n985), .B1(new_n986), .B2(new_n187), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n939), .B1(G898), .B2(new_n187), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n987), .B(new_n988), .Z(G69));
  AOI21_X1  g803(.A(new_n818), .B1(new_n825), .B2(new_n826), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n794), .A2(new_n797), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n857), .A2(new_n735), .ZN(new_n992));
  INV_X1    g806(.A(new_n722), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n790), .A2(new_n702), .A3(new_n993), .ZN(new_n994));
  OR2_X1    g808(.A1(new_n807), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n990), .A2(new_n991), .A3(new_n992), .A4(new_n995), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n996), .A2(G953), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n339), .A2(new_n341), .A3(new_n343), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT124), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(new_n496), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n1000), .B1(G900), .B2(G953), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n992), .A2(new_n724), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(KEYINPUT62), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n846), .A2(new_n381), .A3(new_n710), .A4(new_n780), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n990), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n1002), .A2(KEYINPUT62), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n187), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  AOI22_X1  g821(.A1(new_n997), .A2(new_n1001), .B1(new_n1007), .B2(new_n1000), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n187), .B1(G227), .B2(G900), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1009), .B(KEYINPUT125), .ZN(new_n1010));
  AND3_X1   g824(.A1(new_n1008), .A2(KEYINPUT126), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1009), .ZN(new_n1012));
  OR2_X1    g826(.A1(new_n1008), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(KEYINPUT126), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1011), .B1(new_n1013), .B2(new_n1014), .ZN(G72));
  NAND2_X1  g829(.A1(G472), .A2(G902), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1016), .B(KEYINPUT63), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1017), .B(KEYINPUT127), .ZN(new_n1018));
  OR2_X1    g832(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1018), .B1(new_n1019), .B2(new_n986), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1020), .A2(new_n714), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1018), .B1(new_n996), .B2(new_n986), .ZN(new_n1022));
  AND2_X1   g836(.A1(new_n713), .A2(new_n323), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n945), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  NOR3_X1   g839(.A1(new_n1023), .A2(new_n714), .A3(new_n1017), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1025), .B1(new_n883), .B2(new_n1026), .ZN(G57));
endmodule


