//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 0 0 0 0 0 1 1 1 0 1 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 0 0 0 0 0 0 0 0 1 1 1 1 0 0 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1119, new_n1120, new_n1121,
    new_n1122, new_n1123, new_n1124, new_n1125, new_n1126, new_n1127,
    new_n1128, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238;
  INV_X1    g0000(.A(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G58), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT0), .Z(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n212), .B1(new_n201), .B2(new_n213), .ZN(new_n214));
  AOI21_X1  g0014(.A(new_n214), .B1(G107), .B2(G264), .ZN(new_n215));
  XOR2_X1   g0015(.A(KEYINPUT64), .B(G244), .Z(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G77), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT65), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G50), .A2(G226), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n215), .A2(new_n217), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(new_n208), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT1), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(G58), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(new_n201), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n211), .B(new_n223), .C1(new_n226), .C2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G264), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G226), .B(G232), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n234), .B(new_n239), .Z(G358));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n243), .B(KEYINPUT68), .Z(new_n244));
  NAND2_X1  g0044(.A1(G68), .A2(G77), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n203), .A2(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n246), .B(KEYINPUT67), .Z(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n244), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(G200), .ZN(new_n251));
  INV_X1    g0051(.A(G1), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n252), .B1(G41), .B2(G45), .ZN(new_n253));
  INV_X1    g0053(.A(G274), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1698), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n260), .A2(G222), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT70), .ZN(new_n263));
  AND2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(new_n261), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G223), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(G77), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT70), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n260), .A2(new_n270), .A3(G222), .A4(new_n261), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n263), .A2(new_n268), .A3(new_n269), .A4(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n224), .B1(G33), .B2(G41), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n255), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(G41), .A2(G45), .ZN(new_n275));
  OAI21_X1  g0075(.A(KEYINPUT69), .B1(new_n275), .B2(G1), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT69), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n277), .B(new_n252), .C1(G41), .C2(G45), .ZN(new_n278));
  INV_X1    g0078(.A(new_n224), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G41), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n276), .A2(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G226), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n251), .B1(new_n274), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n274), .A2(G190), .A3(new_n282), .ZN(new_n285));
  OAI21_X1  g0085(.A(G20), .B1(new_n228), .B2(G50), .ZN(new_n286));
  INV_X1    g0086(.A(G150), .ZN(new_n287));
  NOR2_X1   g0087(.A1(G20), .A2(G33), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n225), .A2(G33), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT8), .B(G58), .ZN(new_n291));
  OAI221_X1 g0091(.A(new_n286), .B1(new_n287), .B2(new_n289), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n224), .ZN(new_n294));
  INV_X1    g0094(.A(G50), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n252), .A2(G20), .ZN(new_n296));
  INV_X1    g0096(.A(G13), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AOI22_X1  g0098(.A1(new_n292), .A2(new_n294), .B1(new_n295), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n294), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n296), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G50), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT9), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n304), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT9), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n284), .A2(new_n285), .A3(new_n306), .A4(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT10), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT76), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n284), .A2(new_n311), .A3(new_n285), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n309), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n308), .A2(new_n306), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n274), .A2(new_n282), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n283), .B1(new_n316), .B2(G190), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n314), .B(new_n317), .C1(new_n311), .C2(KEYINPUT10), .ZN(new_n318));
  OAI211_X1 g0118(.A(KEYINPUT71), .B(new_n304), .C1(new_n316), .C2(G169), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT71), .ZN(new_n320));
  AOI21_X1  g0120(.A(G169), .B1(new_n274), .B2(new_n282), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n320), .B1(new_n321), .B2(new_n307), .ZN(new_n322));
  XOR2_X1   g0122(.A(KEYINPUT72), .B(G179), .Z(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n316), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n319), .A2(new_n322), .A3(new_n325), .ZN(new_n326));
  AND3_X1   g0126(.A1(new_n313), .A2(new_n318), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT77), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n261), .A2(G232), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n260), .B(new_n329), .C1(new_n213), .C2(new_n261), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n330), .B(new_n273), .C1(G107), .C2(new_n260), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT73), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n281), .A2(new_n216), .ZN(new_n333));
  INV_X1    g0133(.A(new_n255), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AOI211_X1 g0135(.A(KEYINPUT73), .B(new_n255), .C1(new_n281), .C2(new_n216), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n331), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT74), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n331), .B(KEYINPUT74), .C1(new_n335), .C2(new_n336), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(G190), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n298), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n345), .A2(G77), .ZN(new_n346));
  OR2_X1    g0146(.A1(new_n289), .A2(KEYINPUT75), .ZN(new_n347));
  INV_X1    g0147(.A(new_n291), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n289), .A2(KEYINPUT75), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT15), .B(G87), .ZN(new_n351));
  OAI221_X1 g0151(.A(new_n350), .B1(new_n225), .B2(new_n202), .C1(new_n351), .C2(new_n290), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n346), .B1(new_n352), .B2(new_n294), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(new_n202), .B2(new_n301), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n355), .B1(new_n341), .B2(new_n251), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n344), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n341), .A2(new_n324), .ZN(new_n359));
  INV_X1    g0159(.A(G169), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n339), .A2(new_n360), .A3(new_n340), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n359), .A2(new_n354), .A3(new_n361), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n327), .A2(new_n328), .A3(new_n358), .A4(new_n362), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n313), .A2(new_n318), .A3(new_n326), .A4(new_n362), .ZN(new_n364));
  OAI21_X1  g0164(.A(KEYINPUT77), .B1(new_n364), .B2(new_n357), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n260), .A2(G226), .A3(new_n261), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n260), .A2(G232), .A3(G1698), .ZN(new_n368));
  NAND2_X1  g0168(.A1(G33), .A2(G97), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n255), .B1(new_n370), .B2(new_n273), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT13), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n281), .A2(G238), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n372), .B1(new_n371), .B2(new_n373), .ZN(new_n375));
  OAI21_X1  g0175(.A(G169), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT14), .ZN(new_n377));
  INV_X1    g0177(.A(new_n374), .ZN(new_n378));
  INV_X1    g0178(.A(new_n375), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n378), .A2(G179), .A3(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT14), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n381), .B(G169), .C1(new_n374), .C2(new_n375), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n377), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT78), .ZN(new_n384));
  OAI22_X1  g0184(.A1(new_n289), .A2(new_n295), .B1(new_n225), .B2(G68), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n290), .A2(new_n202), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n294), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n387), .B(KEYINPUT11), .ZN(new_n388));
  OR3_X1    g0188(.A1(new_n345), .A2(KEYINPUT12), .A3(G68), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT12), .B1(new_n345), .B2(G68), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n389), .A2(new_n390), .B1(G68), .B2(new_n302), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT78), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n377), .A2(new_n393), .A3(new_n380), .A4(new_n382), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n384), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n378), .A2(new_n379), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(G200), .ZN(new_n397));
  INV_X1    g0197(.A(new_n392), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n397), .B(new_n398), .C1(new_n343), .C2(new_n396), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT7), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(new_n260), .B2(G20), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n266), .A2(KEYINPUT7), .A3(new_n225), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n201), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G58), .A2(G68), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n225), .B1(new_n228), .B2(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(G159), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n289), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT16), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NOR4_X1   g0214(.A1(new_n405), .A2(new_n413), .A3(new_n410), .A4(new_n407), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n414), .A2(new_n294), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n255), .B1(new_n281), .B2(G232), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n279), .A2(new_n280), .ZN(new_n420));
  INV_X1    g0220(.A(G223), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n261), .ZN(new_n422));
  INV_X1    g0222(.A(G226), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(G1698), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n422), .B(new_n424), .C1(new_n264), .C2(new_n265), .ZN(new_n425));
  NAND2_X1  g0225(.A1(G33), .A2(G87), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n420), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n251), .B1(new_n419), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n425), .A2(new_n426), .ZN(new_n429));
  AOI21_X1  g0229(.A(KEYINPUT80), .B1(new_n429), .B2(new_n273), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT80), .ZN(new_n431));
  AOI211_X1 g0231(.A(new_n431), .B(new_n420), .C1(new_n425), .C2(new_n426), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n343), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n428), .B1(new_n419), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n345), .A2(new_n291), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(new_n302), .B2(new_n291), .ZN(new_n436));
  XNOR2_X1  g0236(.A(new_n436), .B(KEYINPUT79), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n417), .A2(new_n434), .A3(new_n438), .ZN(new_n439));
  XNOR2_X1  g0239(.A(new_n439), .B(KEYINPUT17), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n430), .A2(new_n432), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n418), .A2(new_n324), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT81), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n360), .B1(new_n419), .B2(new_n427), .ZN(new_n445));
  AOI211_X1 g0245(.A(new_n323), .B(new_n255), .C1(new_n281), .C2(G232), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT81), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n446), .B(new_n447), .C1(new_n430), .C2(new_n432), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n444), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT82), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT82), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n444), .A2(new_n448), .A3(new_n451), .A4(new_n445), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n417), .A2(new_n438), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT18), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n453), .A2(KEYINPUT18), .A3(new_n454), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n457), .A2(KEYINPUT83), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT83), .ZN(new_n460));
  AOI221_X4 g0260(.A(new_n456), .B1(new_n417), .B2(new_n438), .C1(new_n450), .C2(new_n452), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT18), .B1(new_n453), .B2(new_n454), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n441), .B1(new_n459), .B2(new_n463), .ZN(new_n464));
  AND3_X1   g0264(.A1(new_n366), .A2(new_n401), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT85), .ZN(new_n466));
  INV_X1    g0266(.A(G45), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n467), .A2(G1), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G274), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  XNOR2_X1  g0270(.A(KEYINPUT5), .B(G41), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(G257), .ZN(new_n474));
  AOI211_X1 g0274(.A(new_n474), .B(new_n273), .C1(new_n471), .C2(new_n468), .ZN(new_n475));
  INV_X1    g0275(.A(G250), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n476), .B1(new_n258), .B2(new_n259), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT4), .ZN(new_n478));
  OAI21_X1  g0278(.A(G1698), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G283), .ZN(new_n480));
  INV_X1    g0280(.A(G244), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n478), .B1(new_n266), .B2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n260), .A2(KEYINPUT4), .A3(G244), .A4(new_n261), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n479), .A2(new_n480), .A3(new_n482), .A4(new_n483), .ZN(new_n484));
  AOI211_X1 g0284(.A(new_n473), .B(new_n475), .C1(new_n484), .C2(new_n273), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n466), .B1(new_n485), .B2(new_n251), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n345), .A2(G97), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n345), .B(new_n300), .C1(G1), .C2(new_n257), .ZN(new_n488));
  INV_X1    g0288(.A(G97), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n403), .A2(new_n404), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(G107), .ZN(new_n492));
  INV_X1    g0292(.A(G107), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n493), .A2(KEYINPUT6), .A3(G97), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n489), .A2(new_n493), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(new_n205), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n494), .B1(new_n496), .B2(KEYINPUT6), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G20), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n288), .A2(G77), .ZN(new_n499));
  XNOR2_X1  g0299(.A(new_n499), .B(KEYINPUT84), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n492), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  AOI211_X1 g0301(.A(new_n487), .B(new_n490), .C1(new_n501), .C2(new_n294), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n484), .A2(new_n273), .ZN(new_n503));
  INV_X1    g0303(.A(new_n475), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n503), .A2(G190), .A3(new_n472), .A4(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n503), .A2(new_n472), .A3(new_n504), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n506), .A2(KEYINPUT85), .A3(G200), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n486), .A2(new_n502), .A3(new_n505), .A4(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT86), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n298), .A2(new_n493), .ZN(new_n511));
  XNOR2_X1  g0311(.A(new_n511), .B(KEYINPUT25), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n260), .A2(new_n225), .A3(G87), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT22), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT22), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n260), .A2(new_n515), .A3(new_n225), .A4(G87), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n225), .A2(G107), .ZN(new_n518));
  XNOR2_X1  g0318(.A(new_n518), .B(KEYINPUT23), .ZN(new_n519));
  INV_X1    g0319(.A(G116), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n257), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n225), .ZN(new_n522));
  AND4_X1   g0322(.A1(KEYINPUT24), .A2(new_n517), .A3(new_n519), .A4(new_n522), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n514), .A2(new_n516), .B1(new_n225), .B2(new_n521), .ZN(new_n524));
  AOI21_X1  g0324(.A(KEYINPUT24), .B1(new_n524), .B2(new_n519), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n512), .B1(new_n526), .B2(new_n294), .ZN(new_n527));
  INV_X1    g0327(.A(new_n488), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(G107), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n267), .A2(G257), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G294), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n477), .A2(new_n261), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n273), .B1(new_n471), .B2(new_n468), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n533), .A2(new_n273), .B1(G264), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n472), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G200), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n535), .A2(new_n472), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G190), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n527), .A2(new_n529), .A3(new_n537), .A4(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n487), .B1(new_n501), .B2(new_n294), .ZN(new_n541));
  INV_X1    g0341(.A(new_n490), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n506), .A2(new_n360), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n543), .B(new_n544), .C1(new_n323), .C2(new_n506), .ZN(new_n545));
  AND3_X1   g0345(.A1(new_n541), .A2(new_n542), .A3(new_n505), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n546), .A2(KEYINPUT86), .A3(new_n486), .A4(new_n507), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n510), .A2(new_n540), .A3(new_n545), .A4(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n260), .A2(G257), .A3(new_n261), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(KEYINPUT87), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n266), .A2(G303), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n260), .A2(G264), .A3(G1698), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT87), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n260), .A2(new_n553), .A3(G257), .A4(new_n261), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n550), .A2(new_n551), .A3(new_n552), .A4(new_n554), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n555), .A2(new_n273), .B1(G270), .B2(new_n534), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n360), .B1(new_n556), .B2(new_n472), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n298), .A2(new_n520), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n480), .B(new_n225), .C1(G33), .C2(new_n489), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n559), .B(new_n294), .C1(new_n225), .C2(G116), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT20), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n560), .A2(new_n561), .ZN(new_n563));
  OAI221_X1 g0363(.A(new_n558), .B1(new_n488), .B2(new_n520), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(KEYINPUT21), .B1(new_n557), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n555), .A2(new_n273), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n534), .A2(G270), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n566), .A2(new_n472), .A3(new_n567), .ZN(new_n568));
  AND4_X1   g0368(.A1(KEYINPUT21), .A2(new_n568), .A3(G169), .A4(new_n564), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n524), .A2(new_n519), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT24), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n524), .A2(KEYINPUT24), .A3(new_n519), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(new_n294), .A3(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n512), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n575), .A2(new_n529), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(G169), .B1(new_n535), .B2(new_n472), .ZN(new_n578));
  INV_X1    g0378(.A(G179), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n578), .B1(new_n579), .B2(new_n538), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n568), .A2(new_n579), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n564), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n568), .A2(G200), .ZN(new_n584));
  INV_X1    g0384(.A(new_n564), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n584), .B(new_n585), .C1(new_n343), .C2(new_n568), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n570), .A2(new_n581), .A3(new_n583), .A4(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(G250), .B1(new_n467), .B2(G1), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n420), .B1(new_n470), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n266), .B1(new_n481), .B2(G1698), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n213), .A2(new_n261), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n521), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n590), .B1(new_n593), .B2(new_n420), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n324), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(new_n360), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n260), .A2(new_n225), .A3(G68), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n369), .A2(new_n225), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n599), .B(KEYINPUT19), .C1(new_n206), .C2(G87), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n369), .A2(G20), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n598), .B(new_n600), .C1(KEYINPUT19), .C2(new_n601), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n602), .A2(new_n294), .B1(new_n298), .B2(new_n351), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(new_n488), .B2(new_n351), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n596), .A2(new_n597), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n528), .A2(G87), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n594), .A2(G200), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(new_n343), .B2(new_n594), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n605), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  NOR3_X1   g0411(.A1(new_n548), .A2(new_n587), .A3(new_n611), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n465), .A2(new_n612), .ZN(G372));
  NOR2_X1   g0413(.A1(new_n548), .A2(new_n611), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n570), .A2(new_n581), .A3(new_n583), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n611), .A2(new_n545), .ZN(new_n617));
  XNOR2_X1  g0417(.A(new_n617), .B(KEYINPUT26), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n616), .A2(new_n605), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n465), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n326), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n399), .A2(new_n354), .A3(new_n359), .A4(new_n361), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n395), .A2(new_n622), .ZN(new_n623));
  OAI22_X1  g0423(.A1(new_n623), .A2(new_n441), .B1(new_n462), .B2(new_n461), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n313), .A2(new_n318), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n621), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n620), .A2(new_n626), .ZN(G369));
  NAND2_X1  g0427(.A1(new_n570), .A2(new_n583), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n297), .A2(G20), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n252), .ZN(new_n630));
  OR2_X1    g0430(.A1(new_n630), .A2(KEYINPUT27), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(KEYINPUT27), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n631), .A2(G213), .A3(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(G343), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n564), .A2(new_n635), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n628), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n628), .A2(new_n636), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(new_n586), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g0439(.A(KEYINPUT88), .B(G330), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n577), .A2(new_n635), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n540), .A2(new_n643), .B1(new_n577), .B2(new_n580), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n581), .A2(new_n635), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT89), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n642), .A2(KEYINPUT89), .A3(new_n646), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n635), .B1(new_n570), .B2(new_n583), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n646), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n654), .A2(new_n645), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n651), .A2(new_n655), .ZN(G399));
  INV_X1    g0456(.A(new_n209), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n657), .A2(G41), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(G1), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(new_n229), .B2(new_n659), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n662), .B(KEYINPUT28), .ZN(new_n663));
  INV_X1    g0463(.A(new_n605), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n664), .B1(new_n614), .B2(new_n615), .ZN(new_n665));
  AOI211_X1 g0465(.A(KEYINPUT29), .B(new_n635), .C1(new_n665), .C2(new_n618), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT29), .ZN(new_n667));
  INV_X1    g0467(.A(new_n635), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n667), .B1(new_n619), .B2(new_n668), .ZN(new_n669));
  AND4_X1   g0469(.A1(new_n535), .A2(new_n595), .A3(new_n503), .A4(new_n504), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n582), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT30), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n538), .A2(new_n485), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n674), .A2(new_n568), .A3(new_n324), .A4(new_n594), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n670), .A2(new_n582), .A3(KEYINPUT30), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n673), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(KEYINPUT31), .B1(new_n677), .B2(new_n635), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n678), .B1(new_n612), .B2(new_n668), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n673), .A2(new_n675), .A3(KEYINPUT90), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n676), .ZN(new_n681));
  AOI21_X1  g0481(.A(KEYINPUT90), .B1(new_n673), .B2(new_n675), .ZN(new_n682));
  OAI211_X1 g0482(.A(KEYINPUT31), .B(new_n635), .C1(new_n681), .C2(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n641), .B1(new_n679), .B2(new_n683), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n666), .A2(new_n669), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n663), .B1(new_n685), .B2(G1), .ZN(G364));
  NAND2_X1  g0486(.A1(new_n629), .A2(G45), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n659), .A2(G1), .A3(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n657), .A2(new_n260), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(new_n467), .B2(new_n230), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(KEYINPUT92), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n692), .A2(KEYINPUT92), .ZN(new_n694));
  OAI211_X1 g0494(.A(new_n693), .B(new_n694), .C1(new_n249), .C2(new_n467), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n260), .A2(new_n209), .ZN(new_n696));
  XOR2_X1   g0496(.A(G355), .B(KEYINPUT91), .Z(new_n697));
  OAI221_X1 g0497(.A(new_n695), .B1(G116), .B2(new_n209), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(G13), .A2(G33), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G20), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n224), .B1(G20), .B2(new_n360), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g0503(.A(new_n703), .B(KEYINPUT93), .Z(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n698), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n225), .A2(new_n343), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n323), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(new_n251), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(G50), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n225), .A2(G190), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n251), .A2(G179), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G107), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n707), .A2(new_n712), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G87), .ZN(new_n718));
  NOR2_X1   g0518(.A1(G179), .A2(G200), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n711), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(G159), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(KEYINPUT32), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n710), .A2(new_n715), .A3(new_n718), .A4(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n323), .A2(new_n711), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G200), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(new_n202), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n225), .B1(new_n719), .B2(G190), .ZN(new_n729));
  OAI22_X1  g0529(.A1(new_n722), .A2(KEYINPUT32), .B1(new_n489), .B2(new_n729), .ZN(new_n730));
  NOR4_X1   g0530(.A1(new_n724), .A2(new_n728), .A3(new_n266), .A4(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n708), .A2(G200), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n725), .A2(new_n251), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  OAI221_X1 g0535(.A(new_n731), .B1(new_n227), .B2(new_n733), .C1(new_n201), .C2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(G303), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n266), .B1(new_n716), .B2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT94), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  AOI22_X1  g0540(.A1(G283), .A2(new_n714), .B1(new_n721), .B2(G329), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n738), .A2(new_n739), .ZN(new_n742));
  INV_X1    g0542(.A(G294), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n741), .B(new_n742), .C1(new_n743), .C2(new_n729), .ZN(new_n744));
  XNOR2_X1  g0544(.A(KEYINPUT33), .B(G317), .ZN(new_n745));
  AOI211_X1 g0545(.A(new_n740), .B(new_n744), .C1(new_n734), .C2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n709), .A2(G326), .ZN(new_n747));
  INV_X1    g0547(.A(G311), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n746), .B(new_n747), .C1(new_n748), .C2(new_n727), .ZN(new_n749));
  INV_X1    g0549(.A(G322), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n733), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n736), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT95), .ZN(new_n753));
  INV_X1    g0553(.A(new_n702), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n689), .B(new_n706), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n755), .B1(new_n639), .B2(new_n701), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n642), .A2(new_n689), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n639), .A2(new_n641), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(G396));
  AOI21_X1  g0560(.A(new_n635), .B1(new_n665), .B2(new_n618), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n362), .A2(new_n635), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n344), .A2(new_n356), .B1(new_n355), .B2(new_n668), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n762), .B1(new_n763), .B2(new_n362), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n761), .B(new_n765), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n766), .A2(new_n684), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n684), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n767), .A2(new_n688), .A3(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n709), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n520), .A2(new_n727), .B1(new_n770), .B2(new_n737), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(G283), .B2(new_n734), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT96), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n773), .B1(G311), .B2(new_n721), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n714), .A2(G87), .ZN(new_n775));
  INV_X1    g0575(.A(new_n729), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n732), .A2(G294), .B1(G97), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n266), .B1(new_n716), .B2(new_n493), .ZN(new_n778));
  XOR2_X1   g0578(.A(new_n778), .B(KEYINPUT97), .Z(new_n779));
  NAND4_X1  g0579(.A1(new_n774), .A2(new_n775), .A3(new_n777), .A4(new_n779), .ZN(new_n780));
  AOI22_X1  g0580(.A1(G143), .A2(new_n732), .B1(new_n726), .B2(G159), .ZN(new_n781));
  AOI22_X1  g0581(.A1(G137), .A2(new_n709), .B1(new_n734), .B2(G150), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n782), .A2(KEYINPUT98), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(KEYINPUT98), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n781), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  XOR2_X1   g0585(.A(new_n785), .B(KEYINPUT34), .Z(new_n786));
  AOI21_X1  g0586(.A(new_n786), .B1(G50), .B2(new_n717), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n714), .A2(G68), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n787), .B(new_n788), .C1(new_n227), .C2(new_n729), .ZN(new_n789));
  INV_X1    g0589(.A(G132), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n260), .B1(new_n720), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n780), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(new_n702), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n702), .A2(new_n699), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n202), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n765), .A2(new_n699), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n793), .A2(new_n689), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n769), .A2(new_n797), .ZN(G384));
  NOR4_X1   g0598(.A1(new_n548), .A2(new_n587), .A3(new_n611), .A4(new_n635), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n677), .A2(KEYINPUT31), .A3(new_n635), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR3_X1   g0601(.A1(new_n799), .A2(new_n678), .A3(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n398), .A2(new_n668), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AND3_X1   g0604(.A1(new_n395), .A2(new_n399), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n804), .B1(new_n395), .B2(new_n399), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n764), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n802), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n459), .A2(new_n463), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n440), .ZN(new_n810));
  INV_X1    g0610(.A(new_n633), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n454), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n455), .A2(new_n439), .A3(new_n812), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(KEYINPUT100), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n454), .B1(new_n453), .B2(new_n811), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT100), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n817), .A2(new_n818), .A3(new_n439), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n816), .A2(KEYINPUT37), .A3(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT37), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n815), .A2(KEYINPUT100), .A3(new_n821), .ZN(new_n822));
  AND2_X1   g0622(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(KEYINPUT38), .B1(new_n814), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n812), .B1(new_n809), .B2(new_n440), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n820), .A2(new_n822), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT38), .ZN(new_n827));
  NOR3_X1   g0627(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n808), .B1(new_n824), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT40), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n821), .B1(new_n817), .B2(KEYINPUT101), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(new_n815), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n461), .A2(new_n462), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n813), .B1(new_n834), .B2(new_n441), .ZN(new_n835));
  AOI21_X1  g0635(.A(KEYINPUT38), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  OAI211_X1 g0636(.A(KEYINPUT40), .B(new_n808), .C1(new_n828), .C2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n831), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n612), .A2(new_n668), .ZN(new_n839));
  INV_X1    g0639(.A(new_n678), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n839), .A2(new_n840), .A3(new_n800), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n465), .A2(new_n841), .ZN(new_n842));
  XOR2_X1   g0642(.A(new_n838), .B(new_n842), .Z(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n640), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT39), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n828), .B2(new_n836), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n814), .A2(KEYINPUT38), .A3(new_n823), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n827), .B1(new_n825), .B2(new_n826), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n847), .A2(KEYINPUT39), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n395), .A2(new_n635), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n846), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n761), .A2(new_n764), .ZN(new_n852));
  INV_X1    g0652(.A(new_n762), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n805), .A2(new_n806), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n854), .B(new_n856), .C1(new_n824), .C2(new_n828), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n834), .A2(new_n633), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n851), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n465), .B1(new_n666), .B2(new_n669), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n626), .ZN(new_n861));
  XOR2_X1   g0661(.A(new_n859), .B(new_n861), .Z(new_n862));
  XNOR2_X1  g0662(.A(new_n844), .B(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n252), .B2(new_n629), .ZN(new_n864));
  OAI211_X1 g0664(.A(G116), .B(new_n226), .C1(new_n497), .C2(KEYINPUT35), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n865), .B(KEYINPUT99), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n497), .A2(KEYINPUT35), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n868), .B(KEYINPUT36), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n406), .A2(G77), .ZN(new_n870));
  OAI22_X1  g0670(.A1(new_n229), .A2(new_n870), .B1(G50), .B2(new_n201), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n871), .A2(G1), .A3(new_n297), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n864), .A2(new_n869), .A3(new_n872), .ZN(G367));
  AOI22_X1  g0673(.A1(new_n726), .A2(G283), .B1(G107), .B2(new_n776), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT46), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(new_n716), .B2(new_n520), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n717), .A2(KEYINPUT46), .A3(G116), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n874), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n878), .B1(G303), .B2(new_n732), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n489), .B2(new_n713), .ZN(new_n880));
  AOI211_X1 g0680(.A(new_n260), .B(new_n880), .C1(G294), .C2(new_n734), .ZN(new_n881));
  INV_X1    g0681(.A(G317), .ZN(new_n882));
  OAI221_X1 g0682(.A(new_n881), .B1(new_n748), .B2(new_n770), .C1(new_n882), .C2(new_n720), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n709), .A2(G143), .B1(G77), .B2(new_n714), .ZN(new_n884));
  AOI22_X1  g0684(.A1(G58), .A2(new_n717), .B1(new_n721), .B2(G137), .ZN(new_n885));
  OAI221_X1 g0685(.A(new_n884), .B1(KEYINPUT105), .B2(new_n885), .C1(new_n201), .C2(new_n729), .ZN(new_n886));
  AOI211_X1 g0686(.A(new_n266), .B(new_n886), .C1(KEYINPUT105), .C2(new_n885), .ZN(new_n887));
  AOI22_X1  g0687(.A1(G50), .A2(new_n726), .B1(new_n734), .B2(G159), .ZN(new_n888));
  XOR2_X1   g0688(.A(new_n888), .B(KEYINPUT104), .Z(new_n889));
  OAI211_X1 g0689(.A(new_n887), .B(new_n889), .C1(new_n287), .C2(new_n733), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n883), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n891), .B(KEYINPUT47), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n702), .ZN(new_n893));
  OAI221_X1 g0693(.A(new_n705), .B1(new_n209), .B2(new_n351), .C1(new_n234), .C2(new_n691), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n607), .A2(new_n668), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n664), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n611), .B2(new_n895), .ZN(new_n897));
  INV_X1    g0697(.A(new_n701), .ZN(new_n898));
  OR2_X1    g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n893), .A2(new_n689), .A3(new_n894), .A4(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n687), .A2(G1), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n543), .A2(new_n635), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n510), .A2(new_n545), .A3(new_n547), .A4(new_n902), .ZN(new_n903));
  OR2_X1    g0703(.A1(new_n545), .A2(new_n668), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n655), .A2(KEYINPUT45), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT45), .B1(new_n655), .B2(new_n905), .ZN(new_n907));
  OR2_X1    g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT44), .B1(new_n655), .B2(new_n905), .ZN(new_n909));
  OR3_X1    g0709(.A1(new_n655), .A2(KEYINPUT44), .A3(new_n905), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n908), .A2(new_n651), .A3(new_n909), .A4(new_n910), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n910), .B(new_n909), .C1(new_n906), .C2(new_n907), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n649), .A2(new_n650), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n646), .A2(new_n652), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n654), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT103), .B1(new_n639), .B2(new_n641), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n917), .A2(new_n918), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n685), .B1(new_n915), .B2(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n658), .B(KEYINPUT41), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n901), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT42), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n654), .A2(new_n926), .A3(new_n905), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n927), .A2(KEYINPUT102), .ZN(new_n928));
  INV_X1    g0728(.A(new_n905), .ZN(new_n929));
  OAI21_X1  g0729(.A(KEYINPUT42), .B1(new_n653), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n545), .B1(new_n903), .B2(new_n581), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n668), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n927), .A2(KEYINPUT102), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n928), .A2(new_n930), .A3(new_n932), .A4(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n897), .A2(KEYINPUT43), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n651), .A2(new_n929), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n934), .B(new_n935), .C1(new_n651), .C2(new_n929), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n897), .A2(KEYINPUT43), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n940), .B(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n900), .B1(new_n925), .B2(new_n943), .ZN(G387));
  NAND2_X1  g0744(.A1(new_n685), .A2(new_n921), .ZN(new_n945));
  INV_X1    g0745(.A(new_n685), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n922), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n945), .A2(new_n658), .A3(new_n947), .ZN(new_n948));
  AOI22_X1  g0748(.A1(G311), .A2(new_n734), .B1(new_n709), .B2(G322), .ZN(new_n949));
  OAI221_X1 g0749(.A(new_n949), .B1(new_n737), .B2(new_n727), .C1(new_n882), .C2(new_n733), .ZN(new_n950));
  XOR2_X1   g0750(.A(KEYINPUT107), .B(KEYINPUT48), .Z(new_n951));
  XNOR2_X1  g0751(.A(new_n950), .B(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(G283), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n952), .B1(new_n953), .B2(new_n729), .C1(new_n743), .C2(new_n716), .ZN(new_n954));
  XOR2_X1   g0754(.A(KEYINPUT108), .B(KEYINPUT49), .Z(new_n955));
  XNOR2_X1  g0755(.A(new_n954), .B(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n260), .B1(new_n721), .B2(G326), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n956), .B(new_n957), .C1(new_n520), .C2(new_n713), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n727), .A2(new_n201), .B1(new_n489), .B2(new_n713), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n733), .A2(new_n295), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n716), .A2(new_n202), .ZN(new_n961));
  XNOR2_X1  g0761(.A(KEYINPUT106), .B(G150), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n720), .A2(new_n962), .ZN(new_n963));
  NOR4_X1   g0763(.A1(new_n959), .A2(new_n960), .A3(new_n961), .A4(new_n963), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n729), .A2(new_n351), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n734), .A2(new_n348), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n266), .B1(new_n709), .B2(G159), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n964), .A2(new_n965), .A3(new_n966), .A4(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n754), .B1(new_n958), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n291), .A2(G50), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT50), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n971), .A2(new_n467), .A3(new_n245), .A4(new_n660), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n691), .B1(new_n239), .B2(G45), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n696), .A2(new_n660), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n657), .A2(new_n493), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n704), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NOR3_X1   g0777(.A1(new_n969), .A2(new_n688), .A3(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n701), .B1(new_n644), .B2(new_n645), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n978), .A2(new_n979), .B1(new_n901), .B2(new_n921), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n948), .A2(new_n980), .ZN(G393));
  NAND2_X1  g0781(.A1(new_n243), .A2(new_n690), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n705), .B(new_n982), .C1(new_n489), .C2(new_n209), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n689), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT109), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n735), .A2(new_n737), .ZN(new_n986));
  AOI22_X1  g0786(.A1(G311), .A2(new_n732), .B1(new_n709), .B2(G317), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT52), .Z(new_n988));
  OAI21_X1  g0788(.A(new_n715), .B1(new_n750), .B2(new_n720), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n260), .B(new_n989), .C1(new_n726), .C2(G294), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n988), .B(new_n990), .C1(new_n953), .C2(new_n716), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n986), .B(new_n991), .C1(G116), .C2(new_n776), .ZN(new_n992));
  AOI22_X1  g0792(.A1(G150), .A2(new_n709), .B1(new_n732), .B2(G159), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n266), .B1(new_n993), .B2(KEYINPUT51), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n201), .B2(new_n716), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n993), .A2(KEYINPUT51), .ZN(new_n996));
  AND2_X1   g0796(.A1(new_n721), .A2(G143), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n729), .A2(new_n202), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(new_n734), .B2(G50), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n999), .B(new_n775), .C1(new_n291), .C2(new_n727), .ZN(new_n1000));
  NOR4_X1   g0800(.A1(new_n995), .A2(new_n996), .A3(new_n997), .A4(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n992), .A2(new_n1001), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT110), .Z(new_n1003));
  OAI221_X1 g0803(.A(new_n985), .B1(new_n898), .B2(new_n905), .C1(new_n1003), .C2(new_n754), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n901), .ZN(new_n1005));
  AND2_X1   g0805(.A1(new_n915), .A2(new_n945), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n658), .B1(new_n915), .B2(new_n945), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1004), .B1(new_n1005), .B2(new_n915), .C1(new_n1006), .C2(new_n1007), .ZN(G390));
  AOI21_X1  g0808(.A(new_n856), .B1(new_n684), .B2(new_n764), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n400), .A2(new_n803), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n395), .A2(new_n399), .A3(new_n804), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n765), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  AND3_X1   g0812(.A1(new_n1012), .A2(new_n841), .A3(G330), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n854), .B1(new_n1009), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n841), .A2(G330), .A3(new_n764), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n855), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n762), .B1(new_n761), .B2(new_n764), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n684), .A2(new_n764), .A3(new_n856), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1014), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n465), .A2(G330), .A3(new_n841), .ZN(new_n1021));
  AND3_X1   g0821(.A1(new_n860), .A2(new_n626), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n850), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n1017), .B2(new_n855), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1026), .A2(new_n846), .A3(new_n849), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n828), .A2(new_n836), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1028), .B(new_n1025), .C1(new_n855), .C2(new_n1017), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1013), .ZN(new_n1030));
  AND3_X1   g0830(.A1(new_n1027), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1018), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1032));
  OR3_X1    g0832(.A1(new_n1024), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1024), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1033), .A2(new_n658), .A3(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n901), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n700), .B1(new_n846), .B2(new_n849), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT111), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n794), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n266), .B1(new_n721), .B2(G125), .ZN(new_n1040));
  INV_X1    g0840(.A(G128), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1040), .B1(new_n409), .B2(new_n729), .C1(new_n770), .C2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n716), .A2(new_n962), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT53), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(KEYINPUT54), .B(G143), .ZN(new_n1045));
  INV_X1    g0845(.A(G137), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1044), .B1(new_n727), .B2(new_n1045), .C1(new_n1046), .C2(new_n735), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n1042), .B(new_n1047), .C1(G50), .C2(new_n714), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n732), .A2(G132), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n260), .B1(new_n709), .B2(G283), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n726), .A2(G97), .ZN(new_n1051));
  AND3_X1   g0851(.A1(new_n1050), .A2(new_n788), .A3(new_n1051), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n718), .B1(new_n743), .B2(new_n720), .C1(new_n733), .C2(new_n520), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n998), .B(new_n1053), .C1(G107), .C2(new_n734), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n1048), .A2(new_n1049), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n689), .B1(new_n348), .B2(new_n1039), .C1(new_n1055), .C2(new_n754), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1037), .B1(new_n1038), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n1038), .B2(new_n1056), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1035), .A2(new_n1036), .A3(new_n1058), .ZN(G378));
  NAND2_X1  g0859(.A1(new_n1012), .A2(new_n841), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n847), .B2(new_n848), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n837), .B(G330), .C1(new_n1061), .C2(KEYINPUT40), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n313), .A2(new_n318), .A3(new_n326), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT114), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n307), .A2(new_n633), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  OR3_X1    g0869(.A1(new_n1066), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1069), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1062), .A2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n831), .A2(G330), .A3(new_n837), .A4(new_n1072), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n859), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1074), .A2(new_n1075), .A3(new_n859), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n901), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1072), .A2(new_n699), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n295), .B1(new_n264), .B2(G41), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n727), .A2(new_n1046), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n733), .A2(new_n1041), .B1(new_n287), .B2(new_n729), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n1084), .B(new_n1085), .C1(G125), .C2(new_n709), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1086), .B1(new_n790), .B2(new_n735), .C1(new_n716), .C2(new_n1045), .ZN(new_n1087));
  OR2_X1    g0887(.A1(new_n1087), .A2(KEYINPUT59), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n714), .A2(G159), .ZN(new_n1089));
  AOI21_X1  g0889(.A(G41), .B1(new_n721), .B2(G124), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1088), .A2(new_n257), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1091));
  AND2_X1   g0891(.A1(new_n1087), .A2(KEYINPUT59), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1083), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  OR3_X1    g0893(.A1(new_n733), .A2(KEYINPUT112), .A3(new_n493), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n961), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n714), .A2(G58), .ZN(new_n1096));
  OAI21_X1  g0896(.A(KEYINPUT112), .B1(new_n733), .B2(new_n493), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(G41), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n729), .B2(new_n201), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n720), .A2(new_n953), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n266), .B1(new_n727), .B2(new_n351), .ZN(new_n1102));
  NOR4_X1   g0902(.A1(new_n1098), .A2(new_n1100), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n1103), .B1(new_n489), .B2(new_n735), .C1(new_n520), .C2(new_n770), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(KEYINPUT113), .B(KEYINPUT58), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1104), .B(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n702), .B1(new_n1093), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n794), .A2(new_n295), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1082), .A2(new_n689), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1081), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1078), .A2(KEYINPUT115), .A3(new_n1079), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1034), .A2(new_n1022), .ZN(new_n1113));
  OR2_X1    g0913(.A1(new_n1079), .A2(KEYINPUT115), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(KEYINPUT57), .B1(new_n1034), .B2(new_n1022), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1115), .A2(KEYINPUT57), .B1(new_n1080), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1111), .B1(new_n1117), .B2(new_n659), .ZN(G375));
  NAND3_X1  g0918(.A1(new_n860), .A2(new_n626), .A3(new_n1021), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1119), .A2(new_n1014), .A3(new_n1019), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1023), .A2(new_n924), .A3(new_n1120), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n856), .A2(new_n700), .B1(G68), .B2(new_n1039), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(G283), .A2(new_n732), .B1(new_n709), .B2(G294), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n266), .B1(new_n713), .B2(new_n202), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1123), .B(new_n965), .C1(KEYINPUT116), .C2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n716), .A2(new_n489), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1124), .A2(KEYINPUT116), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n727), .A2(new_n493), .ZN(new_n1128));
  NOR4_X1   g0928(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1129), .B1(new_n520), .B2(new_n735), .C1(new_n737), .C2(new_n720), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT117), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1096), .B1(new_n409), .B2(new_n716), .C1(new_n770), .C2(new_n790), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n733), .A2(new_n1046), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n735), .A2(new_n1045), .ZN(new_n1134));
  OR4_X1    g0934(.A1(new_n266), .A2(new_n1132), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(G50), .B2(new_n776), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n1136), .B1(new_n1041), .B2(new_n720), .C1(new_n287), .C2(new_n727), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n754), .B1(new_n1131), .B2(new_n1137), .ZN(new_n1138));
  NOR3_X1   g0938(.A1(new_n1122), .A2(new_n688), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(new_n1020), .B2(new_n901), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1121), .A2(new_n1140), .ZN(G381));
  INV_X1    g0941(.A(G378), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1142), .B(new_n1111), .C1(new_n1117), .C2(new_n659), .ZN(new_n1143));
  NOR3_X1   g0943(.A1(new_n1143), .A2(G384), .A3(G381), .ZN(new_n1144));
  OR2_X1    g0944(.A1(G387), .A2(G390), .ZN(new_n1145));
  NOR3_X1   g0945(.A1(new_n1145), .A2(G396), .A3(G393), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1144), .A2(new_n1146), .ZN(G407));
  OAI211_X1 g0947(.A(G407), .B(G213), .C1(G343), .C2(new_n1143), .ZN(G409));
  NAND2_X1  g0948(.A1(new_n1115), .A2(KEYINPUT57), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1116), .A2(new_n1080), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n659), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(G378), .B1(new_n1151), .B2(new_n1110), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1113), .A2(new_n1080), .A3(new_n924), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT118), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT119), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1112), .A2(KEYINPUT119), .A3(new_n1114), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1157), .A2(new_n1158), .A3(new_n901), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1154), .A2(new_n1159), .A3(new_n1142), .A4(new_n1109), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n634), .A2(G213), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT120), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT60), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1120), .A2(new_n1163), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1119), .A2(new_n1014), .A3(KEYINPUT60), .A4(new_n1019), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1164), .A2(new_n658), .A3(new_n1023), .A4(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1166), .A2(G384), .A3(new_n1140), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(G384), .B1(new_n1166), .B2(new_n1140), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1162), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1166), .A2(new_n1140), .ZN(new_n1171));
  INV_X1    g0971(.A(G384), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1173), .A2(KEYINPUT120), .A3(new_n1167), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1170), .A2(new_n1174), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1152), .A2(new_n1160), .A3(new_n1161), .A4(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT124), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT62), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(G375), .A2(G378), .B1(G213), .B2(new_n634), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1181), .A2(new_n1160), .A3(new_n1175), .A4(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1179), .A2(new_n1180), .A3(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n634), .A2(G213), .A3(G2897), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1170), .A2(new_n1185), .A3(new_n1174), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT121), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1173), .A2(new_n1167), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1185), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1187), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1186), .A2(new_n1190), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1170), .A2(new_n1174), .A3(new_n1187), .A4(new_n1185), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n1181), .B2(new_n1160), .ZN(new_n1194));
  OAI21_X1  g0994(.A(KEYINPUT123), .B1(new_n1194), .B2(KEYINPUT61), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT123), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT61), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n1181), .A2(new_n1160), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1196), .B(new_n1197), .C1(new_n1198), .C2(new_n1193), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1184), .A2(new_n1195), .A3(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(G393), .B(new_n759), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(G387), .A2(G390), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(G387), .A2(G390), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1201), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1201), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1145), .A2(new_n1206), .A3(new_n1202), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1205), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1200), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT63), .ZN(new_n1210));
  AOI211_X1 g1010(.A(KEYINPUT61), .B(new_n1208), .C1(new_n1176), .C2(new_n1210), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1193), .B(KEYINPUT122), .Z(new_n1212));
  OAI221_X1 g1012(.A(new_n1211), .B1(new_n1210), .B2(new_n1176), .C1(new_n1212), .C2(new_n1198), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1209), .A2(new_n1213), .ZN(G405));
  NOR2_X1   g1014(.A1(new_n1208), .A2(KEYINPUT126), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1152), .A2(new_n1143), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n1188), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1152), .A2(new_n1143), .A3(new_n1175), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1218), .A2(KEYINPUT125), .A3(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT127), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT126), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n1205), .B2(new_n1207), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1188), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n1152), .B2(new_n1143), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT125), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1223), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n1220), .A2(new_n1221), .A3(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1221), .B1(new_n1220), .B2(new_n1227), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1216), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1152), .A2(new_n1143), .A3(new_n1175), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(new_n1231), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1217), .A2(new_n1226), .A3(new_n1188), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1223), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(KEYINPUT127), .B1(new_n1232), .B2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1220), .A2(new_n1221), .A3(new_n1227), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1236), .A2(new_n1215), .A3(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1230), .A2(new_n1238), .ZN(G402));
endmodule


