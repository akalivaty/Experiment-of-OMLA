//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 1 0 1 0 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:12 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050;
  INV_X1    g000(.A(KEYINPUT82), .ZN(new_n187));
  INV_X1    g001(.A(G143), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT1), .B1(new_n188), .B2(G146), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(G146), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  OAI211_X1 g006(.A(G128), .B(new_n189), .C1(new_n190), .C2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n188), .A2(G146), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n194), .B(new_n195), .C1(KEYINPUT1), .C2(new_n196), .ZN(new_n197));
  AND2_X1   g011(.A1(new_n193), .A2(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n187), .B1(new_n198), .B2(G125), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n193), .A2(new_n197), .ZN(new_n200));
  INV_X1    g014(.A(G125), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(KEYINPUT82), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT0), .ZN(new_n203));
  NOR4_X1   g017(.A1(new_n190), .A2(new_n192), .A3(new_n203), .A4(new_n196), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n206), .B1(new_n194), .B2(new_n195), .ZN(new_n207));
  AND3_X1   g021(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n208));
  AOI21_X1  g022(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AND3_X1   g024(.A1(new_n207), .A2(KEYINPUT65), .A3(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(KEYINPUT65), .B1(new_n207), .B2(new_n210), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n205), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI22_X1  g027(.A1(new_n199), .A2(new_n202), .B1(new_n213), .B2(G125), .ZN(new_n214));
  INV_X1    g028(.A(G953), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G224), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n214), .B(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G104), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT3), .B1(new_n218), .B2(G107), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n220));
  INV_X1    g034(.A(G107), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n221), .A3(G104), .ZN(new_n222));
  INV_X1    g036(.A(G101), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n218), .A2(G107), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n219), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n219), .A2(new_n222), .A3(new_n224), .ZN(new_n226));
  AOI22_X1  g040(.A1(new_n225), .A2(KEYINPUT4), .B1(new_n226), .B2(G101), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n226), .A2(KEYINPUT4), .A3(G101), .ZN(new_n228));
  INV_X1    g042(.A(G119), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G116), .ZN(new_n230));
  INV_X1    g044(.A(G116), .ZN(new_n231));
  AND3_X1   g045(.A1(new_n231), .A2(KEYINPUT68), .A3(G119), .ZN(new_n232));
  AOI21_X1  g046(.A(KEYINPUT68), .B1(new_n231), .B2(G119), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n230), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(KEYINPUT2), .A2(G113), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT67), .B1(KEYINPUT2), .B2(G113), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NOR3_X1   g051(.A1(KEYINPUT67), .A2(KEYINPUT2), .A3(G113), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n235), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n234), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(KEYINPUT2), .A2(G113), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n243), .A2(new_n236), .B1(KEYINPUT2), .B2(G113), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n231), .A2(G119), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n246), .B1(new_n229), .B2(G116), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n231), .A2(KEYINPUT68), .A3(G119), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n245), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n244), .A2(new_n249), .ZN(new_n250));
  OAI22_X1  g064(.A1(new_n227), .A2(new_n228), .B1(new_n240), .B2(new_n250), .ZN(new_n251));
  OAI211_X1 g065(.A(KEYINPUT5), .B(new_n230), .C1(new_n232), .C2(new_n233), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT79), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n253), .B1(new_n230), .B2(KEYINPUT5), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT5), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n255), .A2(new_n229), .A3(KEYINPUT79), .A4(G116), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n252), .A2(new_n257), .A3(G113), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n218), .A2(G107), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n221), .A2(G104), .ZN(new_n260));
  OAI21_X1  g074(.A(G101), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n225), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n244), .A2(new_n249), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n258), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n251), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT80), .ZN(new_n267));
  XNOR2_X1  g081(.A(G110), .B(G122), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT81), .B(KEYINPUT6), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT80), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n251), .A2(new_n271), .A3(new_n265), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n267), .A2(new_n269), .A3(new_n270), .A4(new_n272), .ZN(new_n273));
  AND3_X1   g087(.A1(new_n267), .A2(new_n269), .A3(new_n272), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n251), .A2(new_n265), .A3(new_n268), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(KEYINPUT6), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n217), .B(new_n273), .C1(new_n274), .C2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(G902), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT85), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n216), .A2(KEYINPUT7), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n280), .B1(new_n214), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT65), .ZN(new_n284));
  INV_X1    g098(.A(new_n206), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n285), .B1(new_n190), .B2(new_n192), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT64), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n287), .B1(new_n203), .B2(new_n196), .ZN(new_n288));
  NAND3_X1  g102(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n284), .B1(new_n286), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n207), .A2(new_n210), .A3(KEYINPUT65), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n204), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(KEYINPUT82), .B1(new_n200), .B2(new_n201), .ZN(new_n294));
  AOI211_X1 g108(.A(new_n187), .B(G125), .C1(new_n193), .C2(new_n197), .ZN(new_n295));
  OAI22_X1  g109(.A1(new_n293), .A2(new_n201), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n296), .A2(KEYINPUT85), .A3(new_n281), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n214), .A2(KEYINPUT86), .A3(new_n282), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT86), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n299), .B1(new_n296), .B2(new_n281), .ZN(new_n300));
  AOI22_X1  g114(.A1(new_n283), .A2(new_n297), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n252), .A2(new_n257), .A3(G113), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n225), .B(new_n261), .C1(new_n234), .C2(new_n239), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT83), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(KEYINPUT79), .B1(new_n245), .B2(new_n255), .ZN(new_n305));
  INV_X1    g119(.A(new_n256), .ZN(new_n306));
  OAI21_X1  g120(.A(G113), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AOI221_X4 g121(.A(new_n255), .B1(G116), .B2(new_n229), .C1(new_n247), .C2(new_n248), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n264), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n262), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT83), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n258), .A2(new_n263), .A3(new_n311), .A4(new_n264), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n304), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n268), .B(KEYINPUT8), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT84), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT84), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n313), .A2(new_n317), .A3(new_n314), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n301), .A2(new_n319), .A3(KEYINPUT87), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n275), .ZN(new_n321));
  AOI21_X1  g135(.A(KEYINPUT87), .B1(new_n301), .B2(new_n319), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n279), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT88), .ZN(new_n324));
  OAI21_X1  g138(.A(G210), .B1(G237), .B2(G902), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT87), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n283), .A2(new_n297), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n298), .A2(new_n300), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n313), .A2(new_n317), .A3(new_n314), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n317), .B1(new_n313), .B2(new_n314), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n327), .B1(new_n330), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(new_n275), .A3(new_n320), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT88), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n335), .A2(new_n336), .A3(new_n279), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n324), .A2(new_n326), .A3(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n335), .A2(new_n279), .A3(new_n325), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(G214), .B1(G237), .B2(G902), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT99), .ZN(new_n342));
  NAND2_X1  g156(.A1(KEYINPUT95), .A2(G122), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(KEYINPUT95), .A2(G122), .ZN(new_n345));
  OAI21_X1  g159(.A(G116), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n221), .B1(new_n346), .B2(KEYINPUT14), .ZN(new_n347));
  INV_X1    g161(.A(G122), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n348), .A2(G116), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT95), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n348), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n231), .B1(new_n351), .B2(new_n343), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n347), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n349), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n346), .B(new_n354), .C1(KEYINPUT14), .C2(new_n221), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n188), .A2(G128), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n196), .A2(G143), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n358), .A2(KEYINPUT97), .ZN(new_n359));
  XNOR2_X1  g173(.A(G128), .B(G143), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT97), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G134), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n359), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n358), .A2(KEYINPUT97), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n360), .A2(new_n361), .ZN(new_n366));
  AOI21_X1  g180(.A(G134), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n353), .B(new_n355), .C1(new_n364), .C2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n360), .A2(KEYINPUT13), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n369), .B(G134), .C1(KEYINPUT13), .C2(new_n356), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT98), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n367), .A2(new_n371), .ZN(new_n372));
  AOI211_X1 g186(.A(KEYINPUT98), .B(G134), .C1(new_n365), .C2(new_n366), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n370), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT96), .B1(new_n352), .B2(new_n349), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT96), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n346), .A2(new_n376), .A3(new_n354), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n221), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n375), .A2(G107), .A3(new_n377), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n368), .B1(new_n374), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(KEYINPUT9), .B(G234), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  XOR2_X1   g198(.A(KEYINPUT72), .B(G217), .Z(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n385), .A3(new_n215), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n386), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n368), .B(new_n388), .C1(new_n374), .C2(new_n381), .ZN(new_n389));
  AOI21_X1  g203(.A(G902), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(G478), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n391), .A2(KEYINPUT15), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  AOI211_X1 g208(.A(G902), .B(new_n392), .C1(new_n387), .C2(new_n389), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n342), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n363), .B1(new_n359), .B2(new_n362), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(KEYINPUT98), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n367), .A2(new_n371), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n400), .A2(new_n370), .A3(new_n379), .A4(new_n380), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n388), .B1(new_n401), .B2(new_n368), .ZN(new_n402));
  INV_X1    g216(.A(new_n389), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n278), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n392), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n390), .A2(new_n393), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(KEYINPUT99), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n396), .A2(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(G125), .B(G140), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT16), .ZN(new_n410));
  INV_X1    g224(.A(G140), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G125), .ZN(new_n412));
  OR2_X1    g226(.A1(new_n412), .A2(KEYINPUT16), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n410), .A2(G146), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(G146), .B1(new_n410), .B2(new_n413), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G237), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(new_n215), .A3(G214), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n419), .B1(KEYINPUT89), .B2(new_n188), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT89), .B(G143), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n420), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(G131), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT17), .ZN(new_n424));
  NOR2_X1   g238(.A1(G237), .A2(G953), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n188), .A2(KEYINPUT89), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n188), .A2(KEYINPUT89), .ZN(new_n427));
  OAI211_X1 g241(.A(G214), .B(new_n425), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(G131), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n428), .A2(new_n429), .A3(new_n420), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n423), .A2(new_n424), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n422), .A2(KEYINPUT17), .A3(G131), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT94), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n429), .B1(new_n428), .B2(new_n420), .ZN(new_n435));
  AOI21_X1  g249(.A(KEYINPUT94), .B1(new_n435), .B2(KEYINPUT17), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n417), .B(new_n431), .C1(new_n434), .C2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n201), .A2(G140), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n412), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G146), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n409), .A2(new_n191), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT91), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT18), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n445), .A2(new_n429), .A3(KEYINPUT90), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n422), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n446), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n428), .A2(new_n448), .A3(new_n420), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n440), .A2(new_n441), .A3(KEYINPUT91), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n444), .A2(new_n447), .A3(new_n449), .A4(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(G113), .B(G122), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(new_n218), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(KEYINPUT93), .ZN(new_n454));
  AND3_X1   g268(.A1(new_n437), .A2(new_n451), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n453), .B1(new_n437), .B2(new_n451), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n278), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G475), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT20), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n437), .A2(new_n451), .A3(new_n454), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT19), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n409), .B1(KEYINPUT92), .B2(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n462), .B(new_n191), .C1(new_n409), .C2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n430), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n464), .B1(new_n465), .B2(new_n435), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n414), .A2(KEYINPUT74), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT74), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n410), .A2(new_n468), .A3(new_n413), .A4(G146), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n451), .B1(new_n466), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n453), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n460), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(G475), .A2(G902), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n459), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n475), .ZN(new_n477));
  AOI211_X1 g291(.A(KEYINPUT20), .B(new_n477), .C1(new_n460), .C2(new_n473), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n458), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  OR2_X1    g293(.A1(KEYINPUT100), .A2(G952), .ZN(new_n480));
  NAND2_X1  g294(.A1(KEYINPUT100), .A2(G952), .ZN(new_n481));
  AOI21_X1  g295(.A(G953), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(G234), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n482), .B1(new_n483), .B2(new_n418), .ZN(new_n484));
  OAI211_X1 g298(.A(G902), .B(G953), .C1(new_n483), .C2(new_n418), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n485), .B(KEYINPUT101), .ZN(new_n486));
  XNOR2_X1  g300(.A(KEYINPUT21), .B(G898), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n484), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NOR3_X1   g304(.A1(new_n408), .A2(new_n479), .A3(new_n490), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n340), .A2(new_n341), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(G469), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n293), .B1(new_n227), .B2(new_n228), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT11), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n495), .B1(new_n363), .B2(G137), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n363), .A2(G137), .ZN(new_n497));
  INV_X1    g311(.A(G137), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(KEYINPUT11), .A3(G134), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n496), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(G131), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n496), .A2(new_n499), .A3(new_n429), .A4(new_n497), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n501), .A2(KEYINPUT69), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(KEYINPUT69), .B1(new_n501), .B2(new_n502), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n193), .A2(new_n225), .A3(new_n261), .A4(new_n197), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT10), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n198), .A2(new_n263), .A3(KEYINPUT10), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n494), .A2(new_n505), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  XNOR2_X1  g324(.A(G110), .B(G140), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n215), .A2(G227), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n511), .B(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n501), .A2(new_n502), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT69), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n501), .A2(KEYINPUT69), .A3(new_n502), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n200), .A2(new_n262), .ZN(new_n520));
  AOI22_X1  g334(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n506), .ZN(new_n521));
  OAI21_X1  g335(.A(KEYINPUT78), .B1(new_n521), .B2(KEYINPUT12), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT78), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT12), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n520), .A2(new_n506), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n523), .B(new_n524), .C1(new_n526), .C2(new_n505), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n525), .A2(KEYINPUT12), .A3(new_n516), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n515), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n494), .A2(new_n508), .A3(new_n509), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n518), .A2(new_n519), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n514), .B1(new_n533), .B2(new_n510), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n493), .B(new_n278), .C1(new_n530), .C2(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n493), .A2(new_n278), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n510), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n538), .B1(new_n528), .B2(new_n529), .ZN(new_n539));
  INV_X1    g353(.A(new_n533), .ZN(new_n540));
  OAI22_X1  g354(.A1(new_n539), .A2(new_n514), .B1(new_n540), .B2(new_n515), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n535), .B(new_n537), .C1(new_n541), .C2(new_n493), .ZN(new_n542));
  OAI21_X1  g356(.A(G221), .B1(new_n383), .B2(G902), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT25), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n196), .A2(G119), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT23), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n196), .A2(KEYINPUT23), .A3(G119), .ZN(new_n549));
  INV_X1    g363(.A(G110), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n229), .A2(G128), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n548), .A2(new_n549), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n546), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT24), .B(G110), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI22_X1  g369(.A1(new_n552), .A2(new_n555), .B1(new_n191), .B2(new_n409), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n467), .A2(new_n556), .A3(new_n469), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT75), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n548), .A2(new_n549), .A3(new_n551), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(G110), .ZN(new_n560));
  OAI221_X1 g374(.A(new_n560), .B1(new_n553), .B2(new_n554), .C1(new_n415), .C2(new_n416), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT75), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n467), .A2(new_n556), .A3(new_n562), .A4(new_n469), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n558), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n215), .A2(G221), .A3(G234), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(KEYINPUT76), .ZN(new_n566));
  XNOR2_X1  g380(.A(KEYINPUT22), .B(G137), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n566), .B(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n558), .A2(new_n561), .A3(new_n563), .A4(new_n568), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n545), .B1(new_n572), .B2(new_n278), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n570), .A2(new_n545), .A3(new_n278), .A4(new_n571), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n385), .B1(new_n483), .B2(G902), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(KEYINPUT73), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  OR2_X1    g391(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n576), .A2(G902), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n572), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n578), .A2(KEYINPUT77), .A3(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n580), .B1(new_n573), .B2(new_n577), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT77), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n240), .A2(new_n250), .ZN(new_n586));
  INV_X1    g400(.A(new_n497), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n363), .A2(G137), .ZN(new_n588));
  OAI21_X1  g402(.A(G131), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AND4_X1   g403(.A1(new_n197), .A2(new_n589), .A3(new_n193), .A4(new_n502), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n586), .B(new_n591), .C1(new_n505), .C2(new_n213), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT70), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n532), .A2(new_n293), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n595), .A2(KEYINPUT70), .A3(new_n586), .A4(new_n591), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  AOI22_X1  g411(.A1(new_n213), .A2(KEYINPUT66), .B1(new_n502), .B2(new_n501), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT66), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n205), .B(new_n599), .C1(new_n211), .C2(new_n212), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n590), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n601), .A2(new_n586), .ZN(new_n602));
  OAI21_X1  g416(.A(KEYINPUT28), .B1(new_n597), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT28), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n592), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n425), .A2(G210), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(KEYINPUT27), .ZN(new_n608));
  XNOR2_X1  g422(.A(KEYINPUT26), .B(G101), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n213), .A2(KEYINPUT66), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n612), .A2(new_n600), .A3(new_n516), .ZN(new_n613));
  AOI21_X1  g427(.A(KEYINPUT30), .B1(new_n613), .B2(new_n591), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT30), .ZN(new_n615));
  AOI211_X1 g429(.A(new_n615), .B(new_n590), .C1(new_n532), .C2(new_n293), .ZN(new_n616));
  NOR3_X1   g430(.A1(new_n614), .A2(new_n586), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n594), .A2(new_n596), .A3(new_n610), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT31), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n606), .A2(new_n611), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT71), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n622), .B1(new_n617), .B2(new_n618), .ZN(new_n623));
  INV_X1    g437(.A(new_n597), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n595), .A2(KEYINPUT30), .A3(new_n591), .ZN(new_n625));
  INV_X1    g439(.A(new_n586), .ZN(new_n626));
  OAI211_X1 g440(.A(new_n625), .B(new_n626), .C1(new_n601), .C2(KEYINPUT30), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n624), .A2(new_n627), .A3(KEYINPUT71), .A4(new_n610), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n623), .A2(new_n628), .A3(KEYINPUT31), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n621), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(G472), .A2(G902), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT32), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n605), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n591), .B1(new_n505), .B2(new_n213), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n626), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n594), .A2(new_n596), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n635), .B1(new_n638), .B2(KEYINPUT28), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT29), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n611), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(G902), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n516), .B1(new_n293), .B2(new_n599), .ZN(new_n643));
  INV_X1    g457(.A(new_n600), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n591), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n616), .B1(new_n615), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n597), .B1(new_n646), .B2(new_n626), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n640), .B1(new_n647), .B2(new_n610), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n594), .B(new_n596), .C1(new_n586), .C2(new_n601), .ZN(new_n649));
  AOI211_X1 g463(.A(new_n611), .B(new_n635), .C1(new_n649), .C2(KEYINPUT28), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n642), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n630), .A2(new_n634), .B1(new_n651), .B2(G472), .ZN(new_n652));
  AND3_X1   g466(.A1(new_n623), .A2(new_n628), .A3(KEYINPUT31), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n635), .B1(new_n649), .B2(KEYINPUT28), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n624), .A2(new_n627), .A3(new_n610), .ZN(new_n655));
  OAI22_X1  g469(.A1(new_n654), .A2(new_n610), .B1(new_n655), .B2(KEYINPUT31), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n631), .B1(new_n653), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n633), .ZN(new_n658));
  AOI211_X1 g472(.A(new_n544), .B(new_n585), .C1(new_n652), .C2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n492), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT102), .B(G101), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G3));
  OAI21_X1  g476(.A(new_n278), .B1(new_n653), .B2(new_n656), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(G472), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n657), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n542), .A2(new_n543), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n666), .A2(new_n584), .A3(new_n581), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n335), .A2(new_n279), .A3(new_n325), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n325), .B1(new_n335), .B2(new_n279), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n341), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n671), .A2(new_n490), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n278), .A2(G478), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n387), .A2(new_n389), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(KEYINPUT103), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT33), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n674), .A2(KEYINPUT103), .A3(KEYINPUT33), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n673), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n390), .A2(G478), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n479), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n668), .A2(new_n672), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n683), .B(KEYINPUT104), .Z(new_n684));
  XOR2_X1   g498(.A(KEYINPUT34), .B(G104), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G6));
  NOR3_X1   g500(.A1(new_n476), .A2(new_n478), .A3(KEYINPUT105), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n474), .A2(new_n475), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n688), .A2(KEYINPUT105), .A3(KEYINPUT20), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n458), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n408), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n668), .A2(new_n672), .A3(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(KEYINPUT35), .B(G107), .Z(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G9));
  NOR2_X1   g511(.A1(new_n569), .A2(KEYINPUT36), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n564), .B(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n579), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n700), .B1(new_n573), .B2(new_n577), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n542), .A2(new_n543), .A3(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n665), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n492), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g518(.A(KEYINPUT37), .B(G110), .Z(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G12));
  NAND2_X1  g520(.A1(new_n651), .A2(G472), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n634), .B1(new_n653), .B2(new_n656), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n632), .B1(new_n621), .B2(new_n629), .ZN(new_n709));
  OAI211_X1 g523(.A(new_n707), .B(new_n708), .C1(new_n709), .C2(KEYINPUT32), .ZN(new_n710));
  INV_X1    g524(.A(new_n341), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n323), .A2(new_n326), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n711), .B1(new_n712), .B2(new_n339), .ZN(new_n713));
  XOR2_X1   g527(.A(new_n484), .B(KEYINPUT106), .Z(new_n714));
  OAI21_X1  g528(.A(new_n714), .B1(G900), .B2(new_n486), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n691), .A2(new_n408), .A3(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(new_n702), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n710), .A2(new_n713), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G128), .ZN(G30));
  XNOR2_X1  g533(.A(new_n715), .B(KEYINPUT39), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n666), .A2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n666), .A2(KEYINPUT108), .A3(new_n720), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT40), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n723), .A2(KEYINPUT40), .A3(new_n724), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n340), .B(KEYINPUT38), .ZN(new_n730));
  INV_X1    g544(.A(G472), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n638), .A2(new_n611), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(KEYINPUT107), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT107), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n638), .A2(new_n734), .A3(new_n611), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n623), .A2(new_n733), .A3(new_n628), .A4(new_n735), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n731), .B1(new_n736), .B2(new_n278), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n737), .B1(new_n630), .B2(new_n634), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n658), .ZN(new_n739));
  INV_X1    g553(.A(new_n701), .ZN(new_n740));
  OR2_X1    g554(.A1(new_n476), .A2(new_n478), .ZN(new_n741));
  AOI22_X1  g555(.A1(new_n396), .A2(new_n407), .B1(new_n741), .B2(new_n458), .ZN(new_n742));
  AND4_X1   g556(.A1(new_n341), .A2(new_n739), .A3(new_n740), .A4(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n729), .A2(new_n730), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G143), .ZN(G45));
  OAI211_X1 g559(.A(new_n479), .B(new_n715), .C1(new_n679), .C2(new_n680), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n702), .A2(new_n746), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n710), .A2(new_n713), .A3(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(new_n191), .ZN(G48));
  NOR2_X1   g563(.A1(new_n530), .A2(new_n534), .ZN(new_n750));
  OAI21_X1  g564(.A(G469), .B1(new_n750), .B2(G902), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n751), .A2(new_n543), .A3(new_n535), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(KEYINPUT109), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT109), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n751), .A2(new_n754), .A3(new_n535), .A4(new_n543), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT110), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n753), .A2(KEYINPUT110), .A3(new_n755), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n585), .B1(new_n652), .B2(new_n658), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n760), .A2(new_n672), .A3(new_n761), .A4(new_n682), .ZN(new_n762));
  XNOR2_X1  g576(.A(KEYINPUT41), .B(G113), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n762), .B(new_n763), .ZN(G15));
  NAND4_X1  g578(.A1(new_n760), .A2(new_n672), .A3(new_n761), .A4(new_n694), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G116), .ZN(G18));
  NOR2_X1   g580(.A1(new_n671), .A2(new_n756), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n767), .A2(new_n491), .A3(new_n710), .A4(new_n701), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G119), .ZN(G21));
  AOI21_X1  g583(.A(new_n490), .B1(new_n758), .B2(new_n759), .ZN(new_n770));
  INV_X1    g584(.A(new_n582), .ZN(new_n771));
  OAI22_X1  g585(.A1(new_n655), .A2(KEYINPUT31), .B1(new_n639), .B2(new_n610), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n631), .B1(new_n653), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(G902), .B1(new_n621), .B2(new_n629), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n771), .B(new_n773), .C1(new_n774), .C2(new_n731), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT111), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT111), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n664), .A2(new_n777), .A3(new_n771), .A4(new_n773), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n341), .B(new_n742), .C1(new_n669), .C2(new_n670), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT112), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n712), .A2(new_n339), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n783), .A2(KEYINPUT112), .A3(new_n341), .A4(new_n742), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n770), .A2(new_n779), .A3(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G122), .ZN(G24));
  AOI21_X1  g601(.A(new_n731), .B1(new_n630), .B2(new_n278), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n639), .A2(new_n610), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n617), .A2(KEYINPUT31), .A3(new_n618), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n632), .B1(new_n791), .B2(new_n629), .ZN(new_n792));
  NOR4_X1   g606(.A1(new_n788), .A2(new_n746), .A3(new_n792), .A4(new_n740), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n767), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G125), .ZN(G27));
  INV_X1    g609(.A(KEYINPUT42), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n338), .A2(new_n341), .A3(new_n339), .A4(new_n666), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n746), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n761), .A3(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT113), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n796), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n761), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n803), .A2(new_n797), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT113), .B1(new_n804), .B2(new_n799), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n709), .A2(KEYINPUT32), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(KEYINPUT114), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT114), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n658), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n807), .A2(new_n809), .A3(new_n652), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n771), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n798), .A2(KEYINPUT42), .A3(new_n799), .ZN(new_n812));
  OAI22_X1  g626(.A1(new_n802), .A2(new_n805), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G131), .ZN(G33));
  NAND4_X1  g628(.A1(new_n798), .A2(new_n761), .A3(new_n694), .A4(new_n715), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G134), .ZN(G36));
  INV_X1    g630(.A(KEYINPUT45), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n541), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(KEYINPUT115), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n493), .B1(new_n541), .B2(new_n817), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n536), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n535), .B1(new_n821), .B2(KEYINPUT46), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT46), .ZN(new_n823));
  AOI211_X1 g637(.A(new_n823), .B(new_n536), .C1(new_n819), .C2(new_n820), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n543), .B(new_n720), .C1(new_n822), .C2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n479), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT43), .B1(new_n826), .B2(KEYINPUT116), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n826), .B1(new_n679), .B2(new_n680), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  OAI221_X1 g643(.A(new_n826), .B1(KEYINPUT116), .B2(KEYINPUT43), .C1(new_n679), .C2(new_n680), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n740), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(KEYINPUT44), .B1(new_n831), .B2(new_n665), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n831), .A2(KEYINPUT44), .A3(new_n665), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n338), .A2(new_n341), .A3(new_n339), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n825), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(new_n498), .ZN(G39));
  AOI211_X1 g651(.A(new_n746), .B(new_n710), .C1(new_n584), .C2(new_n581), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(new_n834), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n543), .B1(new_n822), .B2(new_n824), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT47), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI211_X1 g656(.A(KEYINPUT47), .B(new_n543), .C1(new_n822), .C2(new_n824), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n839), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(new_n411), .ZN(G42));
  NOR3_X1   g659(.A1(new_n730), .A2(new_n341), .A3(new_n756), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n714), .B1(new_n829), .B2(new_n830), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n779), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT121), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n851), .A2(KEYINPUT50), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n851), .A2(KEYINPUT50), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n850), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n846), .A2(new_n849), .A3(new_n852), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n751), .A2(new_n535), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n842), .B(new_n843), .C1(new_n543), .C2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n859), .A2(new_n834), .A3(new_n849), .ZN(new_n860));
  INV_X1    g674(.A(new_n834), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n861), .A2(new_n756), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n739), .A2(new_n484), .A3(new_n585), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n679), .A2(new_n479), .A3(new_n680), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT122), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n865), .A2(new_n866), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n788), .A2(new_n740), .A3(new_n792), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n862), .A2(new_n847), .ZN(new_n870));
  AOI22_X1  g684(.A1(new_n867), .A2(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n857), .A2(new_n860), .A3(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT51), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n849), .A2(new_n767), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n862), .A2(new_n682), .A3(new_n863), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n875), .A2(new_n876), .A3(new_n482), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT48), .ZN(new_n879));
  INV_X1    g693(.A(new_n811), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n870), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n879), .B1(new_n870), .B2(new_n880), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n878), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT123), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n857), .A2(KEYINPUT51), .A3(new_n860), .A4(new_n871), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n874), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n715), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n544), .A2(new_n701), .A3(new_n887), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n736), .A2(new_n278), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n708), .B1(new_n889), .B2(new_n731), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n888), .B1(new_n890), .B2(new_n806), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n891), .B1(new_n782), .B2(new_n784), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n753), .A2(new_n755), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n713), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n664), .A2(new_n799), .A3(new_n701), .A4(new_n773), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n718), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NOR4_X1   g710(.A1(new_n892), .A2(new_n896), .A3(KEYINPUT52), .A4(new_n748), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT52), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n666), .A2(new_n740), .A3(new_n715), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n658), .B2(new_n738), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n671), .B1(new_n658), .B2(new_n652), .ZN(new_n901));
  AOI22_X1  g715(.A1(new_n785), .A2(new_n900), .B1(new_n901), .B2(new_n747), .ZN(new_n902));
  INV_X1    g716(.A(new_n896), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n898), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n897), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n492), .B1(new_n659), .B2(new_n703), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n405), .A2(new_n406), .A3(new_n715), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n687), .A2(new_n907), .A3(new_n690), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n908), .A2(new_n543), .A3(new_n542), .A4(new_n701), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n909), .B1(new_n658), .B2(new_n652), .ZN(new_n910));
  AOI22_X1  g724(.A1(new_n798), .A2(new_n793), .B1(new_n834), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n394), .A2(new_n395), .ZN(new_n912));
  OR3_X1    g726(.A1(new_n479), .A2(new_n912), .A3(KEYINPUT119), .ZN(new_n913));
  OAI21_X1  g727(.A(KEYINPUT119), .B1(new_n479), .B2(new_n912), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n913), .A2(new_n681), .A3(new_n914), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n915), .A2(new_n489), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n668), .A2(new_n916), .A3(new_n341), .A4(new_n340), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n906), .A2(new_n911), .A3(new_n815), .A4(new_n917), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n786), .A2(new_n762), .A3(new_n765), .A4(new_n768), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n905), .A2(new_n920), .A3(new_n813), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT53), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(KEYINPUT120), .B1(new_n897), .B2(new_n904), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n785), .A2(new_n900), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n901), .A2(new_n747), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n925), .A2(new_n718), .A3(new_n926), .A4(new_n794), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(KEYINPUT52), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT120), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n902), .A2(new_n903), .A3(new_n898), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n924), .A2(new_n931), .A3(new_n813), .A4(new_n920), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n923), .B1(new_n932), .B2(new_n922), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(KEYINPUT54), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n932), .A2(new_n922), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT54), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n905), .A2(new_n920), .A3(KEYINPUT53), .A4(new_n813), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n934), .A2(new_n938), .ZN(new_n939));
  OAI22_X1  g753(.A1(new_n886), .A2(new_n939), .B1(G952), .B2(G953), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n858), .A2(KEYINPUT49), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT118), .Z(new_n942));
  NAND3_X1  g756(.A1(new_n771), .A2(new_n341), .A3(new_n543), .ZN(new_n943));
  OR3_X1    g757(.A1(new_n943), .A2(new_n828), .A3(KEYINPUT117), .ZN(new_n944));
  OAI21_X1  g758(.A(KEYINPUT117), .B1(new_n943), .B2(new_n828), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n858), .A2(KEYINPUT49), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n942), .A2(new_n944), .A3(new_n945), .A4(new_n946), .ZN(new_n947));
  OR3_X1    g761(.A1(new_n947), .A2(new_n730), .A3(new_n739), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n940), .A2(new_n948), .ZN(G75));
  NOR2_X1   g763(.A1(new_n215), .A2(G952), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n937), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n952), .B1(new_n922), .B2(new_n932), .ZN(new_n953));
  NAND2_X1  g767(.A1(G210), .A2(G902), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n273), .B1(new_n274), .B2(new_n276), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(new_n217), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT55), .Z(new_n958));
  OR2_X1    g772(.A1(new_n958), .A2(KEYINPUT56), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n951), .B1(new_n955), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(KEYINPUT124), .B1(new_n953), .B2(new_n954), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT56), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n935), .A2(new_n937), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT124), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n963), .A2(new_n964), .A3(G210), .A4(G902), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n961), .A2(new_n962), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n960), .B1(new_n966), .B2(new_n958), .ZN(G51));
  XNOR2_X1  g781(.A(new_n536), .B(KEYINPUT57), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n936), .B1(new_n935), .B2(new_n937), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n968), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n750), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n278), .B1(new_n935), .B2(new_n937), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n974), .A2(new_n819), .A3(new_n820), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n950), .B1(new_n973), .B2(new_n975), .ZN(G54));
  NAND2_X1  g790(.A1(KEYINPUT58), .A2(G475), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n974), .A2(new_n474), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n474), .B1(new_n974), .B2(new_n978), .ZN(new_n980));
  NOR3_X1   g794(.A1(new_n979), .A2(new_n980), .A3(new_n950), .ZN(G60));
  NAND2_X1  g795(.A1(new_n677), .A2(new_n678), .ZN(new_n982));
  NAND2_X1  g796(.A1(G478), .A2(G902), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT59), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n982), .B(new_n984), .C1(new_n969), .C2(new_n970), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n951), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n982), .B1(new_n939), .B2(new_n984), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n986), .A2(new_n987), .ZN(G63));
  INV_X1    g802(.A(KEYINPUT61), .ZN(new_n989));
  XOR2_X1   g803(.A(KEYINPUT125), .B(KEYINPUT60), .Z(new_n990));
  NAND2_X1  g804(.A1(G217), .A2(G902), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n990), .B(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n993), .B1(new_n935), .B2(new_n937), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n699), .ZN(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n951), .B1(new_n994), .B2(new_n572), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n989), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(new_n572), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n999), .B1(new_n953), .B2(new_n993), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n1000), .A2(new_n995), .A3(KEYINPUT61), .A4(new_n951), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n998), .A2(new_n1001), .ZN(G66));
  AOI21_X1  g816(.A(new_n215), .B1(new_n488), .B2(G224), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n906), .A2(new_n917), .ZN(new_n1004));
  OR2_X1    g818(.A1(new_n919), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1003), .B1(new_n1005), .B2(new_n215), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n956), .B1(G898), .B2(new_n215), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1006), .B(new_n1007), .Z(G69));
  AOI21_X1  g822(.A(new_n215), .B1(G227), .B2(G900), .ZN(new_n1009));
  INV_X1    g823(.A(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n646), .B(KEYINPUT126), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n462), .B1(new_n409), .B2(new_n463), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1011), .B(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1014), .B1(G900), .B2(G953), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n844), .A2(new_n836), .ZN(new_n1016));
  INV_X1    g830(.A(new_n785), .ZN(new_n1017));
  NOR3_X1   g831(.A1(new_n825), .A2(new_n811), .A3(new_n1017), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n903), .A2(new_n815), .A3(new_n926), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n1016), .A2(new_n813), .A3(new_n1020), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1015), .B1(new_n1021), .B2(G953), .ZN(new_n1022));
  INV_X1    g836(.A(new_n1022), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n744), .A2(new_n926), .A3(new_n903), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1024), .A2(KEYINPUT62), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n861), .A2(new_n725), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n1026), .A2(new_n761), .A3(new_n915), .ZN(new_n1027));
  INV_X1    g841(.A(KEYINPUT62), .ZN(new_n1028));
  NAND4_X1  g842(.A1(new_n744), .A2(new_n1028), .A3(new_n926), .A4(new_n903), .ZN(new_n1029));
  NAND4_X1  g843(.A1(new_n1016), .A2(new_n1025), .A3(new_n1027), .A4(new_n1029), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n1013), .B1(new_n1030), .B2(new_n215), .ZN(new_n1031));
  NOR3_X1   g845(.A1(new_n1023), .A2(new_n1031), .A3(KEYINPUT127), .ZN(new_n1032));
  INV_X1    g846(.A(KEYINPUT127), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1030), .A2(new_n215), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1034), .A2(new_n1014), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1033), .B1(new_n1035), .B2(new_n1022), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1010), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g851(.A(KEYINPUT127), .B1(new_n1023), .B2(new_n1031), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n1035), .A2(new_n1033), .A3(new_n1022), .ZN(new_n1039));
  NAND3_X1  g853(.A1(new_n1038), .A2(new_n1039), .A3(new_n1009), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1037), .A2(new_n1040), .ZN(G72));
  NAND2_X1  g855(.A1(G472), .A2(G902), .ZN(new_n1042));
  XOR2_X1   g856(.A(new_n1042), .B(KEYINPUT63), .Z(new_n1043));
  OAI21_X1  g857(.A(new_n1043), .B1(new_n1030), .B2(new_n1005), .ZN(new_n1044));
  OAI211_X1 g858(.A(new_n1044), .B(new_n610), .C1(new_n617), .C2(new_n597), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n623), .A2(new_n628), .ZN(new_n1046));
  NOR2_X1   g860(.A1(new_n647), .A2(new_n610), .ZN(new_n1047));
  OAI211_X1 g861(.A(new_n933), .B(new_n1043), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g862(.A(new_n1043), .B1(new_n1021), .B2(new_n1005), .ZN(new_n1049));
  NAND3_X1  g863(.A1(new_n1049), .A2(new_n611), .A3(new_n647), .ZN(new_n1050));
  AND4_X1   g864(.A1(new_n951), .A2(new_n1045), .A3(new_n1048), .A4(new_n1050), .ZN(G57));
endmodule


