

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736;

  NOR2_X1 U371 ( .A1(n661), .A2(n662), .ZN(n536) );
  NOR2_X1 U372 ( .A1(n653), .A2(n350), .ZN(n587) );
  XNOR2_X1 U373 ( .A(G902), .B(KEYINPUT15), .ZN(n449) );
  XNOR2_X1 U374 ( .A(n720), .B(n417), .ZN(n471) );
  XNOR2_X1 U375 ( .A(n565), .B(KEYINPUT22), .ZN(n570) );
  INV_X1 U376 ( .A(G953), .ZN(n724) );
  XNOR2_X1 U377 ( .A(n587), .B(KEYINPUT31), .ZN(n633) );
  NOR2_X2 U378 ( .A1(n380), .A2(n615), .ZN(n591) );
  XNOR2_X2 U379 ( .A(n405), .B(KEYINPUT19), .ZN(n557) );
  XOR2_X2 U380 ( .A(KEYINPUT38), .B(n363), .Z(n658) );
  XNOR2_X2 U381 ( .A(n527), .B(n526), .ZN(n642) );
  NOR2_X1 U382 ( .A1(n642), .A2(n641), .ZN(n584) );
  INV_X1 U383 ( .A(KEYINPUT16), .ZN(n409) );
  INV_X1 U384 ( .A(KEYINPUT4), .ZN(n371) );
  XNOR2_X1 U385 ( .A(n382), .B(n381), .ZN(n421) );
  XNOR2_X1 U386 ( .A(n652), .B(n522), .ZN(n579) );
  XNOR2_X1 U387 ( .A(n488), .B(n379), .ZN(n541) );
  OR2_X2 U388 ( .A1(n373), .A2(n372), .ZN(n652) );
  XNOR2_X1 U389 ( .A(n507), .B(n408), .ZN(n705) );
  XNOR2_X1 U390 ( .A(n485), .B(n409), .ZN(n408) );
  XNOR2_X1 U391 ( .A(n704), .B(n411), .ZN(n484) );
  NOR2_X1 U392 ( .A1(n423), .A2(G953), .ZN(n422) );
  XNOR2_X1 U393 ( .A(n371), .B(KEYINPUT64), .ZN(n480) );
  XNOR2_X1 U394 ( .A(n481), .B(G134), .ZN(n493) );
  XOR2_X1 U395 ( .A(G131), .B(G140), .Z(n504) );
  BUF_X1 U396 ( .A(n734), .Z(n349) );
  BUF_X1 U397 ( .A(n586), .Z(n350) );
  XNOR2_X1 U398 ( .A(n577), .B(n578), .ZN(n734) );
  XNOR2_X1 U399 ( .A(n560), .B(n559), .ZN(n586) );
  NAND2_X1 U400 ( .A1(n421), .A2(n419), .ZN(n723) );
  NAND2_X1 U401 ( .A1(n399), .A2(n400), .ZN(n382) );
  NOR2_X1 U402 ( .A1(n418), .A2(n732), .ZN(n393) );
  NOR2_X1 U403 ( .A1(n642), .A2(n641), .ZN(n351) );
  XOR2_X1 U404 ( .A(n439), .B(KEYINPUT62), .Z(n605) );
  NAND2_X1 U405 ( .A1(n407), .A2(n425), .ZN(n352) );
  NAND2_X1 U406 ( .A1(n407), .A2(n425), .ZN(n594) );
  XNOR2_X1 U407 ( .A(n471), .B(n414), .ZN(n439) );
  INV_X1 U408 ( .A(G146), .ZN(n417) );
  AND2_X1 U409 ( .A1(n638), .A2(n364), .ZN(n400) );
  NOR2_X1 U410 ( .A1(n401), .A2(n365), .ZN(n364) );
  XNOR2_X1 U411 ( .A(n370), .B(n493), .ZN(n720) );
  XNOR2_X1 U412 ( .A(n480), .B(G137), .ZN(n370) );
  INV_X1 U413 ( .A(n723), .ZN(n396) );
  NOR2_X1 U414 ( .A1(G902), .A2(G237), .ZN(n440) );
  INV_X1 U415 ( .A(n579), .ZN(n571) );
  NAND2_X1 U416 ( .A1(n374), .A2(n377), .ZN(n373) );
  NAND2_X1 U417 ( .A1(n378), .A2(G902), .ZN(n377) );
  NOR2_X1 U418 ( .A1(G953), .A2(G237), .ZN(n500) );
  INV_X1 U419 ( .A(KEYINPUT79), .ZN(n590) );
  XNOR2_X1 U420 ( .A(KEYINPUT65), .B(n595), .ZN(n596) );
  XNOR2_X1 U421 ( .A(n430), .B(KEYINPUT86), .ZN(n379) );
  NAND2_X1 U422 ( .A1(n585), .A2(n659), .ZN(n441) );
  NAND2_X1 U423 ( .A1(n439), .A2(n378), .ZN(n374) );
  INV_X1 U424 ( .A(KEYINPUT95), .ZN(n434) );
  NOR2_X1 U425 ( .A1(n639), .A2(n420), .ZN(n419) );
  INV_X1 U426 ( .A(n640), .ZN(n420) );
  XNOR2_X1 U427 ( .A(n484), .B(n384), .ZN(n472) );
  XNOR2_X1 U428 ( .A(n469), .B(n468), .ZN(n470) );
  NAND2_X1 U429 ( .A1(n369), .A2(n353), .ZN(n548) );
  INV_X1 U430 ( .A(n524), .ZN(n368) );
  XNOR2_X1 U431 ( .A(n521), .B(n520), .ZN(n522) );
  INV_X1 U432 ( .A(KEYINPUT6), .ZN(n520) );
  XNOR2_X1 U433 ( .A(n719), .B(n402), .ZN(n461) );
  XNOR2_X1 U434 ( .A(n459), .B(n357), .ZN(n460) );
  XNOR2_X1 U435 ( .A(n403), .B(n455), .ZN(n402) );
  NAND2_X1 U436 ( .A1(n530), .A2(n529), .ZN(n365) );
  INV_X1 U437 ( .A(KEYINPUT80), .ZN(n406) );
  INV_X1 U438 ( .A(G224), .ZN(n423) );
  XNOR2_X1 U439 ( .A(n453), .B(n383), .ZN(n645) );
  INV_X1 U440 ( .A(KEYINPUT21), .ZN(n383) );
  XNOR2_X1 U441 ( .A(n645), .B(KEYINPUT94), .ZN(n561) );
  INV_X1 U442 ( .A(KEYINPUT48), .ZN(n381) );
  XNOR2_X1 U443 ( .A(G146), .B(G125), .ZN(n479) );
  XOR2_X1 U444 ( .A(G143), .B(KEYINPUT11), .Z(n502) );
  INV_X1 U445 ( .A(G104), .ZN(n468) );
  INV_X1 U446 ( .A(KEYINPUT69), .ZN(n411) );
  NAND2_X1 U447 ( .A1(G234), .A2(G237), .ZN(n443) );
  INV_X1 U448 ( .A(n588), .ZN(n523) );
  XNOR2_X1 U449 ( .A(n534), .B(n533), .ZN(n662) );
  NAND2_X1 U450 ( .A1(G472), .A2(n376), .ZN(n375) );
  INV_X1 U451 ( .A(G902), .ZN(n376) );
  XNOR2_X1 U452 ( .A(n598), .B(KEYINPUT77), .ZN(n599) );
  INV_X1 U453 ( .A(KEYINPUT45), .ZN(n598) );
  XNOR2_X1 U454 ( .A(n479), .B(KEYINPUT10), .ZN(n719) );
  XNOR2_X1 U455 ( .A(n454), .B(n404), .ZN(n403) );
  INV_X1 U456 ( .A(G140), .ZN(n404) );
  XNOR2_X1 U457 ( .A(KEYINPUT91), .B(KEYINPUT24), .ZN(n454) );
  XNOR2_X1 U458 ( .A(G128), .B(G119), .ZN(n455) );
  XNOR2_X1 U459 ( .A(G137), .B(KEYINPUT90), .ZN(n457) );
  XOR2_X1 U460 ( .A(KEYINPUT23), .B(G110), .Z(n458) );
  XNOR2_X1 U461 ( .A(G116), .B(G107), .ZN(n490) );
  XNOR2_X1 U462 ( .A(n573), .B(n572), .ZN(n413) );
  NOR2_X1 U463 ( .A1(n413), .A2(n586), .ZN(n574) );
  XNOR2_X1 U464 ( .A(n478), .B(KEYINPUT73), .ZN(n542) );
  XNOR2_X1 U465 ( .A(n509), .B(n367), .ZN(n544) );
  XNOR2_X1 U466 ( .A(n508), .B(G475), .ZN(n367) );
  NAND2_X1 U467 ( .A1(n366), .A2(n545), .ZN(n588) );
  INV_X1 U468 ( .A(n544), .ZN(n366) );
  XNOR2_X1 U469 ( .A(n416), .B(n415), .ZN(n414) );
  XNOR2_X1 U470 ( .A(n436), .B(n438), .ZN(n415) );
  XNOR2_X1 U471 ( .A(n609), .B(KEYINPUT120), .ZN(n610) );
  XNOR2_X1 U472 ( .A(n684), .B(n683), .ZN(n685) );
  INV_X1 U473 ( .A(n363), .ZN(n551) );
  XNOR2_X1 U474 ( .A(n538), .B(KEYINPUT42), .ZN(n539) );
  INV_X1 U475 ( .A(KEYINPUT107), .ZN(n538) );
  NAND2_X1 U476 ( .A1(n528), .A2(n569), .ZN(n638) );
  XNOR2_X1 U477 ( .A(n568), .B(KEYINPUT32), .ZN(n428) );
  NOR2_X1 U478 ( .A1(n426), .A2(n581), .ZN(n615) );
  XNOR2_X1 U479 ( .A(n701), .B(n702), .ZN(n387) );
  XNOR2_X1 U480 ( .A(n695), .B(n696), .ZN(n386) );
  AND2_X1 U481 ( .A1(n571), .A2(n368), .ZN(n353) );
  AND2_X1 U482 ( .A1(n652), .A2(n426), .ZN(n354) );
  XOR2_X1 U483 ( .A(KEYINPUT3), .B(KEYINPUT68), .Z(n355) );
  XOR2_X1 U484 ( .A(KEYINPUT85), .B(G107), .Z(n356) );
  XOR2_X1 U485 ( .A(n458), .B(n457), .Z(n357) );
  OR2_X2 U486 ( .A1(n675), .A2(n674), .ZN(n358) );
  NAND2_X1 U487 ( .A1(n394), .A2(n589), .ZN(n359) );
  INV_X1 U488 ( .A(G472), .ZN(n378) );
  NOR2_X1 U489 ( .A1(KEYINPUT44), .A2(n349), .ZN(n360) );
  XNOR2_X1 U490 ( .A(n466), .B(n465), .ZN(n646) );
  XOR2_X1 U491 ( .A(n588), .B(KEYINPUT101), .Z(n630) );
  INV_X1 U492 ( .A(n630), .ZN(n369) );
  NOR2_X1 U493 ( .A1(n676), .A2(n413), .ZN(n361) );
  OR2_X1 U494 ( .A1(n674), .A2(n602), .ZN(n362) );
  INV_X1 U495 ( .A(n703), .ZN(n687) );
  NOR2_X1 U496 ( .A1(G902), .A2(n691), .ZN(n474) );
  XNOR2_X1 U497 ( .A(n721), .B(n470), .ZN(n384) );
  BUF_X2 U498 ( .A(n541), .Z(n363) );
  NOR2_X1 U499 ( .A1(n548), .A2(n405), .ZN(n525) );
  XNOR2_X2 U500 ( .A(G143), .B(G128), .ZN(n481) );
  NOR2_X1 U501 ( .A1(n439), .A2(n375), .ZN(n372) );
  AND2_X2 U502 ( .A1(n603), .A2(n358), .ZN(n694) );
  NAND2_X1 U503 ( .A1(n352), .A2(KEYINPUT44), .ZN(n595) );
  NOR2_X2 U504 ( .A1(n713), .A2(n602), .ZN(n601) );
  XNOR2_X2 U505 ( .A(n600), .B(n599), .ZN(n713) );
  NAND2_X1 U506 ( .A1(n395), .A2(n362), .ZN(n603) );
  XNOR2_X1 U507 ( .A(n594), .B(n406), .ZN(n392) );
  NAND2_X1 U508 ( .A1(n385), .A2(n359), .ZN(n380) );
  XNOR2_X1 U509 ( .A(n532), .B(KEYINPUT40), .ZN(n418) );
  XNOR2_X1 U510 ( .A(n580), .B(KEYINPUT100), .ZN(n427) );
  NAND2_X1 U511 ( .A1(n427), .A2(n354), .ZN(n425) );
  XNOR2_X2 U512 ( .A(n355), .B(n431), .ZN(n485) );
  NAND2_X1 U513 ( .A1(n694), .A2(G475), .ZN(n611) );
  OR2_X2 U514 ( .A1(n570), .A2(n567), .ZN(n429) );
  XNOR2_X2 U515 ( .A(n449), .B(KEYINPUT84), .ZN(n602) );
  NAND2_X1 U516 ( .A1(n734), .A2(KEYINPUT44), .ZN(n385) );
  NOR2_X1 U517 ( .A1(n386), .A2(n703), .ZN(G54) );
  NOR2_X1 U518 ( .A1(n387), .A2(n703), .ZN(G66) );
  XNOR2_X1 U519 ( .A(n388), .B(n479), .ZN(n483) );
  XNOR2_X1 U520 ( .A(n422), .B(n424), .ZN(n388) );
  AND2_X1 U521 ( .A1(n389), .A2(n687), .ZN(G63) );
  XNOR2_X1 U522 ( .A(n697), .B(n390), .ZN(n389) );
  INV_X1 U523 ( .A(n698), .ZN(n390) );
  NAND2_X1 U524 ( .A1(n397), .A2(n396), .ZN(n395) );
  XNOR2_X1 U525 ( .A(n391), .B(n506), .ZN(n608) );
  XNOR2_X1 U526 ( .A(n505), .B(n507), .ZN(n391) );
  NAND2_X1 U527 ( .A1(n392), .A2(n360), .ZN(n593) );
  XNOR2_X1 U528 ( .A(n483), .B(n482), .ZN(n412) );
  XNOR2_X1 U529 ( .A(n601), .B(KEYINPUT76), .ZN(n397) );
  XNOR2_X1 U530 ( .A(n393), .B(KEYINPUT46), .ZN(n399) );
  NAND2_X1 U531 ( .A1(n557), .A2(n558), .ZN(n560) );
  NAND2_X1 U532 ( .A1(n633), .A2(n619), .ZN(n394) );
  NAND2_X1 U533 ( .A1(n398), .A2(n687), .ZN(n607) );
  XNOR2_X1 U534 ( .A(n604), .B(n605), .ZN(n398) );
  INV_X1 U535 ( .A(n736), .ZN(n401) );
  NAND2_X1 U536 ( .A1(n541), .A2(n659), .ZN(n405) );
  INV_X1 U537 ( .A(n733), .ZN(n407) );
  NAND2_X1 U538 ( .A1(n682), .A2(n602), .ZN(n488) );
  XNOR2_X1 U539 ( .A(n410), .B(n705), .ZN(n682) );
  XNOR2_X1 U540 ( .A(n412), .B(n484), .ZN(n410) );
  INV_X1 U541 ( .A(n652), .ZN(n585) );
  NOR2_X1 U542 ( .A1(n666), .A2(n413), .ZN(n667) );
  XNOR2_X1 U543 ( .A(n485), .B(n437), .ZN(n416) );
  XNOR2_X1 U544 ( .A(n418), .B(n735), .ZN(G33) );
  XNOR2_X2 U545 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n424) );
  INV_X1 U546 ( .A(n425), .ZN(n622) );
  INV_X1 U547 ( .A(n646), .ZN(n426) );
  XNOR2_X2 U548 ( .A(n429), .B(n428), .ZN(n733) );
  NOR2_X2 U549 ( .A1(n570), .A2(n569), .ZN(n580) );
  NOR2_X2 U550 ( .A1(n597), .A2(n596), .ZN(n600) );
  AND2_X1 U551 ( .A1(G210), .A2(n487), .ZN(n430) );
  XNOR2_X1 U552 ( .A(n435), .B(n434), .ZN(n436) );
  INV_X1 U553 ( .A(KEYINPUT105), .ZN(n533) );
  NOR2_X1 U554 ( .A1(n661), .A2(n562), .ZN(n563) );
  XNOR2_X1 U555 ( .A(n472), .B(n471), .ZN(n691) );
  INV_X1 U556 ( .A(KEYINPUT1), .ZN(n526) );
  XNOR2_X1 U557 ( .A(n461), .B(n460), .ZN(n699) );
  XOR2_X1 U558 ( .A(KEYINPUT83), .B(n606), .Z(n703) );
  XNOR2_X1 U559 ( .A(n540), .B(n539), .ZN(n732) );
  XNOR2_X1 U560 ( .A(G116), .B(G119), .ZN(n431) );
  XOR2_X1 U561 ( .A(KEYINPUT5), .B(KEYINPUT96), .Z(n433) );
  XNOR2_X1 U562 ( .A(G101), .B(KEYINPUT72), .ZN(n432) );
  XNOR2_X1 U563 ( .A(n433), .B(n432), .ZN(n437) );
  XNOR2_X1 U564 ( .A(G113), .B(G131), .ZN(n435) );
  NAND2_X1 U565 ( .A1(n500), .A2(G210), .ZN(n438) );
  XOR2_X1 U566 ( .A(KEYINPUT30), .B(KEYINPUT102), .Z(n442) );
  XNOR2_X1 U567 ( .A(n440), .B(KEYINPUT71), .ZN(n487) );
  NAND2_X1 U568 ( .A1(G214), .A2(n487), .ZN(n659) );
  XNOR2_X1 U569 ( .A(n442), .B(n441), .ZN(n477) );
  XNOR2_X1 U570 ( .A(n443), .B(KEYINPUT14), .ZN(n445) );
  NAND2_X1 U571 ( .A1(n445), .A2(G952), .ZN(n444) );
  XOR2_X1 U572 ( .A(KEYINPUT87), .B(n444), .Z(n672) );
  NOR2_X1 U573 ( .A1(G953), .A2(n672), .ZN(n554) );
  NAND2_X1 U574 ( .A1(n445), .A2(G902), .ZN(n446) );
  XOR2_X1 U575 ( .A(KEYINPUT88), .B(n446), .Z(n553) );
  NAND2_X1 U576 ( .A1(n553), .A2(G953), .ZN(n447) );
  NOR2_X1 U577 ( .A1(G900), .A2(n447), .ZN(n448) );
  NOR2_X1 U578 ( .A1(n554), .A2(n448), .ZN(n510) );
  XOR2_X1 U579 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n452) );
  NAND2_X1 U580 ( .A1(n602), .A2(G234), .ZN(n450) );
  XNOR2_X1 U581 ( .A(n450), .B(KEYINPUT20), .ZN(n462) );
  NAND2_X1 U582 ( .A1(G221), .A2(n462), .ZN(n451) );
  XNOR2_X1 U583 ( .A(n452), .B(n451), .ZN(n453) );
  NAND2_X1 U584 ( .A1(G234), .A2(n724), .ZN(n456) );
  XOR2_X1 U585 ( .A(KEYINPUT8), .B(n456), .Z(n494) );
  NAND2_X1 U586 ( .A1(G221), .A2(n494), .ZN(n459) );
  NOR2_X1 U587 ( .A1(n699), .A2(G902), .ZN(n466) );
  XOR2_X1 U588 ( .A(KEYINPUT25), .B(KEYINPUT74), .Z(n464) );
  NAND2_X1 U589 ( .A1(G217), .A2(n462), .ZN(n463) );
  XOR2_X1 U590 ( .A(n464), .B(n463), .Z(n465) );
  NAND2_X1 U591 ( .A1(n561), .A2(n646), .ZN(n641) );
  INV_X1 U592 ( .A(n641), .ZN(n475) );
  XNOR2_X1 U593 ( .A(G101), .B(G110), .ZN(n467) );
  XNOR2_X2 U594 ( .A(n356), .B(n467), .ZN(n704) );
  NAND2_X1 U595 ( .A1(G227), .A2(n724), .ZN(n469) );
  XNOR2_X1 U596 ( .A(n504), .B(KEYINPUT89), .ZN(n721) );
  XNOR2_X1 U597 ( .A(KEYINPUT67), .B(G469), .ZN(n473) );
  XNOR2_X2 U598 ( .A(n474), .B(n473), .ZN(n527) );
  NAND2_X1 U599 ( .A1(n475), .A2(n527), .ZN(n582) );
  NOR2_X1 U600 ( .A1(n510), .A2(n582), .ZN(n476) );
  NAND2_X1 U601 ( .A1(n477), .A2(n476), .ZN(n478) );
  XOR2_X1 U602 ( .A(n480), .B(n481), .Z(n482) );
  XOR2_X1 U603 ( .A(G113), .B(G104), .Z(n486) );
  XOR2_X1 U604 ( .A(G122), .B(n486), .Z(n507) );
  AND2_X1 U605 ( .A1(n542), .A2(n658), .ZN(n489) );
  XNOR2_X1 U606 ( .A(n489), .B(KEYINPUT39), .ZN(n531) );
  XOR2_X1 U607 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n491) );
  XNOR2_X1 U608 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U609 ( .A(n493), .B(n492), .ZN(n498) );
  XOR2_X1 U610 ( .A(G122), .B(KEYINPUT98), .Z(n496) );
  NAND2_X1 U611 ( .A1(G217), .A2(n494), .ZN(n495) );
  XNOR2_X1 U612 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U613 ( .A(n498), .B(n497), .ZN(n698) );
  NOR2_X1 U614 ( .A1(G902), .A2(n698), .ZN(n499) );
  XNOR2_X1 U615 ( .A(G478), .B(n499), .ZN(n545) );
  INV_X1 U616 ( .A(n545), .ZN(n515) );
  NAND2_X1 U617 ( .A1(G214), .A2(n500), .ZN(n501) );
  XNOR2_X1 U618 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U619 ( .A(n503), .B(KEYINPUT12), .Z(n506) );
  XNOR2_X1 U620 ( .A(n719), .B(n504), .ZN(n505) );
  NOR2_X1 U621 ( .A1(G902), .A2(n608), .ZN(n509) );
  XNOR2_X1 U622 ( .A(KEYINPUT13), .B(KEYINPUT97), .ZN(n508) );
  NAND2_X1 U623 ( .A1(n515), .A2(n544), .ZN(n634) );
  NOR2_X1 U624 ( .A1(n531), .A2(n634), .ZN(n639) );
  INV_X1 U625 ( .A(KEYINPUT70), .ZN(n519) );
  NOR2_X1 U626 ( .A1(n519), .A2(KEYINPUT47), .ZN(n518) );
  NOR2_X1 U627 ( .A1(n646), .A2(n510), .ZN(n511) );
  NAND2_X1 U628 ( .A1(n645), .A2(n511), .ZN(n524) );
  NOR2_X1 U629 ( .A1(n652), .A2(n524), .ZN(n512) );
  XNOR2_X1 U630 ( .A(KEYINPUT28), .B(n512), .ZN(n513) );
  NAND2_X1 U631 ( .A1(n513), .A2(n527), .ZN(n537) );
  INV_X1 U632 ( .A(n557), .ZN(n514) );
  NOR2_X1 U633 ( .A1(n537), .A2(n514), .ZN(n627) );
  INV_X1 U634 ( .A(n634), .ZN(n623) );
  NOR2_X1 U635 ( .A1(n623), .A2(n523), .ZN(n663) );
  INV_X1 U636 ( .A(n663), .ZN(n516) );
  NAND2_X1 U637 ( .A1(n627), .A2(n516), .ZN(n517) );
  XNOR2_X1 U638 ( .A(n518), .B(n517), .ZN(n530) );
  NAND2_X1 U639 ( .A1(n519), .A2(KEYINPUT47), .ZN(n529) );
  INV_X1 U640 ( .A(KEYINPUT99), .ZN(n521) );
  XNOR2_X1 U641 ( .A(n525), .B(KEYINPUT36), .ZN(n528) );
  INV_X1 U642 ( .A(n642), .ZN(n569) );
  NOR2_X1 U643 ( .A1(n531), .A2(n588), .ZN(n532) );
  NAND2_X1 U644 ( .A1(n545), .A2(n544), .ZN(n661) );
  NAND2_X1 U645 ( .A1(n658), .A2(n659), .ZN(n534) );
  XNOR2_X1 U646 ( .A(KEYINPUT106), .B(KEYINPUT41), .ZN(n535) );
  XNOR2_X1 U647 ( .A(n536), .B(n535), .ZN(n676) );
  NOR2_X1 U648 ( .A1(n537), .A2(n676), .ZN(n540) );
  NAND2_X1 U649 ( .A1(n542), .A2(n363), .ZN(n543) );
  XNOR2_X1 U650 ( .A(KEYINPUT103), .B(n543), .ZN(n546) );
  NOR2_X1 U651 ( .A1(n545), .A2(n544), .ZN(n575) );
  NAND2_X1 U652 ( .A1(n546), .A2(n575), .ZN(n547) );
  XNOR2_X1 U653 ( .A(KEYINPUT104), .B(n547), .ZN(n736) );
  NOR2_X1 U654 ( .A1(n569), .A2(n548), .ZN(n549) );
  NAND2_X1 U655 ( .A1(n549), .A2(n659), .ZN(n550) );
  XNOR2_X1 U656 ( .A(KEYINPUT43), .B(n550), .ZN(n552) );
  NAND2_X1 U657 ( .A1(n552), .A2(n551), .ZN(n640) );
  INV_X1 U658 ( .A(KEYINPUT66), .ZN(n568) );
  NOR2_X1 U659 ( .A1(G898), .A2(n724), .ZN(n708) );
  NAND2_X1 U660 ( .A1(n553), .A2(n708), .ZN(n556) );
  INV_X1 U661 ( .A(n554), .ZN(n555) );
  NAND2_X1 U662 ( .A1(n556), .A2(n555), .ZN(n558) );
  XOR2_X1 U663 ( .A(KEYINPUT81), .B(KEYINPUT0), .Z(n559) );
  INV_X1 U664 ( .A(n586), .ZN(n564) );
  INV_X1 U665 ( .A(n561), .ZN(n562) );
  NAND2_X1 U666 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U667 ( .A1(n646), .A2(n642), .ZN(n566) );
  NAND2_X1 U668 ( .A1(n579), .A2(n566), .ZN(n567) );
  XNOR2_X1 U669 ( .A(KEYINPUT78), .B(KEYINPUT35), .ZN(n578) );
  NAND2_X1 U670 ( .A1(n584), .A2(n571), .ZN(n573) );
  XOR2_X1 U671 ( .A(KEYINPUT82), .B(KEYINPUT33), .Z(n572) );
  XNOR2_X1 U672 ( .A(n574), .B(KEYINPUT34), .ZN(n576) );
  NAND2_X1 U673 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U674 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U675 ( .A1(n350), .A2(n582), .ZN(n583) );
  NAND2_X1 U676 ( .A1(n583), .A2(n652), .ZN(n619) );
  NAND2_X1 U677 ( .A1(n585), .A2(n351), .ZN(n653) );
  NAND2_X1 U678 ( .A1(n588), .A2(n634), .ZN(n589) );
  XNOR2_X1 U679 ( .A(n591), .B(n590), .ZN(n592) );
  NAND2_X1 U680 ( .A1(n593), .A2(n592), .ZN(n597) );
  INV_X1 U681 ( .A(KEYINPUT2), .ZN(n674) );
  OR2_X2 U682 ( .A1(n723), .A2(n713), .ZN(n675) );
  NAND2_X1 U683 ( .A1(n694), .A2(G472), .ZN(n604) );
  NOR2_X1 U684 ( .A1(G952), .A2(n724), .ZN(n606) );
  XNOR2_X1 U685 ( .A(n607), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U686 ( .A(n608), .B(KEYINPUT59), .ZN(n609) );
  XNOR2_X1 U687 ( .A(n611), .B(n610), .ZN(n612) );
  NAND2_X1 U688 ( .A1(n612), .A2(n687), .ZN(n614) );
  INV_X1 U689 ( .A(KEYINPUT60), .ZN(n613) );
  XNOR2_X1 U690 ( .A(n614), .B(n613), .ZN(G60) );
  XOR2_X1 U691 ( .A(G101), .B(n615), .Z(G3) );
  NOR2_X1 U692 ( .A1(n630), .A2(n619), .ZN(n616) );
  XOR2_X1 U693 ( .A(G104), .B(n616), .Z(G6) );
  XOR2_X1 U694 ( .A(KEYINPUT108), .B(KEYINPUT26), .Z(n618) );
  XNOR2_X1 U695 ( .A(G107), .B(KEYINPUT27), .ZN(n617) );
  XNOR2_X1 U696 ( .A(n618), .B(n617), .ZN(n621) );
  NOR2_X1 U697 ( .A1(n634), .A2(n619), .ZN(n620) );
  XOR2_X1 U698 ( .A(n621), .B(n620), .Z(G9) );
  XOR2_X1 U699 ( .A(G110), .B(n622), .Z(G12) );
  XOR2_X1 U700 ( .A(KEYINPUT29), .B(KEYINPUT109), .Z(n625) );
  NAND2_X1 U701 ( .A1(n627), .A2(n623), .ZN(n624) );
  XNOR2_X1 U702 ( .A(n625), .B(n624), .ZN(n626) );
  XOR2_X1 U703 ( .A(G128), .B(n626), .Z(G30) );
  NAND2_X1 U704 ( .A1(n627), .A2(n369), .ZN(n628) );
  XNOR2_X1 U705 ( .A(n628), .B(KEYINPUT110), .ZN(n629) );
  XNOR2_X1 U706 ( .A(G146), .B(n629), .ZN(G48) );
  NOR2_X1 U707 ( .A1(n630), .A2(n633), .ZN(n632) );
  XNOR2_X1 U708 ( .A(G113), .B(KEYINPUT111), .ZN(n631) );
  XNOR2_X1 U709 ( .A(n632), .B(n631), .ZN(G15) );
  NOR2_X1 U710 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U711 ( .A(KEYINPUT112), .B(n635), .Z(n636) );
  XNOR2_X1 U712 ( .A(G116), .B(n636), .ZN(G18) );
  XOR2_X1 U713 ( .A(G125), .B(KEYINPUT37), .Z(n637) );
  XNOR2_X1 U714 ( .A(n638), .B(n637), .ZN(G27) );
  XOR2_X1 U715 ( .A(G134), .B(n639), .Z(G36) );
  XNOR2_X1 U716 ( .A(G140), .B(n640), .ZN(G42) );
  XOR2_X1 U717 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n644) );
  NAND2_X1 U718 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U719 ( .A(n644), .B(n643), .ZN(n650) );
  XOR2_X1 U720 ( .A(KEYINPUT49), .B(KEYINPUT113), .Z(n648) );
  OR2_X1 U721 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U722 ( .A(n648), .B(n647), .ZN(n649) );
  NOR2_X1 U723 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U724 ( .A1(n652), .A2(n651), .ZN(n654) );
  NAND2_X1 U725 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U726 ( .A(n655), .B(KEYINPUT51), .ZN(n656) );
  XOR2_X1 U727 ( .A(KEYINPUT115), .B(n656), .Z(n657) );
  NOR2_X1 U728 ( .A1(n676), .A2(n657), .ZN(n668) );
  NOR2_X1 U729 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U730 ( .A1(n661), .A2(n660), .ZN(n665) );
  NOR2_X1 U731 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U732 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U733 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U734 ( .A(n669), .B(KEYINPUT52), .ZN(n670) );
  XNOR2_X1 U735 ( .A(KEYINPUT116), .B(n670), .ZN(n671) );
  NOR2_X1 U736 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U737 ( .A(KEYINPUT117), .B(n673), .ZN(n679) );
  XOR2_X1 U738 ( .A(n675), .B(n674), .Z(n677) );
  NOR2_X1 U739 ( .A1(n677), .A2(n361), .ZN(n678) );
  NAND2_X1 U740 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U741 ( .A1(n680), .A2(G953), .ZN(n681) );
  XNOR2_X1 U742 ( .A(n681), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U743 ( .A1(n694), .A2(G210), .ZN(n686) );
  XNOR2_X1 U744 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n684) );
  XNOR2_X1 U745 ( .A(n682), .B(KEYINPUT75), .ZN(n683) );
  XNOR2_X1 U746 ( .A(n686), .B(n685), .ZN(n688) );
  NAND2_X1 U747 ( .A1(n688), .A2(n687), .ZN(n690) );
  XOR2_X1 U748 ( .A(KEYINPUT56), .B(KEYINPUT118), .Z(n689) );
  XNOR2_X1 U749 ( .A(n690), .B(n689), .ZN(G51) );
  XNOR2_X1 U750 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n693) );
  XNOR2_X1 U751 ( .A(n691), .B(KEYINPUT57), .ZN(n692) );
  XNOR2_X1 U752 ( .A(n693), .B(n692), .ZN(n696) );
  BUF_X2 U753 ( .A(n694), .Z(n700) );
  NAND2_X1 U754 ( .A1(n700), .A2(G469), .ZN(n695) );
  NAND2_X1 U755 ( .A1(n700), .A2(G478), .ZN(n697) );
  XOR2_X1 U756 ( .A(n699), .B(KEYINPUT121), .Z(n702) );
  NAND2_X1 U757 ( .A1(n700), .A2(G217), .ZN(n701) );
  XNOR2_X1 U758 ( .A(n704), .B(KEYINPUT124), .ZN(n706) );
  XNOR2_X1 U759 ( .A(n706), .B(n705), .ZN(n707) );
  NOR2_X1 U760 ( .A1(n708), .A2(n707), .ZN(n718) );
  NAND2_X1 U761 ( .A1(G224), .A2(G953), .ZN(n709) );
  XNOR2_X1 U762 ( .A(n709), .B(KEYINPUT122), .ZN(n710) );
  XNOR2_X1 U763 ( .A(KEYINPUT61), .B(n710), .ZN(n711) );
  NAND2_X1 U764 ( .A1(n711), .A2(G898), .ZN(n712) );
  XNOR2_X1 U765 ( .A(n712), .B(KEYINPUT123), .ZN(n715) );
  NOR2_X1 U766 ( .A1(n713), .A2(G953), .ZN(n714) );
  NOR2_X1 U767 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U768 ( .A(n716), .B(KEYINPUT125), .ZN(n717) );
  XNOR2_X1 U769 ( .A(n718), .B(n717), .ZN(G69) );
  XNOR2_X1 U770 ( .A(n720), .B(n719), .ZN(n722) );
  XNOR2_X1 U771 ( .A(n722), .B(n721), .ZN(n726) );
  XNOR2_X1 U772 ( .A(n726), .B(n723), .ZN(n725) );
  NAND2_X1 U773 ( .A1(n725), .A2(n724), .ZN(n730) );
  XNOR2_X1 U774 ( .A(G227), .B(n726), .ZN(n727) );
  NAND2_X1 U775 ( .A1(n727), .A2(G900), .ZN(n728) );
  NAND2_X1 U776 ( .A1(G953), .A2(n728), .ZN(n729) );
  NAND2_X1 U777 ( .A1(n730), .A2(n729), .ZN(G72) );
  XOR2_X1 U778 ( .A(G137), .B(KEYINPUT126), .Z(n731) );
  XNOR2_X1 U779 ( .A(n732), .B(n731), .ZN(G39) );
  XOR2_X1 U780 ( .A(n733), .B(G119), .Z(G21) );
  XOR2_X1 U781 ( .A(n349), .B(G122), .Z(G24) );
  XNOR2_X1 U782 ( .A(G131), .B(KEYINPUT127), .ZN(n735) );
  XNOR2_X1 U783 ( .A(G143), .B(n736), .ZN(G45) );
endmodule

