//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 1 0 0 1 1 0 0 0 1 0 0 0 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 0 1 1 1 1 0 0 1 0 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1327,
    new_n1328, new_n1329, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1399, new_n1400, new_n1401,
    new_n1402, new_n1403, new_n1404, new_n1405, new_n1406, new_n1407,
    new_n1408, new_n1409;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  XNOR2_X1  g0013(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n208), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n202), .A2(new_n203), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G50), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(new_n213), .A2(new_n214), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n220), .B1(new_n213), .B2(new_n214), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  INV_X1    g0023(.A(G87), .ZN(new_n224));
  INV_X1    g0024(.A(G250), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n222), .B1(new_n203), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n227));
  INV_X1    g0027(.A(G77), .ZN(new_n228));
  INV_X1    g0028(.A(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G107), .ZN(new_n230));
  INV_X1    g0030(.A(G264), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n227), .B1(new_n228), .B2(new_n229), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n210), .B1(new_n226), .B2(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT1), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n221), .A2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XOR2_X1   g0043(.A(G50), .B(G68), .Z(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(G13), .ZN(new_n251));
  NOR3_X1   g0051(.A1(new_n251), .A2(new_n208), .A3(G1), .ZN(new_n252));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n215), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n208), .A2(G1), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(KEYINPUT67), .A3(G50), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT67), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n259), .B1(new_n256), .B2(new_n201), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n255), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n252), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n261), .B1(G50), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n254), .ZN(new_n264));
  XOR2_X1   g0064(.A(KEYINPUT8), .B(G58), .Z(new_n265));
  NAND2_X1  g0065(.A1(new_n208), .A2(G33), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(G20), .A2(G33), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n265), .A2(new_n267), .B1(G150), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n204), .A2(G20), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n264), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n263), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT9), .ZN(new_n273));
  XNOR2_X1  g0073(.A(new_n272), .B(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT65), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G41), .A2(G45), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n275), .B1(new_n276), .B2(G1), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n207), .B(KEYINPUT65), .C1(G41), .C2(G45), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G274), .ZN(new_n280));
  AND2_X1   g0080(.A1(G1), .A2(G13), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AND2_X1   g0083(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G41), .ZN(new_n285));
  INV_X1    g0085(.A(G45), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n207), .A2(new_n287), .B1(new_n281), .B2(new_n282), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT66), .B(G226), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n284), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT3), .B(G33), .ZN(new_n291));
  INV_X1    g0091(.A(G1698), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n291), .A2(G222), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(G1698), .ZN(new_n294));
  INV_X1    g0094(.A(G223), .ZN(new_n295));
  OAI221_X1 g0095(.A(new_n293), .B1(new_n228), .B2(new_n291), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n290), .A2(new_n298), .A3(G190), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n290), .A2(new_n298), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G200), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n274), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT10), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT10), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n274), .A2(new_n304), .A3(new_n299), .A4(new_n301), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT68), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n255), .A2(G77), .A3(new_n257), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n308), .B1(G77), .B2(new_n262), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n265), .A2(new_n268), .B1(G20), .B2(G77), .ZN(new_n310));
  XNOR2_X1  g0110(.A(KEYINPUT15), .B(G87), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n267), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n264), .B1(new_n310), .B2(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n309), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n284), .B1(G244), .B2(new_n288), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n291), .A2(G232), .A3(new_n292), .ZN(new_n317));
  OAI221_X1 g0117(.A(new_n317), .B1(new_n230), .B2(new_n291), .C1(new_n294), .C2(new_n223), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n297), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G169), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n315), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G179), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n316), .A2(new_n319), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G190), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n315), .B1(new_n320), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G200), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(new_n316), .B2(new_n319), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n307), .B1(new_n326), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n272), .B1(new_n300), .B2(new_n321), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(G179), .B2(new_n300), .ZN(new_n334));
  INV_X1    g0134(.A(new_n331), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n335), .A2(KEYINPUT68), .A3(new_n325), .ZN(new_n336));
  AND4_X1   g0136(.A1(new_n306), .A2(new_n332), .A3(new_n334), .A4(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n255), .A2(G68), .A3(new_n257), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT70), .ZN(new_n339));
  XNOR2_X1  g0139(.A(new_n338), .B(new_n339), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n268), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(new_n228), .B2(new_n266), .ZN(new_n342));
  AND2_X1   g0142(.A1(new_n342), .A2(new_n254), .ZN(new_n343));
  OR2_X1    g0143(.A1(new_n343), .A2(KEYINPUT11), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n252), .A2(new_n203), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n345), .B(KEYINPUT12), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n343), .A2(KEYINPUT11), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n340), .A2(new_n344), .A3(new_n346), .A4(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT14), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n291), .A2(G232), .A3(G1698), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n291), .A2(G226), .A3(new_n292), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT69), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n352), .B1(G33), .B2(G97), .ZN(new_n353));
  NAND2_X1  g0153(.A1(G33), .A2(G97), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n354), .A2(KEYINPUT69), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n350), .A2(new_n351), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n297), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT13), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n279), .A2(new_n283), .B1(new_n288), .B2(G238), .ZN(new_n360));
  AND3_X1   g0160(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n359), .B1(new_n358), .B2(new_n360), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n349), .B(G169), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n358), .A2(new_n360), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT13), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n365), .A2(G179), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n365), .A2(new_n366), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n349), .B1(new_n369), .B2(G169), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n348), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n348), .ZN(new_n373));
  OAI21_X1  g0173(.A(G200), .B1(new_n361), .B2(new_n362), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n365), .A2(G190), .A3(new_n366), .ZN(new_n375));
  AND3_X1   g0175(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n372), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT73), .ZN(new_n378));
  INV_X1    g0178(.A(new_n265), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n379), .A2(new_n256), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n380), .A2(new_n255), .B1(new_n252), .B2(new_n379), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G33), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT3), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT3), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(G33), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT7), .B1(new_n387), .B2(new_n208), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT7), .ZN(new_n389));
  AOI211_X1 g0189(.A(new_n389), .B(G20), .C1(new_n384), .C2(new_n386), .ZN(new_n390));
  OAI21_X1  g0190(.A(G68), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(G159), .ZN(new_n392));
  NOR3_X1   g0192(.A1(new_n392), .A2(G20), .A3(G33), .ZN(new_n393));
  NAND2_X1  g0193(.A1(G58), .A2(G68), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT71), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT71), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n396), .A2(G58), .A3(G68), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n395), .A2(new_n397), .A3(new_n217), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n393), .B1(new_n398), .B2(G20), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n391), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT16), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n264), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n398), .A2(G20), .ZN(new_n403));
  INV_X1    g0203(.A(new_n393), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT72), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT72), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n399), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n406), .A2(KEYINPUT16), .A3(new_n391), .A4(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n382), .B1(new_n402), .B2(new_n409), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n384), .A2(new_n386), .A3(G226), .A4(G1698), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n384), .A2(new_n386), .A3(G223), .A4(new_n292), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G33), .A2(G87), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n297), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n279), .A2(new_n283), .B1(new_n288), .B2(G232), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n321), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n415), .A2(new_n416), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n417), .B1(G179), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(KEYINPUT18), .B1(new_n410), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n389), .B1(new_n291), .B2(G20), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n387), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n401), .B1(new_n423), .B2(G68), .ZN(new_n424));
  AND3_X1   g0224(.A1(new_n424), .A2(new_n406), .A3(new_n408), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n203), .B1(new_n421), .B2(new_n422), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n401), .B1(new_n426), .B2(new_n405), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n254), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n381), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT18), .ZN(new_n430));
  INV_X1    g0230(.A(new_n419), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n378), .B1(new_n420), .B2(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(KEYINPUT73), .A2(KEYINPUT18), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(new_n410), .B2(new_n419), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n409), .A2(new_n254), .A3(new_n427), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n415), .A2(new_n416), .A3(G190), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n329), .B1(new_n415), .B2(new_n416), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n436), .A2(new_n381), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT17), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n436), .A2(new_n439), .A3(KEYINPUT17), .A4(new_n381), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n435), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n433), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n337), .A2(new_n377), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT25), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n262), .A2(new_n448), .A3(G107), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n448), .B1(new_n262), .B2(G107), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n207), .A2(G33), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n255), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n452), .B1(new_n230), .B2(new_n454), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n384), .A2(new_n386), .A3(new_n208), .A4(G87), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT22), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT22), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n291), .A2(new_n458), .A3(new_n208), .A4(G87), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(G33), .A2(G116), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(G20), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT23), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n463), .B1(new_n208), .B2(G107), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n230), .A2(KEYINPUT23), .A3(G20), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n460), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT24), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT24), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n460), .A2(new_n469), .A3(new_n466), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n455), .B1(new_n471), .B2(new_n254), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n384), .A2(new_n386), .A3(G257), .A4(G1698), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(KEYINPUT77), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT77), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n291), .A2(new_n475), .A3(G257), .A4(G1698), .ZN(new_n476));
  NAND2_X1  g0276(.A1(G33), .A2(G294), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n291), .A2(G250), .A3(new_n292), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n474), .A2(new_n476), .A3(new_n477), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n297), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n207), .A2(G45), .ZN(new_n481));
  OR2_X1    g0281(.A1(KEYINPUT5), .A2(G41), .ZN(new_n482));
  NAND2_X1  g0282(.A1(KEYINPUT5), .A2(G41), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NOR3_X1   g0284(.A1(new_n484), .A2(new_n231), .A3(new_n297), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n480), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT78), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n484), .A2(new_n283), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n485), .B1(new_n479), .B2(new_n297), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(KEYINPUT78), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n489), .A2(G179), .A3(new_n490), .A4(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n321), .B1(new_n491), .B2(new_n490), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n472), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n489), .A2(new_n490), .A3(new_n492), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n329), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n491), .A2(new_n327), .A3(new_n490), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n496), .B1(new_n500), .B2(new_n472), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n286), .A2(G1), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n281), .A2(new_n282), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n225), .B1(new_n207), .B2(G45), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n283), .A2(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(G238), .A2(G1698), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n506), .B1(new_n229), .B2(G1698), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n507), .A2(new_n291), .B1(G33), .B2(G116), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n323), .B(new_n505), .C1(new_n508), .C2(new_n503), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT75), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n223), .A2(new_n292), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n229), .A2(G1698), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n384), .A2(new_n511), .A3(new_n386), .A4(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n461), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n297), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT75), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n515), .A2(new_n516), .A3(new_n323), .A4(new_n505), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n503), .A2(new_n504), .ZN(new_n518));
  INV_X1    g0318(.A(new_n283), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n518), .B1(new_n519), .B2(new_n481), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n503), .B1(new_n513), .B2(new_n461), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n321), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n510), .A2(new_n517), .A3(new_n522), .ZN(new_n523));
  NOR3_X1   g0323(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n524));
  OAI21_X1  g0324(.A(KEYINPUT19), .B1(new_n353), .B2(new_n355), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n524), .B1(new_n525), .B2(new_n208), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n384), .A2(new_n386), .A3(new_n208), .A4(G68), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT19), .ZN(new_n528));
  INV_X1    g0328(.A(G97), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n528), .B1(new_n266), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n254), .B1(new_n526), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n312), .A2(new_n262), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n454), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n312), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n532), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT76), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n524), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n354), .A2(KEYINPUT69), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n352), .A2(G33), .A3(G97), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n528), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n540), .B1(new_n543), .B2(G20), .ZN(new_n544));
  AND2_X1   g0344(.A1(new_n527), .A2(new_n530), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n533), .B1(new_n546), .B2(new_n254), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n547), .A2(KEYINPUT76), .A3(new_n536), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n523), .A2(new_n539), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n515), .A2(G190), .A3(new_n505), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n535), .A2(G87), .ZN(new_n551));
  AND4_X1   g0351(.A1(new_n532), .A2(new_n550), .A3(new_n534), .A4(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n520), .A2(new_n521), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n552), .B1(new_n329), .B2(new_n553), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n483), .ZN(new_n556));
  NOR2_X1   g0356(.A1(KEYINPUT5), .A2(G41), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n502), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n558), .A2(G270), .A3(new_n503), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n490), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n384), .A2(new_n386), .A3(G257), .A4(new_n292), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n384), .A2(new_n386), .A3(G264), .A4(G1698), .ZN(new_n563));
  INV_X1    g0363(.A(G303), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n562), .B(new_n563), .C1(new_n564), .C2(new_n291), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n297), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n561), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n255), .A2(G116), .A3(new_n453), .ZN(new_n568));
  INV_X1    g0368(.A(G116), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n252), .A2(new_n569), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n253), .A2(new_n215), .B1(G20), .B2(new_n569), .ZN(new_n571));
  NAND2_X1  g0371(.A1(G33), .A2(G283), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n572), .B(new_n208), .C1(G33), .C2(new_n529), .ZN(new_n573));
  AOI21_X1  g0373(.A(KEYINPUT20), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  AND3_X1   g0374(.A1(new_n571), .A2(KEYINPUT20), .A3(new_n573), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n568), .B(new_n570), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n567), .A2(G169), .A3(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT21), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n576), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n561), .A2(new_n566), .A3(G190), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n560), .B1(new_n297), .B2(new_n565), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n580), .B(new_n581), .C1(new_n582), .C2(new_n329), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(G179), .A3(new_n576), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n567), .A2(KEYINPUT21), .A3(G169), .A4(new_n576), .ZN(new_n585));
  AND4_X1   g0385(.A1(new_n579), .A2(new_n583), .A3(new_n584), .A4(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n268), .A2(G77), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT6), .ZN(new_n588));
  NOR3_X1   g0388(.A1(new_n588), .A2(new_n529), .A3(G107), .ZN(new_n589));
  XNOR2_X1  g0389(.A(G97), .B(G107), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n589), .B1(new_n590), .B2(new_n588), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n587), .B1(new_n591), .B2(new_n208), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n230), .B1(new_n421), .B2(new_n422), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n254), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n262), .A2(G97), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n595), .B1(new_n535), .B2(G97), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n384), .A2(new_n386), .A3(G244), .A4(new_n292), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT4), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n291), .A2(KEYINPUT4), .A3(G244), .A4(new_n292), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n291), .A2(G250), .A3(G1698), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n600), .A2(new_n601), .A3(new_n572), .A4(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n297), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n558), .A2(G257), .A3(new_n503), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n490), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n597), .B1(G200), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(KEYINPUT74), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n606), .B1(new_n603), .B2(new_n297), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT74), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n610), .A2(G190), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  AOI211_X1 g0415(.A(KEYINPUT74), .B(new_n606), .C1(new_n297), .C2(new_n603), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n612), .B1(new_n604), .B2(new_n607), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n321), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n611), .A2(new_n323), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n597), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n586), .A2(new_n615), .A3(new_n621), .ZN(new_n622));
  AND4_X1   g0422(.A1(new_n447), .A2(new_n501), .A3(new_n555), .A4(new_n622), .ZN(G372));
  INV_X1    g0423(.A(new_n334), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n372), .B1(new_n625), .B2(new_n326), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n442), .A2(new_n443), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n420), .B(new_n432), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT80), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n306), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n303), .A2(KEYINPUT80), .A3(new_n305), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n624), .B1(new_n628), .B2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT26), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n597), .A2(new_n619), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n610), .A2(new_n613), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n635), .B1(new_n636), .B2(new_n321), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n634), .B1(new_n555), .B2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT79), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(new_n508), .B2(new_n503), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n521), .A2(KEYINPUT79), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n520), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n537), .B(new_n509), .C1(G169), .C2(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n521), .A2(KEYINPUT79), .ZN(new_n644));
  AOI211_X1 g0444(.A(new_n639), .B(new_n503), .C1(new_n513), .C2(new_n461), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n505), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(G200), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n552), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n618), .A2(new_n648), .A3(new_n620), .A4(new_n643), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n643), .B1(new_n649), .B2(KEYINPUT26), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n638), .A2(new_n650), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n646), .A2(new_n321), .B1(new_n323), .B2(new_n553), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n652), .A2(new_n537), .B1(new_n552), .B2(new_n647), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n615), .A2(new_n621), .A3(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n491), .A2(KEYINPUT78), .ZN(new_n655));
  AOI211_X1 g0455(.A(new_n488), .B(new_n485), .C1(new_n479), .C2(new_n297), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(G200), .B1(new_n657), .B2(new_n490), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n491), .A2(new_n490), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(G190), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n472), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n579), .A2(new_n584), .A3(new_n585), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n654), .B(new_n661), .C1(new_n496), .C2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n651), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n633), .B1(new_n446), .B2(new_n665), .ZN(G369));
  NAND2_X1  g0466(.A1(new_n471), .A2(new_n254), .ZN(new_n667));
  INV_X1    g0467(.A(new_n455), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n490), .A2(G179), .ZN(new_n670));
  NOR3_X1   g0470(.A1(new_n655), .A2(new_n656), .A3(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n669), .B1(new_n671), .B2(new_n494), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT81), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n675));
  INV_X1    g0475(.A(G213), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT82), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(KEYINPUT82), .B1(new_n674), .B2(KEYINPUT27), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n677), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  XOR2_X1   g0482(.A(KEYINPUT83), .B(G343), .Z(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n669), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n660), .B1(new_n497), .B2(new_n329), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n672), .B(new_n685), .C1(new_n686), .C2(new_n669), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT84), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT84), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n661), .A2(new_n689), .A3(new_n672), .A4(new_n685), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n496), .A2(new_n684), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n684), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(new_n580), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n662), .ZN(new_n697));
  INV_X1    g0497(.A(new_n586), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n697), .B1(new_n698), .B2(new_n696), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(G330), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n694), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n662), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(new_n684), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n688), .A2(new_n690), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n496), .A2(new_n695), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n701), .A2(new_n706), .ZN(G399));
  INV_X1    g0507(.A(new_n211), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(G41), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n540), .A2(G116), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n710), .A2(G1), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n218), .B2(new_n710), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT28), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n501), .A2(new_n622), .A3(new_n555), .A4(new_n695), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT30), .ZN(new_n716));
  AND4_X1   g0516(.A1(G179), .A2(new_n553), .A3(new_n566), .A4(new_n561), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n489), .A2(new_n717), .A3(new_n492), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n716), .B1(new_n718), .B2(new_n636), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n616), .A2(new_n617), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n657), .A2(new_n720), .A3(KEYINPUT30), .A4(new_n717), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n642), .A2(new_n582), .A3(G179), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n497), .A2(new_n608), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n719), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(new_n684), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT31), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n724), .A2(KEYINPUT31), .A3(new_n684), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n715), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G330), .ZN(new_n730));
  OAI21_X1  g0530(.A(KEYINPUT85), .B1(new_n496), .B2(new_n662), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT85), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n672), .A2(new_n702), .A3(new_n732), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n731), .A2(new_n654), .A3(new_n733), .A4(new_n661), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n637), .A2(new_n634), .A3(new_n554), .A4(new_n549), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n509), .B1(new_n642), .B2(G169), .ZN(new_n736));
  INV_X1    g0536(.A(new_n537), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n642), .A2(new_n329), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n532), .A2(new_n550), .A3(new_n551), .A4(new_n534), .ZN(new_n739));
  OAI22_X1  g0539(.A1(new_n736), .A2(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(KEYINPUT26), .B1(new_n621), .B2(new_n740), .ZN(new_n741));
  AND3_X1   g0541(.A1(new_n735), .A2(new_n643), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n684), .B1(new_n734), .B2(new_n742), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n743), .A2(KEYINPUT29), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n684), .B1(new_n651), .B2(new_n663), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(KEYINPUT29), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n730), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n714), .B1(new_n748), .B2(G1), .ZN(G364));
  NOR2_X1   g0549(.A1(new_n208), .A2(G179), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n750), .A2(new_n327), .A3(G200), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n291), .B1(new_n752), .B2(G283), .ZN(new_n753));
  INV_X1    g0553(.A(G294), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n327), .A2(G179), .A3(G200), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n208), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n750), .A2(new_n327), .A3(new_n329), .ZN(new_n757));
  OR2_X1    g0557(.A1(new_n757), .A2(KEYINPUT92), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(KEYINPUT92), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G329), .ZN(new_n761));
  OAI221_X1 g0561(.A(new_n753), .B1(new_n754), .B2(new_n756), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n750), .A2(G190), .A3(G200), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT91), .ZN(new_n764));
  OR2_X1    g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n763), .A2(new_n764), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(G20), .A2(G179), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT86), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(new_n327), .A3(G200), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(KEYINPUT33), .B(G317), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n768), .A2(G303), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G326), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n770), .A2(G190), .A3(G200), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT87), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n770), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(G200), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n770), .A2(new_n778), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n780), .A2(G190), .A3(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n762), .B(new_n777), .C1(G322), .C2(new_n783), .ZN(new_n784));
  AND3_X1   g0584(.A1(new_n780), .A2(new_n327), .A3(new_n781), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n785), .A2(KEYINPUT88), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(KEYINPUT88), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G311), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n784), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n782), .A2(new_n202), .B1(new_n201), .B2(new_n776), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n792), .B1(new_n788), .B2(G77), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT89), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n768), .A2(G87), .ZN(new_n795));
  XNOR2_X1  g0595(.A(KEYINPUT90), .B(G159), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n757), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT32), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n756), .A2(new_n529), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n751), .A2(new_n230), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n799), .A2(new_n800), .A3(new_n387), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n772), .A2(G68), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n795), .A2(new_n798), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n791), .B1(new_n794), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n215), .B1(G20), .B2(new_n321), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n251), .A2(G20), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n207), .B1(new_n807), .B2(G45), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n709), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n211), .A2(G355), .A3(new_n291), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n708), .A2(new_n291), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(G45), .B2(new_n218), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n246), .A2(new_n286), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n812), .B1(G116), .B2(new_n211), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(G13), .A2(G33), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(G20), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n819), .A2(new_n805), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n811), .B1(new_n816), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n819), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n806), .B(new_n821), .C1(new_n699), .C2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n700), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(new_n810), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(G330), .B2(new_n699), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n823), .A2(new_n826), .ZN(G396));
  NOR2_X1   g0627(.A1(new_n805), .A2(new_n817), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n811), .B1(new_n228), .B2(new_n828), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n829), .B(KEYINPUT93), .Z(new_n830));
  OAI21_X1  g0630(.A(new_n291), .B1(new_n751), .B2(new_n203), .ZN(new_n831));
  INV_X1    g0631(.A(new_n756), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n831), .B1(G58), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(G132), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n833), .B1(new_n767), .B2(new_n201), .C1(new_n834), .C2(new_n760), .ZN(new_n835));
  INV_X1    g0635(.A(G137), .ZN(new_n836));
  INV_X1    g0636(.A(G150), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n836), .A2(new_n776), .B1(new_n771), .B2(new_n837), .ZN(new_n838));
  XOR2_X1   g0638(.A(KEYINPUT95), .B(G143), .Z(new_n839));
  AOI21_X1  g0639(.A(new_n838), .B1(new_n783), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n789), .B2(new_n796), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT34), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n835), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n842), .B2(new_n841), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n751), .A2(new_n224), .ZN(new_n845));
  INV_X1    g0645(.A(new_n760), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n799), .B(new_n845), .C1(new_n846), .C2(G311), .ZN(new_n847));
  INV_X1    g0647(.A(G283), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n847), .B1(new_n848), .B2(new_n771), .C1(new_n564), .C2(new_n776), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n387), .B1(new_n767), .B2(new_n230), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n850), .B(KEYINPUT94), .Z(new_n851));
  NOR2_X1   g0651(.A1(new_n782), .A2(new_n754), .ZN(new_n852));
  NOR3_X1   g0652(.A1(new_n849), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n569), .B2(new_n789), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n844), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n805), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n830), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OR2_X1    g0657(.A1(new_n857), .A2(KEYINPUT96), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(KEYINPUT96), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n684), .B1(new_n314), .B2(new_n309), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n326), .B1(new_n335), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n325), .A2(new_n684), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n817), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n858), .A2(new_n859), .A3(new_n865), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n745), .B(new_n864), .ZN(new_n867));
  INV_X1    g0667(.A(new_n730), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XOR2_X1   g0669(.A(new_n869), .B(KEYINPUT97), .Z(new_n870));
  OAI21_X1  g0670(.A(new_n811), .B1(new_n867), .B2(new_n868), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n866), .B1(new_n870), .B2(new_n871), .ZN(G384));
  INV_X1    g0672(.A(new_n591), .ZN(new_n873));
  OR2_X1    g0673(.A1(new_n873), .A2(KEYINPUT35), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(KEYINPUT35), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n874), .A2(G116), .A3(new_n216), .A4(new_n875), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n876), .B(KEYINPUT36), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n219), .A2(G77), .A3(new_n397), .A4(new_n395), .ZN(new_n878));
  OAI22_X1  g0678(.A1(new_n878), .A2(KEYINPUT98), .B1(G50), .B2(new_n203), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(KEYINPUT98), .B2(new_n878), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n251), .A2(G1), .ZN(new_n881));
  INV_X1    g0681(.A(G330), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT101), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n407), .B1(new_n403), .B2(new_n404), .ZN(new_n884));
  AOI211_X1 g0684(.A(KEYINPUT72), .B(new_n393), .C1(new_n398), .C2(G20), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n264), .B1(new_n886), .B2(new_n424), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n406), .A2(new_n408), .A3(new_n391), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n401), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n382), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n440), .B1(new_n890), .B2(new_n419), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n682), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT37), .ZN(new_n894));
  INV_X1    g0694(.A(new_n682), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n429), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n429), .A2(new_n431), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n440), .B(new_n896), .C1(new_n897), .C2(KEYINPUT100), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT100), .B1(new_n410), .B2(new_n419), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n894), .ZN(new_n900));
  OAI22_X1  g0700(.A1(new_n893), .A2(new_n894), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n892), .B1(new_n433), .B2(new_n444), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n901), .A2(KEYINPUT38), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT38), .B1(new_n901), .B2(new_n902), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n883), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT38), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n409), .A2(new_n254), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT16), .B1(new_n886), .B2(new_n391), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n381), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n895), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n420), .A2(new_n432), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT73), .ZN(new_n912));
  AND3_X1   g0712(.A1(new_n435), .A2(new_n442), .A3(new_n443), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n440), .B1(new_n410), .B2(new_n682), .ZN(new_n915));
  NOR3_X1   g0715(.A1(new_n410), .A2(KEYINPUT100), .A3(new_n419), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT37), .B1(new_n897), .B2(KEYINPUT100), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n909), .A2(new_n431), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n910), .A2(new_n919), .A3(new_n440), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n917), .A2(new_n918), .B1(new_n920), .B2(KEYINPUT37), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n906), .B1(new_n914), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n901), .A2(new_n902), .A3(KEYINPUT38), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n922), .A2(KEYINPUT101), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n905), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n695), .A2(new_n373), .ZN(new_n926));
  OAI21_X1  g0726(.A(G169), .B1(new_n361), .B2(new_n362), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(KEYINPUT14), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n928), .A2(new_n367), .A3(new_n363), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n926), .B1(new_n929), .B2(new_n376), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(KEYINPUT99), .ZN(new_n931));
  INV_X1    g0731(.A(new_n926), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n371), .A2(new_n932), .A3(new_n625), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT99), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n934), .B(new_n926), .C1(new_n929), .C2(new_n376), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n931), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n863), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n715), .A2(new_n728), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT104), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n725), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n724), .A2(KEYINPUT104), .A3(new_n684), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n941), .A2(new_n726), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n937), .B1(new_n939), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT40), .B1(new_n925), .B2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT40), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n420), .A2(new_n442), .A3(new_n432), .A4(new_n443), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n682), .B1(new_n436), .B2(new_n381), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT103), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n947), .A2(KEYINPUT103), .A3(new_n948), .ZN(new_n952));
  AND3_X1   g0752(.A1(new_n436), .A2(new_n381), .A3(new_n439), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n953), .A2(new_n948), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n419), .B1(new_n436), .B2(new_n381), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT100), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n954), .A2(new_n894), .A3(new_n957), .A4(new_n899), .ZN(new_n958));
  OAI21_X1  g0758(.A(KEYINPUT37), .B1(new_n915), .B2(new_n955), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n951), .A2(new_n952), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n906), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n946), .B1(new_n962), .B2(new_n923), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n945), .B1(new_n944), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n446), .B1(new_n939), .B2(new_n943), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n882), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n964), .B2(new_n965), .ZN(new_n967));
  INV_X1    g0767(.A(new_n936), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n745), .A2(new_n863), .ZN(new_n969));
  INV_X1    g0769(.A(new_n862), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n968), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n925), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT39), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n949), .A2(new_n950), .B1(new_n958), .B2(new_n959), .ZN(new_n974));
  AOI21_X1  g0774(.A(KEYINPUT38), .B1(new_n974), .B2(new_n952), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n973), .B1(new_n975), .B2(new_n903), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n372), .A2(new_n695), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT102), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n922), .A2(KEYINPUT39), .A3(new_n923), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n976), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n911), .A2(new_n682), .ZN(new_n981));
  AND3_X1   g0781(.A1(new_n972), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n743), .A2(KEYINPUT29), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n447), .B(new_n983), .C1(KEYINPUT29), .C2(new_n745), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n633), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n982), .B(new_n985), .Z(new_n986));
  NAND2_X1  g0786(.A1(new_n967), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n207), .B2(new_n807), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n967), .A2(new_n986), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n877), .B1(new_n880), .B2(new_n881), .C1(new_n988), .C2(new_n989), .ZN(G367));
  INV_X1    g0790(.A(KEYINPUT46), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n767), .B2(new_n569), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT107), .Z(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(G303), .B2(new_n783), .ZN(new_n994));
  NOR3_X1   g0794(.A1(new_n767), .A2(new_n991), .A3(new_n569), .ZN(new_n995));
  INV_X1    g0795(.A(G317), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n387), .B1(new_n757), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(G107), .B2(new_n832), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n998), .B1(new_n529), .B2(new_n751), .C1(new_n790), .C2(new_n776), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n995), .B(new_n999), .C1(G294), .C2(new_n772), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n994), .B(new_n1000), .C1(new_n848), .C2(new_n789), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n767), .A2(new_n202), .B1(new_n771), .B2(new_n796), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n776), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n839), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n752), .A2(G77), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n832), .A2(G68), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n757), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n387), .B1(new_n1007), .B2(G137), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .A4(new_n1008), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n1002), .B(new_n1009), .C1(G150), .C2(new_n783), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n789), .B2(new_n201), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1001), .A2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT47), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n805), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n820), .B1(new_n211), .B2(new_n311), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(new_n813), .B2(new_n242), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n811), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n695), .B1(new_n547), .B2(new_n551), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n643), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n653), .B2(new_n1018), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT105), .Z(new_n1021));
  OAI211_X1 g0821(.A(new_n1014), .B(new_n1017), .C1(new_n822), .C2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n684), .A2(new_n597), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n615), .A2(new_n621), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n637), .A2(new_n684), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n704), .A2(new_n705), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT45), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n704), .A2(KEYINPUT45), .A3(new_n705), .A4(new_n1026), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1026), .ZN(new_n1032));
  AOI21_X1  g0832(.A(KEYINPUT44), .B1(new_n706), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT44), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n1034), .B(new_n1026), .C1(new_n704), .C2(new_n705), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1031), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n701), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n704), .B1(new_n693), .B2(new_n703), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n1038), .A2(new_n824), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n824), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n747), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n701), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1031), .B(new_n1042), .C1(new_n1033), .C2(new_n1035), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1037), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n748), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n709), .B(KEYINPUT41), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n809), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1042), .A2(new_n1032), .ZN(new_n1048));
  AND2_X1   g0848(.A1(new_n1021), .A2(KEYINPUT43), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1021), .A2(KEYINPUT43), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n688), .A2(new_n690), .A3(new_n703), .A4(new_n1026), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n1052), .A2(KEYINPUT42), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n621), .B1(new_n1024), .B2(new_n672), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n1052), .A2(KEYINPUT42), .B1(new_n695), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(KEYINPUT106), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT106), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1053), .A2(new_n1055), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1051), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1061), .A2(new_n1050), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1048), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1061), .B1(new_n1050), .B2(new_n1049), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1048), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1064), .B(new_n1065), .C1(new_n1061), .C2(new_n1050), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1022), .B1(new_n1047), .B2(new_n1067), .ZN(G387));
  OAI221_X1 g0868(.A(new_n387), .B1(new_n757), .B2(new_n775), .C1(new_n569), .C2(new_n751), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n768), .A2(G294), .B1(G283), .B2(new_n832), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G311), .A2(new_n772), .B1(new_n1003), .B2(G322), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n782), .B2(new_n996), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(new_n788), .B2(G303), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1070), .B1(new_n1073), .B2(KEYINPUT48), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(KEYINPUT48), .B2(new_n1073), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT49), .ZN(new_n1076));
  OR2_X1    g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1069), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n783), .A2(G50), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n772), .A2(new_n265), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n291), .B1(new_n757), .B2(new_n837), .C1(new_n529), .C2(new_n751), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n312), .B2(new_n832), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n768), .A2(G77), .B1(G159), .B2(new_n1003), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1080), .A2(new_n1081), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n788), .B2(G68), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n805), .B1(new_n1079), .B2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n239), .A2(new_n286), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n265), .A2(new_n201), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT50), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n711), .B(new_n286), .C1(new_n203), .C2(new_n228), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n813), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1088), .B1(KEYINPUT108), .B2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(KEYINPUT108), .B2(new_n1092), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n211), .A2(new_n291), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n1094), .B1(G107), .B2(new_n211), .C1(new_n711), .C2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n811), .B1(new_n1096), .B2(new_n820), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1087), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n694), .B2(new_n819), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1099), .B1(new_n809), .B2(new_n1100), .ZN(new_n1101));
  OR3_X1    g0901(.A1(new_n1100), .A2(KEYINPUT109), .A3(new_n748), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1041), .ZN(new_n1103));
  OAI21_X1  g0903(.A(KEYINPUT109), .B1(new_n1100), .B2(new_n748), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1102), .A2(new_n709), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1101), .A2(new_n1105), .ZN(G393));
  NAND2_X1  g0906(.A1(new_n1037), .A2(new_n1043), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n1103), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1108), .A2(new_n709), .A3(new_n1044), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1037), .A2(new_n1043), .A3(new_n809), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT111), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n813), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n820), .B1(new_n529), .B2(new_n211), .C1(new_n1112), .C2(new_n249), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n810), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n789), .A2(new_n379), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n782), .A2(new_n392), .B1(new_n837), .B2(new_n776), .ZN(new_n1116));
  XOR2_X1   g0916(.A(new_n1116), .B(KEYINPUT51), .Z(new_n1117));
  AOI211_X1 g0917(.A(new_n387), .B(new_n845), .C1(new_n1007), .C2(new_n839), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n832), .A2(G77), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1120), .B1(new_n201), .B2(new_n771), .C1(new_n203), .C2(new_n767), .ZN(new_n1121));
  OR3_X1    g0921(.A1(new_n1115), .A2(new_n1117), .A3(new_n1121), .ZN(new_n1122));
  OR2_X1    g0922(.A1(new_n1122), .A2(KEYINPUT110), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n782), .A2(new_n790), .B1(new_n996), .B2(new_n776), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT52), .ZN(new_n1125));
  INV_X1    g0925(.A(G322), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n387), .B1(new_n757), .B2(new_n1126), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n800), .B(new_n1127), .C1(G116), .C2(new_n832), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n564), .B2(new_n771), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(G283), .B2(new_n768), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1125), .B(new_n1130), .C1(new_n789), .C2(new_n754), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1122), .A2(KEYINPUT110), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1123), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1114), .B1(new_n1133), .B2(new_n805), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1134), .B1(new_n822), .B2(new_n1026), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n1110), .A2(new_n1111), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1111), .B1(new_n1110), .B2(new_n1135), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1109), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT112), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1109), .B(KEYINPUT112), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(G390));
  NAND3_X1  g0942(.A1(new_n729), .A2(G330), .A3(new_n863), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1143), .A2(new_n968), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n976), .A2(new_n979), .ZN(new_n1146));
  XOR2_X1   g0946(.A(new_n977), .B(KEYINPUT102), .Z(new_n1147));
  AOI21_X1  g0947(.A(new_n862), .B1(new_n745), .B2(new_n863), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1147), .B1(new_n1148), .B2(new_n968), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1146), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1147), .B1(new_n975), .B2(new_n903), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n734), .A2(new_n742), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n861), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1152), .A2(new_n695), .A3(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n968), .B1(new_n1154), .B2(new_n970), .ZN(new_n1155));
  NOR3_X1   g0955(.A1(new_n1151), .A2(new_n1155), .A3(KEYINPUT113), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT113), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n978), .B1(new_n962), .B2(new_n923), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n684), .B(new_n861), .C1(new_n734), .C2(new_n742), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n936), .B1(new_n1159), .B2(new_n862), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1157), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1145), .B(new_n1150), .C1(new_n1156), .C2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(KEYINPUT113), .B1(new_n1151), .B2(new_n1155), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1158), .A2(new_n1160), .A3(new_n1157), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n1163), .A2(new_n1164), .B1(new_n1146), .B2(new_n1149), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n935), .A2(new_n933), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n864), .B1(new_n1166), .B2(new_n931), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n941), .A2(new_n726), .A3(new_n942), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1167), .B(G330), .C1(new_n1168), .C2(new_n938), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1162), .B(new_n809), .C1(new_n1165), .C2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(KEYINPUT115), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n1150), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1169), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT115), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1175), .A2(new_n1176), .A3(new_n809), .A4(new_n1162), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1171), .A2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1162), .B1(new_n1165), .B2(new_n1169), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1148), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1143), .A2(KEYINPUT114), .A3(new_n968), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n1169), .ZN(new_n1182));
  AOI21_X1  g0982(.A(KEYINPUT114), .B1(new_n1143), .B2(new_n968), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1180), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(G330), .B1(new_n1168), .B2(new_n938), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n968), .B1(new_n1185), .B2(new_n864), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1159), .A2(new_n862), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1186), .A2(new_n1145), .A3(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1184), .A2(new_n1188), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n984), .B(new_n633), .C1(new_n446), .C2(new_n1185), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1179), .A2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1190), .B1(new_n1184), .B2(new_n1188), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1175), .A2(new_n1162), .A3(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1193), .A2(new_n1195), .A3(new_n709), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(KEYINPUT54), .B(G143), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n789), .A2(new_n1197), .B1(new_n836), .B2(new_n771), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n1198), .A2(KEYINPUT116), .B1(G159), .B2(new_n832), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(KEYINPUT116), .B2(new_n1198), .ZN(new_n1200));
  XOR2_X1   g1000(.A(new_n1200), .B(KEYINPUT117), .Z(new_n1201));
  NOR2_X1   g1001(.A1(new_n767), .A2(new_n837), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1202), .B(KEYINPUT53), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n291), .B1(new_n751), .B2(new_n201), .ZN(new_n1204));
  INV_X1    g1004(.A(G128), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n776), .A2(new_n1205), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1204), .B(new_n1206), .C1(new_n846), .C2(G125), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1203), .B(new_n1207), .C1(new_n834), .C2(new_n782), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1201), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT118), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n760), .A2(new_n754), .B1(new_n203), .B2(new_n751), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT119), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n795), .A2(new_n387), .A3(new_n1119), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n230), .A2(new_n771), .B1(new_n776), .B2(new_n848), .ZN(new_n1215));
  NOR3_X1   g1015(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1216), .B1(new_n569), .B2(new_n782), .C1(new_n789), .C2(new_n529), .ZN(new_n1217));
  OAI21_X1  g1017(.A(KEYINPUT118), .B1(new_n1201), .B2(new_n1208), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1211), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n805), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1146), .A2(new_n817), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n811), .B1(new_n379), .B2(new_n828), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1178), .A2(new_n1196), .A3(new_n1223), .ZN(G378));
  NOR2_X1   g1024(.A1(new_n291), .A2(G41), .ZN(new_n1225));
  AOI211_X1 g1025(.A(G50), .B(new_n1225), .C1(new_n383), .C2(new_n285), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n1006), .A2(new_n1225), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1227), .B1(new_n202), .B2(new_n751), .C1(new_n848), .C2(new_n760), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n768), .A2(G77), .B1(G97), .B2(new_n772), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n569), .B2(new_n776), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n1228), .B(new_n1230), .C1(G107), .C2(new_n783), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n789), .B2(new_n311), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1226), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  AOI211_X1 g1034(.A(G33), .B(G41), .C1(new_n1007), .C2(G124), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n796), .B2(new_n751), .ZN(new_n1236));
  XOR2_X1   g1036(.A(new_n1236), .B(KEYINPUT121), .Z(new_n1237));
  NOR2_X1   g1037(.A1(new_n782), .A2(new_n1205), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n772), .A2(G132), .B1(G150), .B2(new_n832), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1003), .A2(G125), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1239), .B(new_n1240), .C1(new_n767), .C2(new_n1197), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n1238), .B(new_n1241), .C1(new_n788), .C2(G137), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT59), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1237), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1242), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1245), .A2(KEYINPUT59), .ZN(new_n1246));
  OAI221_X1 g1046(.A(new_n1234), .B1(new_n1233), .B2(new_n1232), .C1(new_n1244), .C2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n805), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n811), .B1(new_n201), .B2(new_n828), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n630), .A2(new_n334), .A3(new_n631), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n682), .A2(new_n272), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1252), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n630), .A2(new_n334), .A3(new_n631), .A4(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1250), .B1(new_n1253), .B2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1253), .A2(new_n1255), .A3(new_n1250), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1248), .B(new_n1249), .C1(new_n1259), .C2(new_n818), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n982), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n925), .A2(new_n944), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n946), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n882), .B1(new_n963), .B2(new_n944), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1259), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(KEYINPUT40), .B1(new_n975), .B2(new_n903), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1167), .B1(new_n1168), .B2(new_n938), .ZN(new_n1268));
  OAI21_X1  g1068(.A(G330), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1253), .A2(new_n1255), .A3(new_n1250), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1270), .A2(new_n1256), .ZN(new_n1271));
  NOR3_X1   g1071(.A1(new_n945), .A2(new_n1269), .A3(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1262), .B1(new_n1266), .B2(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1271), .B1(new_n945), .B2(new_n1269), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1268), .B1(new_n905), .B2(new_n924), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1265), .B(new_n1259), .C1(new_n1275), .C2(KEYINPUT40), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1274), .A2(new_n1276), .A3(new_n982), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1273), .A2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1261), .B1(new_n1278), .B2(new_n809), .ZN(new_n1279));
  AOI221_X4 g1079(.A(new_n1144), .B1(new_n1146), .B2(new_n1149), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1169), .B1(new_n1172), .B2(new_n1150), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1190), .B1(new_n1282), .B2(new_n1189), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1274), .A2(new_n1276), .A3(new_n982), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n982), .B1(new_n1274), .B2(new_n1276), .ZN(new_n1285));
  OAI21_X1  g1085(.A(KEYINPUT57), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n709), .B1(new_n1283), .B2(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1191), .B1(new_n1179), .B2(new_n1192), .ZN(new_n1288));
  AOI21_X1  g1088(.A(KEYINPUT57), .B1(new_n1288), .B2(new_n1278), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1279), .B1(new_n1287), .B2(new_n1289), .ZN(G375));
  NAND3_X1  g1090(.A1(new_n1184), .A2(new_n1190), .A3(new_n1188), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1192), .A2(new_n1046), .A3(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n968), .A2(new_n817), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n291), .B1(new_n751), .B2(new_n202), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1294), .B1(G50), .B2(new_n832), .ZN(new_n1295));
  OAI221_X1 g1095(.A(new_n1295), .B1(new_n767), .B2(new_n392), .C1(new_n1205), .C2(new_n760), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1296), .B1(new_n788), .B2(G150), .ZN(new_n1297));
  XOR2_X1   g1097(.A(new_n1297), .B(KEYINPUT122), .Z(new_n1298));
  OAI22_X1  g1098(.A1(new_n834), .A2(new_n776), .B1(new_n771), .B2(new_n1197), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1299), .B1(new_n783), .B2(G137), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n291), .B1(new_n752), .B2(G77), .ZN(new_n1302));
  OAI221_X1 g1102(.A(new_n1302), .B1(new_n311), .B2(new_n756), .C1(new_n760), .C2(new_n564), .ZN(new_n1303));
  AOI22_X1  g1103(.A1(new_n768), .A2(G97), .B1(G116), .B2(new_n772), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1304), .B1(new_n754), .B2(new_n776), .ZN(new_n1305));
  AOI211_X1 g1105(.A(new_n1303), .B(new_n1305), .C1(G283), .C2(new_n783), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1306), .B1(new_n789), .B2(new_n230), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n856), .B1(new_n1301), .B2(new_n1307), .ZN(new_n1308));
  AOI211_X1 g1108(.A(new_n811), .B(new_n1308), .C1(new_n203), .C2(new_n828), .ZN(new_n1309));
  AOI22_X1  g1109(.A1(new_n1189), .A2(new_n809), .B1(new_n1293), .B2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1292), .A2(new_n1310), .ZN(G381));
  OAI21_X1  g1111(.A(new_n809), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n1260), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1288), .A2(new_n1278), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT57), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1315), .B1(new_n1273), .B2(new_n1277), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n710), .B1(new_n1317), .B2(new_n1288), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1313), .B1(new_n1316), .B2(new_n1318), .ZN(new_n1319));
  AND3_X1   g1119(.A1(new_n1178), .A2(new_n1196), .A3(new_n1223), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1101), .A2(new_n1105), .A3(new_n826), .A4(new_n823), .ZN(new_n1322));
  OR3_X1    g1122(.A1(new_n1322), .A2(G384), .A3(G381), .ZN(new_n1323));
  NOR3_X1   g1123(.A1(new_n1323), .A2(G390), .A3(G387), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1321), .B1(new_n1324), .B2(KEYINPUT123), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1325), .B1(KEYINPUT123), .B2(new_n1324), .ZN(G407));
  NAND2_X1  g1126(.A1(new_n683), .A2(G213), .ZN(new_n1327));
  XNOR2_X1  g1127(.A(new_n1327), .B(KEYINPUT124), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1328), .ZN(new_n1329));
  OAI211_X1 g1129(.A(G407), .B(G213), .C1(new_n1321), .C2(new_n1329), .ZN(G409));
  AOI21_X1  g1130(.A(new_n710), .B1(new_n1179), .B2(new_n1192), .ZN(new_n1331));
  AND2_X1   g1131(.A1(new_n1220), .A2(new_n1222), .ZN(new_n1332));
  AOI22_X1  g1132(.A1(new_n1195), .A2(new_n1331), .B1(new_n1332), .B2(new_n1221), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1288), .A2(new_n1046), .A3(new_n1278), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1333), .A2(new_n1178), .A3(new_n1279), .A4(new_n1334), .ZN(new_n1335));
  OAI211_X1 g1135(.A(new_n1329), .B(new_n1335), .C1(new_n1319), .C2(new_n1320), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT60), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1291), .A2(new_n1337), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1184), .A2(new_n1190), .A3(new_n1188), .A4(KEYINPUT60), .ZN(new_n1339));
  NAND4_X1  g1139(.A1(new_n1338), .A2(new_n1192), .A3(new_n709), .A4(new_n1339), .ZN(new_n1340));
  AND3_X1   g1140(.A1(new_n1340), .A2(G384), .A3(new_n1310), .ZN(new_n1341));
  AOI21_X1  g1141(.A(G384), .B1(new_n1340), .B2(new_n1310), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1343), .ZN(new_n1344));
  OAI21_X1  g1144(.A(KEYINPUT62), .B1(new_n1336), .B2(new_n1344), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT125), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1328), .A2(G2897), .ZN(new_n1347));
  INV_X1    g1147(.A(new_n1347), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1344), .A2(new_n1346), .A3(new_n1348), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1346), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1350));
  NOR3_X1   g1150(.A1(new_n1341), .A2(new_n1342), .A3(new_n1346), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1350), .B1(new_n1351), .B2(new_n1347), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1336), .A2(new_n1349), .A3(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT61), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(G375), .A2(G378), .ZN(new_n1355));
  AND2_X1   g1155(.A1(new_n1334), .A2(new_n1279), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1328), .B1(new_n1356), .B2(new_n1320), .ZN(new_n1357));
  INV_X1    g1157(.A(KEYINPUT62), .ZN(new_n1358));
  NAND4_X1  g1158(.A1(new_n1355), .A2(new_n1357), .A3(new_n1358), .A4(new_n1343), .ZN(new_n1359));
  NAND4_X1  g1159(.A1(new_n1345), .A2(new_n1353), .A3(new_n1354), .A4(new_n1359), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(G393), .A2(G396), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1361), .A2(new_n1322), .ZN(new_n1362));
  AOI21_X1  g1162(.A(G387), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1363));
  INV_X1    g1163(.A(KEYINPUT126), .ZN(new_n1364));
  OAI21_X1  g1164(.A(new_n1362), .B1(new_n1363), .B2(new_n1364), .ZN(new_n1365));
  INV_X1    g1165(.A(G387), .ZN(new_n1366));
  INV_X1    g1166(.A(new_n1137), .ZN(new_n1367));
  NAND3_X1  g1167(.A1(new_n1110), .A2(new_n1111), .A3(new_n1135), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1367), .A2(new_n1368), .ZN(new_n1369));
  AOI21_X1  g1169(.A(KEYINPUT112), .B1(new_n1369), .B2(new_n1109), .ZN(new_n1370));
  INV_X1    g1170(.A(new_n1141), .ZN(new_n1371));
  OAI21_X1  g1171(.A(new_n1366), .B1(new_n1370), .B2(new_n1371), .ZN(new_n1372));
  NAND3_X1  g1172(.A1(new_n1140), .A2(G387), .A3(new_n1141), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1372), .A2(new_n1373), .ZN(new_n1374));
  AND2_X1   g1174(.A1(new_n1365), .A2(new_n1374), .ZN(new_n1375));
  NAND4_X1  g1175(.A1(new_n1372), .A2(new_n1364), .A3(new_n1373), .A4(new_n1362), .ZN(new_n1376));
  INV_X1    g1176(.A(new_n1376), .ZN(new_n1377));
  NOR2_X1   g1177(.A1(new_n1375), .A2(new_n1377), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1360), .A2(new_n1378), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(new_n1316), .A2(new_n1318), .ZN(new_n1380));
  AOI21_X1  g1180(.A(new_n1320), .B1(new_n1380), .B2(new_n1279), .ZN(new_n1381));
  NAND2_X1  g1181(.A1(new_n1334), .A2(new_n1279), .ZN(new_n1382));
  OAI21_X1  g1182(.A(new_n1329), .B1(new_n1382), .B2(G378), .ZN(new_n1383));
  NOR3_X1   g1183(.A1(new_n1381), .A2(new_n1344), .A3(new_n1383), .ZN(new_n1384));
  NAND2_X1  g1184(.A1(new_n1365), .A2(new_n1374), .ZN(new_n1385));
  AOI22_X1  g1185(.A1(new_n1384), .A2(KEYINPUT63), .B1(new_n1385), .B2(new_n1376), .ZN(new_n1386));
  NAND2_X1  g1186(.A1(new_n1340), .A2(new_n1310), .ZN(new_n1387));
  INV_X1    g1187(.A(G384), .ZN(new_n1388));
  NAND2_X1  g1188(.A1(new_n1387), .A2(new_n1388), .ZN(new_n1389));
  NAND3_X1  g1189(.A1(new_n1340), .A2(G384), .A3(new_n1310), .ZN(new_n1390));
  NAND3_X1  g1190(.A1(new_n1389), .A2(KEYINPUT125), .A3(new_n1390), .ZN(new_n1391));
  NAND2_X1  g1191(.A1(new_n1391), .A2(new_n1348), .ZN(new_n1392));
  AOI22_X1  g1192(.A1(new_n1355), .A2(new_n1357), .B1(new_n1392), .B2(new_n1350), .ZN(new_n1393));
  AOI21_X1  g1193(.A(KEYINPUT61), .B1(new_n1393), .B2(new_n1349), .ZN(new_n1394));
  INV_X1    g1194(.A(KEYINPUT63), .ZN(new_n1395));
  OAI21_X1  g1195(.A(new_n1395), .B1(new_n1336), .B2(new_n1344), .ZN(new_n1396));
  NAND3_X1  g1196(.A1(new_n1386), .A2(new_n1394), .A3(new_n1396), .ZN(new_n1397));
  NAND2_X1  g1197(.A1(new_n1379), .A2(new_n1397), .ZN(G405));
  INV_X1    g1198(.A(KEYINPUT127), .ZN(new_n1399));
  OAI21_X1  g1199(.A(new_n1399), .B1(new_n1375), .B2(new_n1377), .ZN(new_n1400));
  NAND3_X1  g1200(.A1(new_n1385), .A2(KEYINPUT127), .A3(new_n1376), .ZN(new_n1401));
  NAND3_X1  g1201(.A1(new_n1355), .A2(new_n1321), .A3(new_n1343), .ZN(new_n1402));
  NAND2_X1  g1202(.A1(new_n1355), .A2(new_n1321), .ZN(new_n1403));
  NAND2_X1  g1203(.A1(new_n1403), .A2(new_n1344), .ZN(new_n1404));
  NAND4_X1  g1204(.A1(new_n1400), .A2(new_n1401), .A3(new_n1402), .A4(new_n1404), .ZN(new_n1405));
  NAND2_X1  g1205(.A1(new_n1404), .A2(new_n1402), .ZN(new_n1406));
  AND3_X1   g1206(.A1(new_n1385), .A2(KEYINPUT127), .A3(new_n1376), .ZN(new_n1407));
  AOI21_X1  g1207(.A(KEYINPUT127), .B1(new_n1385), .B2(new_n1376), .ZN(new_n1408));
  OAI21_X1  g1208(.A(new_n1406), .B1(new_n1407), .B2(new_n1408), .ZN(new_n1409));
  NAND2_X1  g1209(.A1(new_n1405), .A2(new_n1409), .ZN(G402));
endmodule


