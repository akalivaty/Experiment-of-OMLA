//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 0 1 0 1 1 1 0 1 0 1 1 0 1 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 1 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 1 0 1 0 1 1 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:52 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1113, new_n1114, new_n1115,
    new_n1116, new_n1117, new_n1118, new_n1119, new_n1120, new_n1121,
    new_n1122, new_n1123, new_n1124, new_n1125, new_n1126, new_n1127,
    new_n1128, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1207, new_n1208, new_n1209;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n202), .A2(new_n203), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT65), .Z(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n209), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  INV_X1    g0022(.A(G87), .ZN(new_n223));
  INV_X1    g0023(.A(G250), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n221), .B1(new_n203), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n226));
  INV_X1    g0026(.A(G77), .ZN(new_n227));
  INV_X1    g0027(.A(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G107), .ZN(new_n229));
  INV_X1    g0029(.A(G264), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n226), .B1(new_n227), .B2(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n211), .B1(new_n225), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n214), .B(new_n220), .C1(KEYINPUT1), .C2(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT66), .ZN(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n247), .B(new_n248), .Z(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  OAI21_X1  g0050(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n251));
  INV_X1    g0051(.A(G274), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G1), .A3(G13), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n251), .ZN(new_n256));
  XOR2_X1   g0056(.A(new_n256), .B(KEYINPUT67), .Z(new_n257));
  AOI21_X1  g0057(.A(new_n253), .B1(new_n257), .B2(G226), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT3), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G1698), .ZN(new_n264));
  INV_X1    g0064(.A(G223), .ZN(new_n265));
  OAI22_X1  g0065(.A1(new_n264), .A2(new_n265), .B1(new_n227), .B2(new_n263), .ZN(new_n266));
  AND2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(G1698), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n266), .B1(G222), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n258), .B1(new_n255), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G190), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n275), .A2(G50), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n210), .A2(G33), .B1(G1), .B2(G13), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT8), .B(G58), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n209), .A2(G33), .ZN(new_n279));
  OR2_X1    g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G20), .A2(G33), .ZN(new_n281));
  AOI22_X1  g0081(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n277), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n218), .B1(new_n211), .B2(new_n260), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n209), .A2(G1), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI211_X1 g0086(.A(new_n276), .B(new_n283), .C1(G50), .C2(new_n286), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n287), .A2(KEYINPUT9), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n287), .A2(KEYINPUT9), .ZN(new_n289));
  NOR4_X1   g0089(.A1(new_n274), .A2(new_n288), .A3(new_n289), .A4(KEYINPUT72), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT71), .B(G200), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n272), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT73), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  OR2_X1    g0094(.A1(new_n294), .A2(KEYINPUT10), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(KEYINPUT10), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n272), .A2(G179), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n297), .B(KEYINPUT68), .ZN(new_n298));
  INV_X1    g0098(.A(G169), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n287), .B1(new_n272), .B2(new_n299), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n295), .A2(new_n296), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  NOR3_X1   g0101(.A1(new_n201), .A2(G20), .A3(G33), .ZN(new_n302));
  OAI22_X1  g0102(.A1(new_n279), .A2(new_n227), .B1(new_n209), .B2(G68), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n284), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT11), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n305), .ZN(new_n307));
  OAI21_X1  g0107(.A(KEYINPUT12), .B1(new_n275), .B2(G68), .ZN(new_n308));
  OR3_X1    g0108(.A1(new_n275), .A2(KEYINPUT12), .A3(G68), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n286), .A2(G68), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AND3_X1   g0110(.A1(new_n306), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n270), .A2(G226), .ZN(new_n312));
  XNOR2_X1  g0112(.A(new_n312), .B(KEYINPUT74), .ZN(new_n313));
  INV_X1    g0113(.A(G97), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n260), .A2(new_n314), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n263), .A2(G232), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n315), .B1(new_n316), .B2(G1698), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n255), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n253), .B1(new_n257), .B2(G238), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT13), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT13), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n320), .A2(new_n324), .A3(new_n321), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n311), .B1(new_n326), .B2(new_n273), .ZN(new_n327));
  INV_X1    g0127(.A(G200), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n328), .B1(new_n323), .B2(new_n325), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n326), .A2(G169), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT75), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT14), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n323), .A2(G179), .A3(new_n325), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n332), .A2(new_n333), .ZN(new_n337));
  AND2_X1   g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n326), .B(G169), .C1(new_n332), .C2(new_n333), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n335), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  XNOR2_X1  g0140(.A(new_n311), .B(KEYINPUT76), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n330), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT69), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n257), .A2(G244), .ZN(new_n344));
  INV_X1    g0144(.A(G1698), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n263), .A2(G232), .A3(new_n345), .ZN(new_n346));
  OAI221_X1 g0146(.A(new_n346), .B1(new_n229), .B2(new_n263), .C1(new_n264), .C2(new_n222), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n319), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n208), .B(G274), .C1(G41), .C2(G45), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n344), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n343), .B1(new_n350), .B2(new_n291), .ZN(new_n351));
  INV_X1    g0151(.A(new_n350), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n351), .B1(G190), .B2(new_n352), .ZN(new_n353));
  NOR3_X1   g0153(.A1(new_n350), .A2(new_n343), .A3(new_n273), .ZN(new_n354));
  INV_X1    g0154(.A(new_n278), .ZN(new_n355));
  OR2_X1    g0155(.A1(new_n281), .A2(KEYINPUT70), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n281), .A2(KEYINPUT70), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  XNOR2_X1  g0158(.A(KEYINPUT15), .B(G87), .ZN(new_n359));
  OAI221_X1 g0159(.A(new_n358), .B1(new_n209), .B2(new_n227), .C1(new_n279), .C2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n284), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n286), .A2(G77), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n361), .B(new_n362), .C1(G77), .C2(new_n275), .ZN(new_n363));
  NOR3_X1   g0163(.A1(new_n353), .A2(new_n354), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G179), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n352), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n350), .A2(new_n299), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(new_n363), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n364), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n301), .A2(new_n342), .A3(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n261), .A2(new_n209), .A3(new_n262), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT7), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT7), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n261), .A2(new_n374), .A3(new_n209), .A4(new_n262), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n373), .A2(G68), .A3(new_n375), .ZN(new_n376));
  XNOR2_X1  g0176(.A(G58), .B(G68), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n377), .A2(G20), .B1(G159), .B2(new_n281), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT77), .ZN(new_n380));
  AOI21_X1  g0180(.A(KEYINPUT16), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n376), .B(new_n378), .C1(new_n380), .C2(KEYINPUT16), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n382), .A2(new_n284), .A3(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n355), .B1(new_n284), .B2(new_n285), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n278), .A2(new_n275), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n265), .A2(new_n345), .ZN(new_n389));
  INV_X1    g0189(.A(G226), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(G1698), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n389), .B(new_n391), .C1(new_n267), .C2(new_n268), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G33), .A2(G87), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n319), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n255), .A2(G232), .A3(new_n251), .ZN(new_n396));
  AND2_X1   g0196(.A1(new_n396), .A2(new_n349), .ZN(new_n397));
  AOI21_X1  g0197(.A(G169), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n255), .B1(new_n392), .B2(new_n393), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n396), .A2(new_n349), .ZN(new_n400));
  NOR3_X1   g0200(.A1(new_n399), .A2(new_n400), .A3(G179), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT78), .B1(new_n398), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n395), .A2(new_n365), .A3(new_n397), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT78), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n299), .B1(new_n399), .B2(new_n400), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n402), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT18), .ZN(new_n408));
  AND3_X1   g0208(.A1(new_n388), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n408), .B1(new_n388), .B2(new_n407), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT79), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n399), .A2(new_n400), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n273), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(G200), .B2(new_n412), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n384), .A2(new_n414), .A3(new_n387), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT80), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT17), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g0219(.A1(KEYINPUT80), .A2(KEYINPUT17), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n387), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n277), .B1(new_n379), .B2(new_n381), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n422), .B1(new_n423), .B2(new_n383), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n421), .B1(new_n424), .B2(new_n414), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT81), .B1(new_n419), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n415), .B1(new_n420), .B2(new_n418), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT81), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n424), .B(new_n414), .C1(new_n416), .C2(new_n417), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n404), .B1(new_n403), .B2(new_n405), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT18), .B1(new_n433), .B2(new_n424), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT79), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n388), .A2(new_n407), .A3(new_n408), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n411), .A2(new_n426), .A3(new_n430), .A4(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n371), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g0239(.A(KEYINPUT5), .B(G41), .ZN(new_n440));
  INV_X1    g0240(.A(G45), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n441), .A2(G1), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NOR3_X1   g0243(.A1(new_n443), .A2(new_n252), .A3(new_n319), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n319), .B1(new_n442), .B2(new_n440), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(G270), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n270), .A2(G257), .B1(G303), .B2(new_n269), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n449), .B1(new_n230), .B2(new_n264), .ZN(new_n450));
  OR2_X1    g0250(.A1(new_n450), .A2(KEYINPUT89), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n255), .B1(new_n450), .B2(KEYINPUT89), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n448), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G33), .A2(G283), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n454), .B(new_n209), .C1(G33), .C2(new_n314), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n284), .B(new_n455), .C1(new_n209), .C2(G116), .ZN(new_n456));
  XNOR2_X1  g0256(.A(new_n456), .B(KEYINPUT20), .ZN(new_n457));
  INV_X1    g0257(.A(new_n275), .ZN(new_n458));
  INV_X1    g0258(.A(G116), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n277), .B(new_n275), .C1(G1), .C2(new_n260), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n460), .B1(new_n461), .B2(new_n459), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n457), .A2(new_n462), .ZN(new_n463));
  NOR3_X1   g0263(.A1(new_n453), .A2(new_n463), .A3(new_n299), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT21), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT21), .ZN(new_n466));
  OR2_X1    g0266(.A1(new_n457), .A2(new_n462), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(G169), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n466), .B1(new_n468), .B2(new_n453), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n453), .A2(new_n467), .A3(G179), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n465), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n463), .B1(new_n453), .B2(new_n328), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n472), .B1(G190), .B2(new_n453), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n263), .A2(new_n209), .A3(G87), .ZN(new_n475));
  XNOR2_X1  g0275(.A(new_n475), .B(KEYINPUT22), .ZN(new_n476));
  NOR3_X1   g0276(.A1(new_n260), .A2(new_n459), .A3(G20), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT23), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n478), .B1(new_n209), .B2(G107), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n229), .A2(KEYINPUT23), .A3(G20), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g0282(.A(new_n482), .B(KEYINPUT24), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n284), .ZN(new_n484));
  INV_X1    g0284(.A(new_n461), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT25), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n486), .B1(new_n275), .B2(G107), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n458), .A2(KEYINPUT25), .A3(new_n229), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n485), .A2(G107), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n269), .A2(new_n345), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n491), .A2(G257), .B1(G33), .B2(G294), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n263), .A2(new_n345), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n492), .B1(new_n224), .B2(new_n493), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n494), .A2(new_n319), .B1(G264), .B2(new_n446), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n445), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G200), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n495), .A2(G190), .A3(new_n445), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(KEYINPUT90), .B1(new_n490), .B2(new_n499), .ZN(new_n500));
  AND2_X1   g0300(.A1(new_n497), .A2(new_n498), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT90), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n501), .A2(new_n502), .A3(new_n484), .A4(new_n489), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n496), .A2(new_n299), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n495), .A2(new_n365), .A3(new_n445), .ZN(new_n505));
  AND2_X1   g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n500), .A2(new_n503), .B1(new_n490), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n359), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n508), .A2(new_n275), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n263), .A2(new_n209), .A3(G68), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n279), .A2(new_n314), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n511), .B1(KEYINPUT19), .B2(new_n512), .ZN(new_n513));
  XOR2_X1   g0313(.A(KEYINPUT86), .B(G87), .Z(new_n514));
  NOR2_X1   g0314(.A1(G97), .A2(G107), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g0316(.A(new_n516), .B(KEYINPUT87), .ZN(new_n517));
  AOI21_X1  g0317(.A(G20), .B1(new_n315), .B2(KEYINPUT19), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n513), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  OAI221_X1 g0320(.A(new_n510), .B1(new_n359), .B2(new_n461), .C1(new_n520), .C2(new_n277), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT85), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n522), .B1(new_n270), .B2(G238), .ZN(new_n523));
  NOR3_X1   g0323(.A1(new_n493), .A2(KEYINPUT85), .A3(new_n222), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI22_X1  g0325(.A1(new_n264), .A2(new_n228), .B1(new_n260), .B2(new_n459), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n319), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR3_X1   g0327(.A1(new_n319), .A2(new_n224), .A3(new_n442), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n528), .B1(G274), .B2(new_n442), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n299), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n521), .B(new_n531), .C1(G179), .C2(new_n530), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n527), .A2(G190), .A3(new_n529), .ZN(new_n533));
  XNOR2_X1  g0333(.A(new_n533), .B(KEYINPUT88), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n520), .A2(new_n277), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n535), .A2(new_n509), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n530), .A2(new_n291), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n485), .A2(G87), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n532), .B1(new_n534), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n515), .A2(KEYINPUT6), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(KEYINPUT6), .B2(new_n314), .ZN(new_n542));
  XNOR2_X1  g0342(.A(KEYINPUT82), .B(G107), .ZN(new_n543));
  XNOR2_X1  g0343(.A(new_n542), .B(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G20), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n281), .A2(G77), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(KEYINPUT83), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n373), .A2(G107), .A3(new_n375), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT83), .B1(new_n545), .B2(new_n546), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n284), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT4), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n493), .B2(new_n228), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n491), .A2(G250), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(new_n454), .A3(new_n554), .ZN(new_n555));
  NOR3_X1   g0355(.A1(new_n493), .A2(new_n552), .A3(new_n228), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n319), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n444), .B1(new_n446), .B2(G257), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(G190), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n458), .A2(G97), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n562), .B1(new_n461), .B2(G97), .ZN(new_n563));
  XNOR2_X1  g0363(.A(new_n563), .B(KEYINPUT84), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n559), .A2(G200), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n551), .A2(new_n561), .A3(new_n564), .A4(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n559), .A2(new_n299), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(G179), .B2(new_n559), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n569), .B1(new_n551), .B2(new_n564), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n540), .A2(new_n567), .A3(new_n570), .ZN(new_n571));
  AND4_X1   g0371(.A1(new_n439), .A2(new_n474), .A3(new_n507), .A4(new_n571), .ZN(G372));
  NAND2_X1  g0372(.A1(new_n426), .A2(new_n430), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n340), .A2(new_n341), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n369), .B1(new_n327), .B2(new_n329), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n409), .A2(new_n410), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  OR2_X1    g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n295), .A2(new_n296), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n579), .A2(new_n580), .B1(new_n298), .B2(new_n300), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n551), .A2(new_n564), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n582), .B(new_n568), .C1(G179), .C2(new_n559), .ZN(new_n583));
  OAI21_X1  g0383(.A(KEYINPUT26), .B1(new_n540), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT26), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n536), .A2(new_n537), .A3(new_n538), .A4(new_n533), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n570), .A2(new_n585), .A3(new_n532), .A4(new_n586), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n584), .A2(new_n587), .A3(new_n532), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n532), .A2(new_n586), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n589), .B1(new_n500), .B2(new_n503), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n567), .A2(new_n570), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n490), .A2(new_n504), .A3(new_n505), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n592), .A2(new_n469), .A3(new_n465), .A4(new_n470), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n590), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n588), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n439), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n581), .A2(new_n596), .ZN(G369));
  NAND3_X1  g0397(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n598));
  OR2_X1    g0398(.A1(new_n598), .A2(KEYINPUT27), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(KEYINPUT27), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n599), .A2(G213), .A3(new_n600), .ZN(new_n601));
  XOR2_X1   g0401(.A(new_n601), .B(KEYINPUT91), .Z(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT92), .ZN(new_n604));
  OR2_X1    g0404(.A1(new_n604), .A2(G343), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(G343), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n603), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n608), .A2(new_n463), .ZN(new_n609));
  MUX2_X1   g0409(.A(new_n474), .B(new_n471), .S(new_n609), .Z(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(G330), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n490), .A2(new_n607), .ZN(new_n612));
  XOR2_X1   g0412(.A(new_n612), .B(KEYINPUT93), .Z(new_n613));
  AND2_X1   g0413(.A1(new_n500), .A2(new_n503), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n592), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n592), .A2(new_n607), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n611), .A2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n471), .A2(new_n608), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n616), .B1(new_n615), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n620), .A2(new_n623), .ZN(G399));
  NOR2_X1   g0424(.A1(new_n517), .A2(G116), .ZN(new_n625));
  INV_X1    g0425(.A(new_n212), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n626), .A2(G41), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n625), .A2(G1), .A3(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT94), .ZN(new_n630));
  OAI22_X1  g0430(.A1(new_n629), .A2(new_n630), .B1(new_n216), .B2(new_n628), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n630), .B2(new_n629), .ZN(new_n632));
  XOR2_X1   g0432(.A(new_n632), .B(KEYINPUT28), .Z(new_n633));
  INV_X1    g0433(.A(KEYINPUT31), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n474), .A2(new_n507), .A3(new_n571), .A4(new_n608), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT30), .ZN(new_n636));
  INV_X1    g0436(.A(new_n530), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n637), .A2(new_n495), .A3(new_n560), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n453), .A2(G179), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n636), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n496), .A2(new_n530), .A3(new_n365), .A4(new_n559), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n640), .B1(new_n453), .B2(new_n641), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n638), .A2(new_n639), .A3(new_n636), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n607), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n634), .B1(new_n635), .B2(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n644), .A2(new_n634), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(G330), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n540), .A2(new_n583), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n585), .ZN(new_n650));
  OAI21_X1  g0450(.A(KEYINPUT26), .B1(new_n583), .B2(new_n589), .ZN(new_n651));
  XOR2_X1   g0451(.A(new_n532), .B(KEYINPUT96), .Z(new_n652));
  NAND3_X1  g0452(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n590), .A2(new_n591), .A3(new_n593), .ZN(new_n654));
  OAI211_X1 g0454(.A(KEYINPUT29), .B(new_n608), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n607), .B1(new_n588), .B2(new_n594), .ZN(new_n656));
  XNOR2_X1  g0456(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n655), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n648), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n633), .B1(new_n660), .B2(G1), .ZN(G364));
  AND2_X1   g0461(.A1(new_n209), .A2(G13), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n208), .B1(new_n662), .B2(G45), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n627), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(G13), .A2(G33), .ZN(new_n667));
  XOR2_X1   g0467(.A(new_n667), .B(KEYINPUT97), .Z(new_n668));
  OR2_X1    g0468(.A1(new_n668), .A2(G20), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n669), .B(KEYINPUT98), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n218), .B1(G20), .B2(new_n299), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n217), .A2(new_n441), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n626), .A2(new_n263), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n674), .B(new_n675), .C1(new_n249), .C2(new_n441), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n626), .A2(new_n269), .ZN(new_n677));
  AOI22_X1  g0477(.A1(new_n677), .A2(G355), .B1(new_n459), .B2(new_n626), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n666), .B1(new_n673), .B2(new_n679), .ZN(new_n680));
  XOR2_X1   g0480(.A(new_n680), .B(KEYINPUT99), .Z(new_n681));
  NOR2_X1   g0481(.A1(new_n209), .A2(G190), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n365), .A2(G200), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(G179), .A2(G200), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(G159), .ZN(new_n688));
  OAI221_X1 g0488(.A(new_n263), .B1(new_n227), .B2(new_n684), .C1(new_n688), .C2(KEYINPUT32), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n689), .B1(KEYINPUT32), .B2(new_n688), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n291), .A2(new_n365), .A3(new_n682), .ZN(new_n691));
  XOR2_X1   g0491(.A(new_n691), .B(KEYINPUT100), .Z(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G107), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n209), .B1(new_n685), .B2(G190), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n694), .A2(KEYINPUT101), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(KEYINPUT101), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G97), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n209), .A2(new_n273), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n683), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n365), .A2(new_n328), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n682), .ZN(new_n703));
  OAI22_X1  g0503(.A1(new_n202), .A2(new_n701), .B1(new_n703), .B2(new_n203), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n291), .A2(new_n365), .A3(new_n700), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(new_n514), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n700), .A2(new_n702), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  AOI211_X1 g0508(.A(new_n704), .B(new_n706), .C1(G50), .C2(new_n708), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n690), .A2(new_n693), .A3(new_n699), .A4(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(G303), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n705), .A2(new_n711), .ZN(new_n712));
  XOR2_X1   g0512(.A(KEYINPUT33), .B(G317), .Z(new_n713));
  INV_X1    g0513(.A(G329), .ZN(new_n714));
  OAI22_X1  g0514(.A1(new_n713), .A2(new_n703), .B1(new_n686), .B2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(G326), .ZN(new_n716));
  INV_X1    g0516(.A(G311), .ZN(new_n717));
  OAI22_X1  g0517(.A1(new_n707), .A2(new_n716), .B1(new_n684), .B2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(G322), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n269), .B1(new_n701), .B2(new_n719), .ZN(new_n720));
  NOR4_X1   g0520(.A1(new_n712), .A2(new_n715), .A3(new_n718), .A4(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(G294), .ZN(new_n722));
  INV_X1    g0522(.A(new_n692), .ZN(new_n723));
  INV_X1    g0523(.A(G283), .ZN(new_n724));
  OAI221_X1 g0524(.A(new_n721), .B1(new_n722), .B2(new_n697), .C1(new_n723), .C2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n710), .A2(new_n725), .A3(KEYINPUT102), .ZN(new_n726));
  AOI21_X1  g0526(.A(KEYINPUT102), .B1(new_n710), .B2(new_n725), .ZN(new_n727));
  INV_X1    g0527(.A(new_n672), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n681), .B1(new_n726), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(new_n610), .B2(new_n670), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n611), .A2(new_n666), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n610), .A2(G330), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n731), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n734), .B(KEYINPUT103), .ZN(G396));
  INV_X1    g0535(.A(new_n701), .ZN(new_n736));
  AOI22_X1  g0536(.A1(G294), .A2(new_n736), .B1(new_n687), .B2(G311), .ZN(new_n737));
  OAI221_X1 g0537(.A(new_n737), .B1(new_n459), .B2(new_n684), .C1(new_n711), .C2(new_n707), .ZN(new_n738));
  INV_X1    g0538(.A(new_n703), .ZN(new_n739));
  AOI211_X1 g0539(.A(new_n263), .B(new_n738), .C1(G283), .C2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n692), .A2(G87), .ZN(new_n741));
  INV_X1    g0541(.A(new_n705), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G107), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n740), .A2(new_n699), .A3(new_n741), .A4(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n684), .ZN(new_n745));
  AOI22_X1  g0545(.A1(G143), .A2(new_n736), .B1(new_n745), .B2(G159), .ZN(new_n746));
  INV_X1    g0546(.A(G137), .ZN(new_n747));
  INV_X1    g0547(.A(G150), .ZN(new_n748));
  OAI221_X1 g0548(.A(new_n746), .B1(new_n747), .B2(new_n707), .C1(new_n748), .C2(new_n703), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT34), .ZN(new_n750));
  INV_X1    g0550(.A(G132), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n263), .B1(new_n686), .B2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n752), .B1(new_n742), .B2(G50), .ZN(new_n753));
  OAI211_X1 g0553(.A(new_n750), .B(new_n753), .C1(new_n202), .C2(new_n697), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n723), .A2(new_n203), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n744), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(new_n672), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n672), .A2(new_n667), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n666), .B1(new_n227), .B2(new_n758), .ZN(new_n759));
  AND2_X1   g0559(.A1(new_n607), .A2(new_n363), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n368), .B1(new_n364), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n369), .A2(new_n608), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n757), .B(new_n759), .C1(new_n764), .C2(new_n668), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n656), .B(new_n763), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n665), .B1(new_n767), .B2(new_n648), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n767), .A2(new_n648), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n765), .B1(new_n769), .B2(new_n770), .ZN(G384));
  INV_X1    g0571(.A(new_n544), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT35), .ZN(new_n773));
  OAI211_X1 g0573(.A(G116), .B(new_n219), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n774), .B1(new_n773), .B2(new_n772), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT36), .ZN(new_n776));
  INV_X1    g0576(.A(new_n216), .ZN(new_n777));
  OAI211_X1 g0577(.A(new_n777), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n201), .A2(G68), .ZN(new_n779));
  AOI211_X1 g0579(.A(new_n208), .B(G13), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n424), .A2(new_n603), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n434), .B(new_n436), .C1(new_n419), .C2(new_n425), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n415), .B1(new_n433), .B2(new_n424), .ZN(new_n784));
  OAI21_X1  g0584(.A(KEYINPUT37), .B1(new_n784), .B2(new_n782), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n388), .A2(new_n407), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n388), .A2(new_n602), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT37), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n786), .A2(new_n787), .A3(new_n788), .A4(new_n415), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n782), .A2(new_n783), .B1(new_n785), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(KEYINPUT107), .B1(new_n790), .B2(KEYINPUT38), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT104), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT16), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n277), .B1(new_n379), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n376), .A2(KEYINPUT16), .A3(new_n378), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n422), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n415), .B1(new_n603), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n433), .A2(new_n796), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n792), .B(KEYINPUT37), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n799), .A2(new_n789), .ZN(new_n800));
  OAI21_X1  g0600(.A(KEYINPUT37), .B1(new_n797), .B2(new_n798), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(KEYINPUT104), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n796), .A2(new_n603), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n800), .A2(new_n802), .B1(new_n438), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n791), .B1(new_n805), .B2(KEYINPUT38), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT107), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n438), .A2(new_n804), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n802), .A2(new_n799), .A3(new_n789), .ZN(new_n809));
  AND4_X1   g0609(.A1(new_n807), .A2(new_n808), .A3(KEYINPUT38), .A4(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n806), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n341), .A2(new_n607), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n342), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n341), .B(new_n607), .C1(new_n340), .C2(new_n330), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n763), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n647), .A2(KEYINPUT40), .A3(new_n811), .A4(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(KEYINPUT38), .B1(new_n808), .B2(new_n809), .ZN(new_n817));
  AND3_X1   g0617(.A1(new_n808), .A2(KEYINPUT38), .A3(new_n809), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT105), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n805), .A2(KEYINPUT38), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(KEYINPUT105), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n820), .A2(KEYINPUT106), .A3(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT106), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n808), .A2(new_n809), .A3(new_n819), .A4(KEYINPUT38), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(KEYINPUT38), .B2(new_n805), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n819), .B1(new_n805), .B2(KEYINPUT38), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n824), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n823), .A2(new_n828), .ZN(new_n829));
  AND3_X1   g0629(.A1(new_n829), .A2(new_n647), .A3(new_n815), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n816), .B1(new_n830), .B2(KEYINPUT40), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n647), .A2(new_n439), .ZN(new_n832));
  OR2_X1    g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n831), .A2(new_n832), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n833), .A2(G330), .A3(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n762), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(new_n656), .B2(new_n764), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n813), .A2(new_n814), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n840), .A2(new_n829), .B1(new_n578), .B2(new_n603), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT39), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(new_n820), .B2(new_n822), .ZN(new_n843));
  INV_X1    g0643(.A(new_n791), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n821), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n818), .A2(new_n807), .ZN(new_n846));
  AOI21_X1  g0646(.A(KEYINPUT39), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(KEYINPUT108), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n340), .A2(new_n341), .A3(new_n608), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(KEYINPUT39), .B1(new_n826), .B2(new_n827), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n842), .B1(new_n806), .B2(new_n810), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT108), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n848), .A2(new_n850), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n841), .A2(new_n855), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n439), .B(new_n655), .C1(new_n656), .C2(new_n658), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n581), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n856), .B(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n835), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n208), .B2(new_n662), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n835), .A2(new_n859), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n781), .B1(new_n861), .B2(new_n862), .ZN(G367));
  NAND3_X1  g0663(.A1(new_n615), .A2(new_n617), .A3(new_n622), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n582), .A2(new_n607), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n591), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n583), .B2(new_n608), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  OR2_X1    g0668(.A1(new_n864), .A2(new_n868), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n869), .A2(KEYINPUT42), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(KEYINPUT42), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n583), .B1(new_n866), .B2(new_n592), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n608), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n870), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n608), .B1(new_n536), .B2(new_n538), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n875), .B(KEYINPUT109), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n876), .A2(new_n532), .A3(new_n586), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n877), .B1(new_n532), .B2(new_n876), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT110), .ZN(new_n879));
  OR2_X1    g0679(.A1(new_n879), .A2(KEYINPUT43), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(KEYINPUT43), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n878), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(KEYINPUT43), .B2(new_n878), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n874), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n870), .A2(new_n871), .A3(new_n873), .A4(new_n882), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n620), .A2(new_n868), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n886), .B(new_n887), .ZN(new_n888));
  XOR2_X1   g0688(.A(new_n627), .B(KEYINPUT41), .Z(new_n889));
  NAND2_X1  g0689(.A1(new_n623), .A2(new_n867), .ZN(new_n890));
  XOR2_X1   g0690(.A(new_n890), .B(KEYINPUT45), .Z(new_n891));
  NOR2_X1   g0691(.A1(new_n623), .A2(new_n867), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n892), .B(KEYINPUT44), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n619), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n618), .A2(new_n621), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n896), .A2(new_n611), .A3(new_n864), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n611), .B1(new_n896), .B2(new_n864), .ZN(new_n898));
  OR2_X1    g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n660), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT111), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n899), .A2(new_n660), .A3(KEYINPUT111), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n891), .A2(new_n620), .A3(new_n893), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n895), .A2(new_n902), .A3(new_n903), .A4(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n889), .B1(new_n905), .B2(new_n660), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n888), .B1(new_n906), .B2(new_n664), .ZN(new_n907));
  INV_X1    g0707(.A(new_n673), .ZN(new_n908));
  INV_X1    g0708(.A(new_n675), .ZN(new_n909));
  OAI22_X1  g0709(.A1(new_n909), .A2(new_n241), .B1(new_n212), .B2(new_n359), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n665), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  AOI22_X1  g0711(.A1(G159), .A2(new_n739), .B1(new_n687), .B2(G137), .ZN(new_n912));
  OAI221_X1 g0712(.A(new_n912), .B1(new_n201), .B2(new_n684), .C1(new_n748), .C2(new_n701), .ZN(new_n913));
  AOI211_X1 g0713(.A(new_n269), .B(new_n913), .C1(G143), .C2(new_n708), .ZN(new_n914));
  OAI221_X1 g0714(.A(new_n914), .B1(new_n202), .B2(new_n705), .C1(new_n227), .C2(new_n691), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n697), .A2(new_n203), .ZN(new_n916));
  AOI22_X1  g0716(.A1(G294), .A2(new_n739), .B1(new_n736), .B2(G303), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n708), .A2(G311), .B1(new_n745), .B2(G283), .ZN(new_n918));
  INV_X1    g0718(.A(new_n691), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(G97), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n263), .B1(new_n687), .B2(G317), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n917), .A2(new_n918), .A3(new_n920), .A4(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n742), .A2(KEYINPUT46), .A3(G116), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT46), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n705), .B2(new_n459), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n923), .B(new_n925), .C1(new_n229), .C2(new_n697), .ZN(new_n926));
  OAI22_X1  g0726(.A1(new_n915), .A2(new_n916), .B1(new_n922), .B2(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT47), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n911), .B1(new_n928), .B2(new_n672), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n878), .B2(new_n670), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n907), .A2(new_n930), .ZN(G387));
  NAND2_X1  g0731(.A1(new_n902), .A2(new_n903), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n932), .B(new_n627), .C1(new_n660), .C2(new_n899), .ZN(new_n933));
  INV_X1    g0733(.A(new_n625), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n934), .A2(new_n677), .B1(new_n229), .B2(new_n626), .ZN(new_n935));
  AND3_X1   g0735(.A1(new_n355), .A2(KEYINPUT50), .A3(new_n201), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT50), .B1(new_n355), .B2(new_n201), .ZN(new_n937));
  OAI221_X1 g0737(.A(new_n441), .B1(new_n203), .B2(new_n227), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n675), .B1(new_n934), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n238), .A2(new_n441), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n935), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n908), .B1(new_n941), .B2(KEYINPUT112), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(KEYINPUT112), .B2(new_n941), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n698), .A2(new_n508), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n355), .A2(new_n739), .B1(new_n745), .B2(G68), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n708), .A2(G159), .B1(new_n687), .B2(G150), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n269), .B1(new_n736), .B2(G50), .ZN(new_n947));
  AND3_X1   g0747(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n944), .B(new_n948), .C1(new_n227), .C2(new_n705), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(G97), .B2(new_n692), .ZN(new_n950));
  AOI22_X1  g0750(.A1(G317), .A2(new_n736), .B1(new_n745), .B2(G303), .ZN(new_n951));
  OAI221_X1 g0751(.A(new_n951), .B1(new_n717), .B2(new_n703), .C1(new_n719), .C2(new_n707), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT48), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n953), .B1(new_n724), .B2(new_n697), .C1(new_n722), .C2(new_n705), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT49), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n269), .B1(new_n686), .B2(new_n716), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(new_n919), .B2(G116), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n950), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n665), .B(new_n943), .C1(new_n958), .C2(new_n728), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(new_n618), .B2(new_n671), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(new_n899), .B2(new_n664), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n933), .A2(new_n961), .ZN(G393));
  OAI21_X1  g0762(.A(new_n673), .B1(new_n314), .B2(new_n212), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n246), .A2(new_n675), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n665), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  AOI22_X1  g0765(.A1(G150), .A2(new_n708), .B1(new_n736), .B2(G159), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n966), .A2(KEYINPUT51), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n263), .B1(new_n703), .B2(new_n201), .ZN(new_n968));
  INV_X1    g0768(.A(G143), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n684), .A2(new_n278), .B1(new_n686), .B2(new_n969), .ZN(new_n970));
  NOR3_X1   g0770(.A1(new_n967), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n698), .A2(G77), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n966), .A2(KEYINPUT51), .B1(G68), .B2(new_n742), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n971), .A2(new_n741), .A3(new_n972), .A4(new_n973), .ZN(new_n974));
  AOI22_X1  g0774(.A1(G317), .A2(new_n708), .B1(new_n736), .B2(G311), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT52), .Z(new_n976));
  AOI21_X1  g0776(.A(new_n263), .B1(new_n745), .B2(G294), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n705), .A2(new_n724), .B1(new_n719), .B2(new_n686), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT113), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n976), .A2(new_n693), .A3(new_n977), .A4(new_n979), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n697), .A2(new_n459), .B1(new_n711), .B2(new_n703), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT114), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n974), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n965), .B1(new_n983), .B2(new_n672), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n867), .B2(new_n670), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n895), .A2(new_n904), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n985), .B1(new_n986), .B2(new_n663), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n905), .A2(new_n627), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(new_n932), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n987), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(G390));
  NAND3_X1  g0791(.A1(new_n647), .A2(G330), .A3(new_n439), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n581), .A2(new_n992), .A3(new_n857), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n647), .A2(G330), .A3(new_n815), .ZN(new_n994));
  OAI211_X1 g0794(.A(G330), .B(new_n764), .C1(new_n645), .C2(new_n646), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n839), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n584), .A2(new_n587), .A3(new_n532), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n608), .B(new_n764), .C1(new_n654), .C2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n762), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n608), .B(new_n761), .C1(new_n653), .C2(new_n654), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n994), .A2(new_n996), .A3(new_n762), .A4(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n993), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n994), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n850), .B1(new_n1000), .B2(new_n838), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(new_n848), .B2(new_n854), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n811), .A2(new_n849), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1002), .A2(new_n762), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1009), .B1(new_n838), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1006), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n849), .B1(new_n837), .B2(new_n839), .ZN(new_n1013));
  AND3_X1   g0813(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n853), .B1(new_n851), .B2(new_n852), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1013), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1011), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1016), .A2(new_n994), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1012), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1005), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1004), .A2(new_n1012), .A3(new_n1018), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1020), .A2(new_n627), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT117), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1012), .A2(new_n664), .A3(new_n1018), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT115), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1012), .A2(new_n1018), .A3(KEYINPUT115), .A4(new_n664), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n668), .B1(new_n848), .B2(new_n854), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n705), .A2(new_n748), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT53), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n698), .A2(G159), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n919), .A2(G50), .ZN(new_n1033));
  INV_X1    g0833(.A(G128), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n707), .A2(new_n1034), .B1(new_n701), .B2(new_n751), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(KEYINPUT54), .B(G143), .ZN(new_n1036));
  INV_X1    g0836(.A(G125), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n684), .A2(new_n1036), .B1(new_n686), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n263), .B1(new_n703), .B2(new_n747), .ZN(new_n1039));
  NOR3_X1   g0839(.A1(new_n1035), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .A4(new_n1040), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n703), .A2(new_n229), .B1(new_n686), .B2(new_n722), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n701), .A2(new_n459), .B1(new_n684), .B2(new_n314), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1042), .B(new_n1043), .C1(G283), .C2(new_n708), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n972), .B(new_n1044), .C1(new_n723), .C2(new_n203), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n269), .B1(new_n705), .B2(new_n223), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT116), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1041), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n672), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n758), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1049), .B(new_n665), .C1(new_n355), .C2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1029), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1023), .B1(new_n1028), .B2(new_n1053), .ZN(new_n1054));
  AOI211_X1 g0854(.A(KEYINPUT117), .B(new_n1052), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1022), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT118), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  OAI211_X1 g0858(.A(KEYINPUT118), .B(new_n1022), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n1058), .A2(new_n1059), .ZN(G378));
  INV_X1    g0860(.A(KEYINPUT120), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT57), .ZN(new_n1062));
  OAI211_X1 g0862(.A(G330), .B(new_n816), .C1(new_n830), .C2(KEYINPUT40), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n603), .A2(new_n287), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n301), .B(new_n1064), .Z(new_n1065));
  XNOR2_X1  g0865(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1065), .B(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1068), .A2(new_n841), .A3(new_n855), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1068), .B1(new_n855), .B2(new_n841), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1063), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1063), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1068), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n856), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1073), .A2(new_n1075), .A3(new_n1069), .ZN(new_n1076));
  AND2_X1   g0876(.A1(new_n1072), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n993), .ZN(new_n1078));
  AND2_X1   g0878(.A1(new_n1021), .A2(new_n1078), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1061), .B(new_n1062), .C1(new_n1077), .C2(new_n1079), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n1072), .A2(new_n1076), .B1(new_n1021), .B2(new_n1078), .ZN(new_n1081));
  OAI21_X1  g0881(.A(KEYINPUT120), .B1(new_n1081), .B2(KEYINPUT57), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n628), .B1(new_n1081), .B2(KEYINPUT57), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1080), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n663), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n665), .B1(G50), .B2(new_n1050), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1068), .A2(new_n668), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n916), .ZN(new_n1088));
  AOI211_X1 g0888(.A(G41), .B(new_n263), .C1(new_n736), .C2(G107), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n707), .A2(new_n459), .B1(new_n703), .B2(new_n314), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n684), .A2(new_n359), .B1(new_n686), .B2(new_n724), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(G58), .A2(new_n919), .B1(new_n742), .B2(G77), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1088), .A2(new_n1089), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT58), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n201), .B1(new_n267), .B2(G41), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n1034), .A2(new_n701), .B1(new_n703), .B2(new_n751), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n707), .A2(new_n1037), .B1(new_n684), .B2(new_n747), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n1099), .B1(new_n697), .B2(new_n748), .C1(new_n705), .C2(new_n1036), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1100), .A2(KEYINPUT59), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(KEYINPUT59), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n919), .A2(G159), .ZN(new_n1103));
  AOI211_X1 g0903(.A(G33), .B(G41), .C1(new_n687), .C2(G124), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1102), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1095), .B(new_n1096), .C1(new_n1101), .C2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT119), .ZN(new_n1107));
  OR2_X1    g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n728), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1086), .B(new_n1087), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1085), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1084), .A2(new_n1111), .ZN(G375));
  INV_X1    g0912(.A(new_n1001), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1003), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n993), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n889), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1116), .A2(new_n1117), .A3(new_n1005), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n839), .A2(new_n667), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT121), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n707), .A2(new_n751), .B1(new_n701), .B2(new_n747), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n703), .A2(new_n1036), .B1(new_n686), .B2(new_n1034), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n263), .B1(new_n684), .B2(new_n748), .ZN(new_n1123));
  NOR3_X1   g0923(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(G58), .A2(new_n919), .B1(new_n742), .B2(G159), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1124), .B(new_n1125), .C1(new_n201), .C2(new_n697), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n708), .A2(G294), .B1(new_n745), .B2(G107), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n1127), .B1(new_n459), .B2(new_n703), .C1(new_n724), .C2(new_n701), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n263), .B(new_n1128), .C1(G303), .C2(new_n687), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1129), .B(new_n944), .C1(new_n314), .C2(new_n705), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n723), .A2(new_n227), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1126), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n672), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n666), .B1(new_n203), .B2(new_n758), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1120), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n1115), .B2(new_n663), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1118), .A2(new_n1137), .ZN(G381));
  NOR2_X1   g0938(.A1(G375), .A2(new_n1056), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n990), .A2(new_n907), .A3(new_n930), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  NOR4_X1   g0941(.A1(G393), .A2(G381), .A3(G396), .A4(G384), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1139), .A2(new_n1141), .A3(new_n1142), .ZN(G407));
  NAND3_X1  g0943(.A1(new_n605), .A2(new_n606), .A3(G213), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n1139), .A2(KEYINPUT122), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(KEYINPUT122), .B1(new_n1139), .B2(new_n1145), .ZN(new_n1147));
  OAI211_X1 g0947(.A(G213), .B(G407), .C1(new_n1146), .C2(new_n1147), .ZN(G409));
  AOI21_X1  g0948(.A(new_n990), .B1(new_n907), .B2(new_n930), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT126), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1150), .A2(new_n1151), .A3(new_n1140), .ZN(new_n1152));
  OAI21_X1  g0952(.A(KEYINPUT126), .B1(new_n1141), .B2(new_n1149), .ZN(new_n1153));
  XOR2_X1   g0953(.A(G393), .B(G396), .Z(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1152), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1154), .B(KEYINPUT126), .C1(new_n1141), .C2(new_n1149), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1058), .A2(new_n1059), .A3(new_n1111), .A4(new_n1084), .ZN(new_n1159));
  OR3_X1    g0959(.A1(new_n1085), .A2(KEYINPUT123), .A3(new_n1110), .ZN(new_n1160));
  OAI21_X1  g0960(.A(KEYINPUT123), .B1(new_n1085), .B2(new_n1110), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1081), .A2(new_n1117), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1056), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1145), .B1(new_n1159), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT60), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1116), .B1(new_n1167), .B2(new_n1004), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1115), .A2(KEYINPUT60), .A3(new_n993), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1168), .A2(new_n627), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n1137), .ZN(new_n1171));
  INV_X1    g0971(.A(G384), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1170), .A2(G384), .A3(new_n1137), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n1176), .A2(KEYINPUT62), .ZN(new_n1177));
  AND2_X1   g0977(.A1(new_n1166), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1159), .A2(new_n1165), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(KEYINPUT124), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT124), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1159), .A2(new_n1181), .A3(new_n1165), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1180), .A2(new_n1144), .A3(new_n1176), .A4(new_n1182), .ZN(new_n1183));
  XOR2_X1   g0983(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1184));
  AOI21_X1  g0984(.A(new_n1178), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT61), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1145), .A2(G2897), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1175), .A2(KEYINPUT125), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT125), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1188), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n1188), .B2(new_n1191), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1186), .B1(new_n1193), .B2(new_n1166), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1158), .B1(new_n1185), .B2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1156), .A2(new_n1186), .A3(new_n1157), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT63), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1175), .A2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1196), .B1(new_n1166), .B2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1180), .A2(new_n1144), .A3(new_n1182), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1191), .A2(new_n1188), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1192), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1197), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1183), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1199), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1195), .A2(new_n1205), .ZN(G405));
  NAND2_X1  g1006(.A1(G375), .A2(new_n1164), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1159), .A2(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(new_n1176), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(new_n1158), .ZN(G402));
endmodule


