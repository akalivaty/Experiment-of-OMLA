

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589;

  NOR2_X1 U326 ( .A1(n568), .A2(n387), .ZN(n388) );
  INV_X1 U327 ( .A(KEYINPUT112), .ZN(n383) );
  XNOR2_X1 U328 ( .A(n370), .B(n369), .ZN(n372) );
  XNOR2_X1 U329 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U330 ( .A(n434), .B(n433), .ZN(n452) );
  XOR2_X1 U331 ( .A(n362), .B(n361), .Z(n294) );
  NOR2_X1 U332 ( .A1(n415), .A2(n519), .ZN(n575) );
  XNOR2_X1 U333 ( .A(G99GAT), .B(G85GAT), .ZN(n334) );
  XOR2_X1 U334 ( .A(n334), .B(G106GAT), .Z(n377) );
  XNOR2_X1 U335 ( .A(KEYINPUT48), .B(n391), .ZN(n548) );
  XOR2_X1 U336 ( .A(KEYINPUT36), .B(n568), .Z(n587) );
  XOR2_X1 U337 ( .A(n343), .B(n340), .Z(n580) );
  XNOR2_X1 U338 ( .A(n378), .B(n377), .ZN(n568) );
  XNOR2_X1 U339 ( .A(n457), .B(G183GAT), .ZN(n458) );
  XNOR2_X1 U340 ( .A(n459), .B(n458), .ZN(G1350GAT) );
  XOR2_X1 U341 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n296) );
  NAND2_X1 U342 ( .A1(G226GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U343 ( .A(n296), .B(n295), .ZN(n306) );
  XOR2_X1 U344 ( .A(KEYINPUT21), .B(KEYINPUT82), .Z(n298) );
  XNOR2_X1 U345 ( .A(G197GAT), .B(G218GAT), .ZN(n297) );
  XNOR2_X1 U346 ( .A(n298), .B(n297), .ZN(n420) );
  XOR2_X1 U347 ( .A(G204GAT), .B(G64GAT), .Z(n300) );
  XNOR2_X1 U348 ( .A(G176GAT), .B(G92GAT), .ZN(n299) );
  XNOR2_X1 U349 ( .A(n300), .B(n299), .ZN(n332) );
  XOR2_X1 U350 ( .A(n420), .B(n332), .Z(n304) );
  XNOR2_X1 U351 ( .A(G36GAT), .B(G190GAT), .ZN(n301) );
  XNOR2_X1 U352 ( .A(n301), .B(KEYINPUT74), .ZN(n367) );
  XNOR2_X1 U353 ( .A(G8GAT), .B(G183GAT), .ZN(n302) );
  XNOR2_X1 U354 ( .A(n302), .B(G211GAT), .ZN(n352) );
  XNOR2_X1 U355 ( .A(n367), .B(n352), .ZN(n303) );
  XNOR2_X1 U356 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U357 ( .A(n306), .B(n305), .ZN(n311) );
  XOR2_X1 U358 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n308) );
  XNOR2_X1 U359 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n307) );
  XNOR2_X1 U360 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U361 ( .A(KEYINPUT80), .B(n309), .ZN(n447) );
  INV_X1 U362 ( .A(n447), .ZN(n310) );
  XOR2_X1 U363 ( .A(n311), .B(n310), .Z(n523) );
  XNOR2_X1 U364 ( .A(KEYINPUT120), .B(n523), .ZN(n392) );
  XOR2_X1 U365 ( .A(G22GAT), .B(G15GAT), .Z(n341) );
  XOR2_X1 U366 ( .A(G197GAT), .B(G36GAT), .Z(n313) );
  XNOR2_X1 U367 ( .A(G29GAT), .B(G50GAT), .ZN(n312) );
  XNOR2_X1 U368 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U369 ( .A(n341), .B(n314), .Z(n316) );
  NAND2_X1 U370 ( .A1(G229GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U371 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U372 ( .A(n317), .B(KEYINPUT29), .Z(n320) );
  XNOR2_X1 U373 ( .A(G43GAT), .B(KEYINPUT7), .ZN(n318) );
  XNOR2_X1 U374 ( .A(n318), .B(KEYINPUT8), .ZN(n371) );
  XNOR2_X1 U375 ( .A(G169GAT), .B(n371), .ZN(n319) );
  XNOR2_X1 U376 ( .A(n320), .B(n319), .ZN(n328) );
  XOR2_X1 U377 ( .A(KEYINPUT67), .B(KEYINPUT68), .Z(n322) );
  XNOR2_X1 U378 ( .A(G1GAT), .B(G8GAT), .ZN(n321) );
  XNOR2_X1 U379 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U380 ( .A(KEYINPUT66), .B(G113GAT), .Z(n324) );
  XNOR2_X1 U381 ( .A(KEYINPUT30), .B(G141GAT), .ZN(n323) );
  XNOR2_X1 U382 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U383 ( .A(n326), .B(n325), .Z(n327) );
  XOR2_X1 U384 ( .A(n328), .B(n327), .Z(n551) );
  XOR2_X1 U385 ( .A(G71GAT), .B(KEYINPUT13), .Z(n329) );
  XOR2_X1 U386 ( .A(G78GAT), .B(n329), .Z(n343) );
  XOR2_X1 U387 ( .A(KEYINPUT69), .B(KEYINPUT32), .Z(n331) );
  NAND2_X1 U388 ( .A1(G230GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U389 ( .A(n331), .B(n330), .ZN(n333) );
  XOR2_X1 U390 ( .A(n333), .B(n332), .Z(n336) );
  XOR2_X1 U391 ( .A(n377), .B(G57GAT), .Z(n335) );
  XNOR2_X1 U392 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U393 ( .A(n337), .B(KEYINPUT31), .Z(n339) );
  XOR2_X1 U394 ( .A(G120GAT), .B(G148GAT), .Z(n402) );
  XNOR2_X1 U395 ( .A(KEYINPUT33), .B(n402), .ZN(n338) );
  XNOR2_X1 U396 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U397 ( .A(KEYINPUT45), .B(KEYINPUT111), .ZN(n380) );
  XNOR2_X1 U398 ( .A(n341), .B(G64GAT), .ZN(n342) );
  XNOR2_X1 U399 ( .A(n342), .B(KEYINPUT12), .ZN(n356) );
  XOR2_X1 U400 ( .A(n343), .B(KEYINPUT77), .Z(n345) );
  NAND2_X1 U401 ( .A1(G231GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U402 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U403 ( .A(KEYINPUT14), .B(KEYINPUT76), .Z(n347) );
  XNOR2_X1 U404 ( .A(KEYINPUT15), .B(KEYINPUT78), .ZN(n346) );
  XNOR2_X1 U405 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U406 ( .A(n349), .B(n348), .Z(n354) );
  XOR2_X1 U407 ( .A(G155GAT), .B(G57GAT), .Z(n351) );
  XNOR2_X1 U408 ( .A(G1GAT), .B(G127GAT), .ZN(n350) );
  XNOR2_X1 U409 ( .A(n351), .B(n350), .ZN(n408) );
  XNOR2_X1 U410 ( .A(n408), .B(n352), .ZN(n353) );
  XNOR2_X1 U411 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U412 ( .A(n356), .B(n355), .Z(n560) );
  INV_X1 U413 ( .A(n560), .ZN(n584) );
  XOR2_X1 U414 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n358) );
  XNOR2_X1 U415 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n357) );
  XNOR2_X1 U416 ( .A(n358), .B(n357), .ZN(n362) );
  XOR2_X1 U417 ( .A(KEYINPUT64), .B(KEYINPUT72), .Z(n360) );
  XNOR2_X1 U418 ( .A(KEYINPUT75), .B(KEYINPUT71), .ZN(n359) );
  XNOR2_X1 U419 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U420 ( .A(G162GAT), .B(G92GAT), .Z(n364) );
  NAND2_X1 U421 ( .A1(G232GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U422 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U423 ( .A(KEYINPUT73), .B(n365), .ZN(n366) );
  XNOR2_X1 U424 ( .A(n294), .B(n366), .ZN(n370) );
  XOR2_X1 U425 ( .A(G29GAT), .B(G134GAT), .Z(n403) );
  XOR2_X1 U426 ( .A(G50GAT), .B(KEYINPUT70), .Z(n417) );
  XOR2_X1 U427 ( .A(n403), .B(n417), .Z(n368) );
  NAND2_X1 U428 ( .A1(n371), .A2(n372), .ZN(n376) );
  INV_X1 U429 ( .A(n371), .ZN(n374) );
  INV_X1 U430 ( .A(n372), .ZN(n373) );
  NAND2_X1 U431 ( .A1(n374), .A2(n373), .ZN(n375) );
  AND2_X1 U432 ( .A1(n376), .A2(n375), .ZN(n378) );
  NOR2_X1 U433 ( .A1(n584), .A2(n587), .ZN(n379) );
  XOR2_X1 U434 ( .A(n380), .B(n379), .Z(n381) );
  NAND2_X1 U435 ( .A1(n580), .A2(n381), .ZN(n382) );
  NOR2_X1 U436 ( .A1(n551), .A2(n382), .ZN(n384) );
  XNOR2_X1 U437 ( .A(n384), .B(n383), .ZN(n390) );
  XOR2_X1 U438 ( .A(KEYINPUT41), .B(n580), .Z(n453) );
  INV_X1 U439 ( .A(n453), .ZN(n555) );
  NAND2_X1 U440 ( .A1(n551), .A2(n555), .ZN(n385) );
  XNOR2_X1 U441 ( .A(n385), .B(KEYINPUT46), .ZN(n386) );
  XOR2_X1 U442 ( .A(KEYINPUT110), .B(n560), .Z(n539) );
  NAND2_X1 U443 ( .A1(n386), .A2(n539), .ZN(n387) );
  XNOR2_X1 U444 ( .A(KEYINPUT47), .B(n388), .ZN(n389) );
  NAND2_X1 U445 ( .A1(n390), .A2(n389), .ZN(n391) );
  NAND2_X1 U446 ( .A1(n392), .A2(n548), .ZN(n393) );
  XNOR2_X1 U447 ( .A(n393), .B(KEYINPUT54), .ZN(n415) );
  XOR2_X1 U448 ( .A(KEYINPUT6), .B(KEYINPUT84), .Z(n395) );
  XNOR2_X1 U449 ( .A(KEYINPUT88), .B(KEYINPUT89), .ZN(n394) );
  XNOR2_X1 U450 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U451 ( .A(n396), .B(KEYINPUT87), .Z(n398) );
  XOR2_X1 U452 ( .A(G113GAT), .B(KEYINPUT0), .Z(n440) );
  XNOR2_X1 U453 ( .A(n440), .B(G85GAT), .ZN(n397) );
  XNOR2_X1 U454 ( .A(n398), .B(n397), .ZN(n401) );
  XOR2_X1 U455 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n400) );
  XNOR2_X1 U456 ( .A(G141GAT), .B(G162GAT), .ZN(n399) );
  XNOR2_X1 U457 ( .A(n400), .B(n399), .ZN(n416) );
  XOR2_X1 U458 ( .A(n401), .B(n416), .Z(n405) );
  XNOR2_X1 U459 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U460 ( .A(n405), .B(n404), .ZN(n414) );
  XOR2_X1 U461 ( .A(KEYINPUT86), .B(KEYINPUT1), .Z(n407) );
  XNOR2_X1 U462 ( .A(KEYINPUT85), .B(KEYINPUT4), .ZN(n406) );
  XNOR2_X1 U463 ( .A(n407), .B(n406), .ZN(n412) );
  XOR2_X1 U464 ( .A(KEYINPUT5), .B(n408), .Z(n410) );
  NAND2_X1 U465 ( .A1(G225GAT), .A2(G233GAT), .ZN(n409) );
  XNOR2_X1 U466 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U467 ( .A(n412), .B(n411), .Z(n413) );
  XNOR2_X1 U468 ( .A(n414), .B(n413), .ZN(n467) );
  XOR2_X1 U469 ( .A(KEYINPUT90), .B(n467), .Z(n550) );
  INV_X1 U470 ( .A(n550), .ZN(n519) );
  XOR2_X1 U471 ( .A(n416), .B(G204GAT), .Z(n419) );
  XNOR2_X1 U472 ( .A(G106GAT), .B(n417), .ZN(n418) );
  XNOR2_X1 U473 ( .A(n419), .B(n418), .ZN(n424) );
  XOR2_X1 U474 ( .A(n420), .B(KEYINPUT23), .Z(n422) );
  NAND2_X1 U475 ( .A1(G228GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U476 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U477 ( .A(n424), .B(n423), .Z(n432) );
  XOR2_X1 U478 ( .A(G148GAT), .B(G78GAT), .Z(n426) );
  XNOR2_X1 U479 ( .A(G22GAT), .B(G155GAT), .ZN(n425) );
  XNOR2_X1 U480 ( .A(n426), .B(n425), .ZN(n430) );
  XOR2_X1 U481 ( .A(KEYINPUT83), .B(KEYINPUT22), .Z(n428) );
  XNOR2_X1 U482 ( .A(G211GAT), .B(KEYINPUT24), .ZN(n427) );
  XNOR2_X1 U483 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U485 ( .A(n432), .B(n431), .ZN(n468) );
  NAND2_X1 U486 ( .A1(n575), .A2(n468), .ZN(n434) );
  XOR2_X1 U487 ( .A(KEYINPUT55), .B(KEYINPUT121), .Z(n433) );
  XOR2_X1 U488 ( .A(G183GAT), .B(G127GAT), .Z(n436) );
  XNOR2_X1 U489 ( .A(G15GAT), .B(G120GAT), .ZN(n435) );
  XNOR2_X1 U490 ( .A(n436), .B(n435), .ZN(n451) );
  XOR2_X1 U491 ( .A(G71GAT), .B(G176GAT), .Z(n438) );
  XNOR2_X1 U492 ( .A(G134GAT), .B(G99GAT), .ZN(n437) );
  XNOR2_X1 U493 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U494 ( .A(n439), .B(G190GAT), .Z(n442) );
  XNOR2_X1 U495 ( .A(G43GAT), .B(n440), .ZN(n441) );
  XNOR2_X1 U496 ( .A(n442), .B(n441), .ZN(n446) );
  XOR2_X1 U497 ( .A(KEYINPUT20), .B(KEYINPUT81), .Z(n444) );
  NAND2_X1 U498 ( .A1(G227GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U499 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U500 ( .A(n446), .B(n445), .Z(n449) );
  XOR2_X1 U501 ( .A(n447), .B(KEYINPUT79), .Z(n448) );
  XNOR2_X1 U502 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X2 U503 ( .A(n451), .B(n450), .Z(n531) );
  NAND2_X1 U504 ( .A1(n452), .A2(n531), .ZN(n569) );
  NOR2_X1 U505 ( .A1(n569), .A2(n453), .ZN(n456) );
  XNOR2_X1 U506 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n454) );
  XNOR2_X1 U507 ( .A(n454), .B(G176GAT), .ZN(n455) );
  XNOR2_X1 U508 ( .A(n456), .B(n455), .ZN(G1349GAT) );
  NOR2_X1 U509 ( .A1(n539), .A2(n569), .ZN(n459) );
  XNOR2_X1 U510 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n457) );
  XNOR2_X1 U511 ( .A(KEYINPUT34), .B(KEYINPUT94), .ZN(n480) );
  XOR2_X1 U512 ( .A(G1GAT), .B(KEYINPUT95), .Z(n478) );
  NAND2_X1 U513 ( .A1(n551), .A2(n580), .ZN(n493) );
  NOR2_X1 U514 ( .A1(n568), .A2(n584), .ZN(n460) );
  XNOR2_X1 U515 ( .A(n460), .B(KEYINPUT16), .ZN(n475) );
  XOR2_X1 U516 ( .A(KEYINPUT27), .B(n523), .Z(n470) );
  NOR2_X1 U517 ( .A1(n468), .A2(n531), .ZN(n461) );
  XNOR2_X1 U518 ( .A(n461), .B(KEYINPUT26), .ZN(n576) );
  INV_X1 U519 ( .A(n576), .ZN(n462) );
  NOR2_X1 U520 ( .A1(n470), .A2(n462), .ZN(n547) );
  NAND2_X1 U521 ( .A1(n531), .A2(n523), .ZN(n463) );
  NAND2_X1 U522 ( .A1(n468), .A2(n463), .ZN(n464) );
  XNOR2_X1 U523 ( .A(KEYINPUT25), .B(n464), .ZN(n465) );
  NOR2_X1 U524 ( .A1(n547), .A2(n465), .ZN(n466) );
  NOR2_X1 U525 ( .A1(n467), .A2(n466), .ZN(n473) );
  XNOR2_X1 U526 ( .A(n468), .B(KEYINPUT65), .ZN(n469) );
  XNOR2_X1 U527 ( .A(n469), .B(KEYINPUT28), .ZN(n527) );
  NOR2_X1 U528 ( .A1(n527), .A2(n470), .ZN(n471) );
  NAND2_X1 U529 ( .A1(n519), .A2(n471), .ZN(n533) );
  NOR2_X1 U530 ( .A1(n531), .A2(n533), .ZN(n472) );
  NOR2_X1 U531 ( .A1(n473), .A2(n472), .ZN(n490) );
  INV_X1 U532 ( .A(n490), .ZN(n474) );
  NAND2_X1 U533 ( .A1(n475), .A2(n474), .ZN(n506) );
  NOR2_X1 U534 ( .A1(n493), .A2(n506), .ZN(n476) );
  XOR2_X1 U535 ( .A(KEYINPUT93), .B(n476), .Z(n485) );
  NAND2_X1 U536 ( .A1(n485), .A2(n519), .ZN(n477) );
  XNOR2_X1 U537 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U538 ( .A(n480), .B(n479), .ZN(G1324GAT) );
  NAND2_X1 U539 ( .A1(n523), .A2(n485), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n481), .B(KEYINPUT96), .ZN(n482) );
  XNOR2_X1 U541 ( .A(G8GAT), .B(n482), .ZN(G1325GAT) );
  XOR2_X1 U542 ( .A(G15GAT), .B(KEYINPUT35), .Z(n484) );
  NAND2_X1 U543 ( .A1(n485), .A2(n531), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n484), .B(n483), .ZN(G1326GAT) );
  XOR2_X1 U545 ( .A(G22GAT), .B(KEYINPUT97), .Z(n487) );
  NAND2_X1 U546 ( .A1(n485), .A2(n527), .ZN(n486) );
  XNOR2_X1 U547 ( .A(n487), .B(n486), .ZN(G1327GAT) );
  XOR2_X1 U548 ( .A(KEYINPUT98), .B(KEYINPUT101), .Z(n489) );
  XNOR2_X1 U549 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n489), .B(n488), .ZN(n498) );
  NOR2_X1 U551 ( .A1(n587), .A2(n490), .ZN(n491) );
  NAND2_X1 U552 ( .A1(n491), .A2(n584), .ZN(n492) );
  XOR2_X1 U553 ( .A(KEYINPUT37), .B(n492), .Z(n518) );
  NOR2_X1 U554 ( .A1(n518), .A2(n493), .ZN(n495) );
  XNOR2_X1 U555 ( .A(KEYINPUT100), .B(KEYINPUT38), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U557 ( .A(KEYINPUT99), .B(n496), .Z(n504) );
  NAND2_X1 U558 ( .A1(n504), .A2(n519), .ZN(n497) );
  XOR2_X1 U559 ( .A(n498), .B(n497), .Z(G1328GAT) );
  NAND2_X1 U560 ( .A1(n523), .A2(n504), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n499), .B(KEYINPUT102), .ZN(n500) );
  XNOR2_X1 U562 ( .A(G36GAT), .B(n500), .ZN(G1329GAT) );
  XOR2_X1 U563 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n502) );
  NAND2_X1 U564 ( .A1(n504), .A2(n531), .ZN(n501) );
  XNOR2_X1 U565 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U566 ( .A(G43GAT), .B(n503), .ZN(G1330GAT) );
  NAND2_X1 U567 ( .A1(n504), .A2(n527), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n505), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n509) );
  INV_X1 U570 ( .A(n551), .ZN(n577) );
  NAND2_X1 U571 ( .A1(n577), .A2(n555), .ZN(n517) );
  NOR2_X1 U572 ( .A1(n517), .A2(n506), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n507), .B(KEYINPUT104), .ZN(n513) );
  NAND2_X1 U574 ( .A1(n519), .A2(n513), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n509), .B(n508), .ZN(G1332GAT) );
  XOR2_X1 U576 ( .A(G64GAT), .B(KEYINPUT105), .Z(n511) );
  NAND2_X1 U577 ( .A1(n513), .A2(n523), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n511), .B(n510), .ZN(G1333GAT) );
  NAND2_X1 U579 ( .A1(n513), .A2(n531), .ZN(n512) );
  XNOR2_X1 U580 ( .A(n512), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n515) );
  NAND2_X1 U582 ( .A1(n527), .A2(n513), .ZN(n514) );
  XNOR2_X1 U583 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U584 ( .A(G78GAT), .B(n516), .ZN(G1335GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n521) );
  NOR2_X1 U586 ( .A1(n518), .A2(n517), .ZN(n528) );
  NAND2_X1 U587 ( .A1(n528), .A2(n519), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U589 ( .A(G85GAT), .B(n522), .ZN(G1336GAT) );
  NAND2_X1 U590 ( .A1(n523), .A2(n528), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n524), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U592 ( .A(G99GAT), .B(KEYINPUT109), .Z(n526) );
  NAND2_X1 U593 ( .A1(n528), .A2(n531), .ZN(n525) );
  XNOR2_X1 U594 ( .A(n526), .B(n525), .ZN(G1338GAT) );
  NAND2_X1 U595 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n529), .B(KEYINPUT44), .ZN(n530) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(n530), .ZN(G1339GAT) );
  NAND2_X1 U598 ( .A1(n531), .A2(n548), .ZN(n532) );
  NOR2_X1 U599 ( .A1(n533), .A2(n532), .ZN(n543) );
  NAND2_X1 U600 ( .A1(n543), .A2(n551), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n534), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT113), .B(KEYINPUT49), .Z(n536) );
  NAND2_X1 U603 ( .A1(n543), .A2(n555), .ZN(n535) );
  XNOR2_X1 U604 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U605 ( .A(G120GAT), .B(n537), .Z(G1341GAT) );
  INV_X1 U606 ( .A(n543), .ZN(n538) );
  NOR2_X1 U607 ( .A1(n539), .A2(n538), .ZN(n541) );
  XNOR2_X1 U608 ( .A(KEYINPUT114), .B(KEYINPUT50), .ZN(n540) );
  XNOR2_X1 U609 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U610 ( .A(G127GAT), .B(n542), .Z(G1342GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n545) );
  NAND2_X1 U612 ( .A1(n543), .A2(n568), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U614 ( .A(G134GAT), .B(n546), .Z(G1343GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n553) );
  NAND2_X1 U616 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n563) );
  NAND2_X1 U618 ( .A1(n563), .A2(n551), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G141GAT), .B(n554), .ZN(G1344GAT) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n559) );
  XOR2_X1 U622 ( .A(KEYINPUT52), .B(KEYINPUT118), .Z(n557) );
  NAND2_X1 U623 ( .A1(n563), .A2(n555), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(G1345GAT) );
  XOR2_X1 U626 ( .A(G155GAT), .B(KEYINPUT119), .Z(n562) );
  NAND2_X1 U627 ( .A1(n563), .A2(n560), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1346GAT) );
  NAND2_X1 U629 ( .A1(n563), .A2(n568), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U631 ( .A1(n577), .A2(n569), .ZN(n565) );
  XOR2_X1 U632 ( .A(G169GAT), .B(n565), .Z(G1348GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n567) );
  XNOR2_X1 U634 ( .A(G190GAT), .B(KEYINPUT125), .ZN(n566) );
  XNOR2_X1 U635 ( .A(n567), .B(n566), .ZN(n572) );
  INV_X1 U636 ( .A(n568), .ZN(n570) );
  NOR2_X1 U637 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U638 ( .A(n572), .B(n571), .Z(G1351GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n574) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n573) );
  XNOR2_X1 U641 ( .A(n574), .B(n573), .ZN(n579) );
  NAND2_X1 U642 ( .A1(n575), .A2(n576), .ZN(n586) );
  NOR2_X1 U643 ( .A1(n577), .A2(n586), .ZN(n578) );
  XOR2_X1 U644 ( .A(n579), .B(n578), .Z(G1352GAT) );
  NOR2_X1 U645 ( .A1(n580), .A2(n586), .ZN(n582) );
  XNOR2_X1 U646 ( .A(KEYINPUT61), .B(KEYINPUT127), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XOR2_X1 U648 ( .A(G204GAT), .B(n583), .Z(G1353GAT) );
  NOR2_X1 U649 ( .A1(n584), .A2(n586), .ZN(n585) );
  XOR2_X1 U650 ( .A(G211GAT), .B(n585), .Z(G1354GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U652 ( .A(KEYINPUT62), .B(n588), .Z(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

