//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1191, new_n1192, new_n1193, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G250), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT65), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  INV_X1    g0014(.A(G264), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n209), .B(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(KEYINPUT0), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G20), .ZN(new_n220));
  INV_X1    g0020(.A(G58), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(G50), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n217), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G58), .B2(G232), .ZN(new_n226));
  INV_X1    g0026(.A(G238), .ZN(new_n227));
  INV_X1    g0027(.A(G244), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n226), .B1(new_n222), .B2(new_n227), .C1(new_n202), .C2(new_n228), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n230), .B1(new_n205), .B2(new_n214), .C1(new_n206), .C2(new_n215), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n211), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT1), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n216), .A2(KEYINPUT0), .ZN(new_n234));
  NOR3_X1   g0034(.A1(new_n225), .A2(new_n233), .A3(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G226), .ZN(new_n238));
  INV_X1    g0038(.A(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT66), .ZN(new_n246));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(G1), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G13), .A3(G20), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT69), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND4_X1  g0056(.A1(new_n253), .A2(KEYINPUT69), .A3(G13), .A4(G20), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n218), .B1(new_n210), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G20), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n258), .B(new_n261), .C1(G1), .C2(new_n262), .ZN(new_n263));
  OR2_X1    g0063(.A1(new_n263), .A2(new_n202), .ZN(new_n264));
  AND2_X1   g0064(.A1(new_n256), .A2(new_n257), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n202), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT8), .B(G58), .ZN(new_n267));
  NOR3_X1   g0067(.A1(new_n267), .A2(G20), .A3(G33), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT15), .B(G87), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n262), .A2(G33), .ZN(new_n270));
  OAI22_X1  g0070(.A1(new_n269), .A2(new_n270), .B1(new_n262), .B2(new_n202), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n260), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n264), .A2(new_n266), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n218), .B1(G33), .B2(G41), .ZN(new_n274));
  INV_X1    g0074(.A(G274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n253), .B1(G41), .B2(G45), .ZN(new_n276));
  NOR3_X1   g0076(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(new_n276), .B(KEYINPUT67), .ZN(new_n279));
  INV_X1    g0079(.A(G41), .ZN(new_n280));
  OAI211_X1 g0080(.A(G1), .B(G13), .C1(new_n259), .C2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n278), .B1(new_n282), .B2(new_n228), .ZN(new_n283));
  XNOR2_X1  g0083(.A(new_n283), .B(KEYINPUT70), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT3), .B(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G1698), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT68), .ZN(new_n287));
  XNOR2_X1  g0087(.A(new_n286), .B(new_n287), .ZN(new_n288));
  AND2_X1   g0088(.A1(new_n288), .A2(G238), .ZN(new_n289));
  INV_X1    g0089(.A(G1698), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n285), .A2(new_n290), .ZN(new_n291));
  OR3_X1    g0091(.A1(new_n291), .A2(KEYINPUT71), .A3(new_n239), .ZN(new_n292));
  OAI21_X1  g0092(.A(KEYINPUT71), .B1(new_n291), .B2(new_n239), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n292), .B(new_n293), .C1(new_n206), .C2(new_n285), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n274), .B1(new_n289), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n284), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n273), .B1(new_n297), .B2(G190), .ZN(new_n298));
  INV_X1    g0098(.A(G200), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n298), .B1(new_n299), .B2(new_n297), .ZN(new_n300));
  INV_X1    g0100(.A(G179), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G169), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n296), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n302), .A2(new_n304), .A3(new_n273), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT16), .ZN(new_n307));
  NAND2_X1  g0107(.A1(G58), .A2(G68), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT74), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n308), .B(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n223), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G20), .ZN(new_n312));
  NOR2_X1   g0112(.A1(G20), .A2(G33), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G159), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT7), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n316), .B1(new_n285), .B2(G20), .ZN(new_n317));
  AND2_X1   g0117(.A1(KEYINPUT3), .A2(G33), .ZN(new_n318));
  NOR2_X1   g0118(.A1(KEYINPUT3), .A2(G33), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n320), .A2(KEYINPUT7), .A3(new_n262), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n222), .B1(new_n317), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n307), .B1(new_n315), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n322), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n324), .A2(KEYINPUT16), .A3(new_n314), .A4(new_n312), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n323), .A2(new_n325), .A3(new_n260), .ZN(new_n326));
  INV_X1    g0126(.A(G226), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G1698), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n328), .B1(G223), .B2(G1698), .ZN(new_n329));
  INV_X1    g0129(.A(G87), .ZN(new_n330));
  OAI22_X1  g0130(.A1(new_n329), .A2(new_n320), .B1(new_n259), .B2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n277), .B1(new_n331), .B2(new_n274), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n279), .A2(G232), .A3(new_n281), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G200), .ZN(new_n335));
  INV_X1    g0135(.A(new_n267), .ZN(new_n336));
  MUX2_X1   g0136(.A(new_n258), .B(new_n263), .S(new_n336), .Z(new_n337));
  INV_X1    g0137(.A(new_n334), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(G190), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n326), .A2(new_n335), .A3(new_n337), .A4(new_n339), .ZN(new_n340));
  XNOR2_X1  g0140(.A(new_n340), .B(KEYINPUT17), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n326), .A2(new_n337), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n334), .A2(G179), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n343), .B1(new_n303), .B2(new_n334), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT18), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT18), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n342), .A2(new_n344), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n306), .A2(new_n341), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n288), .A2(G223), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n320), .A2(G1698), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n353), .A2(G222), .B1(G77), .B2(new_n320), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n281), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n278), .B1(new_n282), .B2(new_n327), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n357), .A2(new_n299), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n358), .B1(G190), .B2(new_n357), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT72), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT10), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n313), .A2(G150), .ZN(new_n362));
  OAI221_X1 g0162(.A(new_n362), .B1(new_n201), .B2(new_n262), .C1(new_n267), .C2(new_n270), .ZN(new_n363));
  INV_X1    g0163(.A(G50), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n363), .A2(new_n260), .B1(new_n265), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(new_n364), .B2(new_n263), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n366), .B(KEYINPUT9), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n359), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n361), .A2(new_n368), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n359), .B(new_n367), .C1(new_n360), .C2(KEYINPUT10), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n357), .A2(new_n301), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n303), .B1(new_n355), .B2(new_n356), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n371), .A2(new_n366), .A3(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n369), .A2(new_n370), .A3(new_n373), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n313), .A2(G50), .B1(G20), .B2(new_n222), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(new_n202), .B2(new_n270), .ZN(new_n376));
  AND2_X1   g0176(.A1(new_n376), .A2(new_n260), .ZN(new_n377));
  OR2_X1    g0177(.A1(new_n377), .A2(KEYINPUT11), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(KEYINPUT11), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n265), .A2(KEYINPUT12), .A3(new_n222), .ZN(new_n380));
  OR2_X1    g0180(.A1(new_n265), .A2(KEYINPUT12), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n378), .A2(new_n379), .A3(new_n380), .A4(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n222), .B1(new_n263), .B2(KEYINPUT12), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT73), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(new_n259), .B2(new_n205), .ZN(new_n387));
  NAND3_X1  g0187(.A1(KEYINPUT73), .A2(G33), .A3(G97), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n239), .A2(G1698), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(G226), .B2(G1698), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n389), .B1(new_n391), .B2(new_n320), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n277), .B1(new_n392), .B2(new_n274), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(new_n227), .B2(new_n282), .ZN(new_n394));
  XNOR2_X1  g0194(.A(new_n394), .B(KEYINPUT13), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(G169), .ZN(new_n396));
  OAI22_X1  g0196(.A1(new_n396), .A2(KEYINPUT14), .B1(new_n301), .B2(new_n395), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n396), .A2(KEYINPUT14), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n385), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n395), .A2(G200), .ZN(new_n400));
  INV_X1    g0200(.A(G190), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n400), .B(new_n384), .C1(new_n401), .C2(new_n395), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  NOR3_X1   g0203(.A1(new_n351), .A2(new_n374), .A3(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT82), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n265), .A2(new_n405), .A3(new_n206), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT25), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT82), .B1(new_n258), .B2(G107), .ZN(new_n408));
  AND3_X1   g0208(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n407), .B1(new_n406), .B2(new_n408), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n253), .A2(G33), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n258), .A2(new_n261), .A3(new_n411), .ZN(new_n412));
  OAI22_X1  g0212(.A1(new_n409), .A2(new_n410), .B1(new_n206), .B2(new_n412), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n262), .B(G87), .C1(new_n318), .C2(new_n319), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT22), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT22), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n285), .A2(new_n416), .A3(new_n262), .A4(G87), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT24), .ZN(new_n419));
  AOI21_X1  g0219(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT23), .ZN(new_n421));
  OAI22_X1  g0221(.A1(new_n420), .A2(G20), .B1(new_n421), .B2(new_n206), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n421), .A2(new_n206), .A3(G20), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT80), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n421), .A2(new_n206), .A3(KEYINPUT80), .A4(G20), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n422), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n418), .A2(new_n419), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n419), .B1(new_n418), .B2(new_n427), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n260), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT81), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT81), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n432), .B(new_n260), .C1(new_n428), .C2(new_n429), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n413), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  OAI211_X1 g0234(.A(G257), .B(G1698), .C1(new_n318), .C2(new_n319), .ZN(new_n435));
  OAI211_X1 g0235(.A(G250), .B(new_n290), .C1(new_n318), .C2(new_n319), .ZN(new_n436));
  NAND2_X1  g0236(.A1(G33), .A2(G294), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT83), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT83), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n435), .A2(new_n436), .A3(new_n440), .A4(new_n437), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n439), .A2(new_n274), .A3(new_n441), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n253), .B(G45), .C1(new_n280), .C2(KEYINPUT5), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n280), .A2(KEYINPUT5), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n281), .B(G264), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  XNOR2_X1  g0245(.A(new_n445), .B(KEYINPUT84), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n443), .A2(new_n444), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n447), .A2(G274), .A3(new_n281), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n442), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n303), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(G179), .B2(new_n449), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n434), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n431), .A2(new_n433), .ZN(new_n454));
  INV_X1    g0254(.A(new_n413), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n449), .A2(new_n299), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n442), .A2(new_n446), .A3(new_n401), .A4(new_n448), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AND4_X1   g0258(.A1(KEYINPUT85), .A2(new_n454), .A3(new_n455), .A4(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(KEYINPUT85), .B1(new_n434), .B2(new_n458), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n453), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT86), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT86), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n453), .B(new_n463), .C1(new_n459), .C2(new_n460), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(G264), .A2(G1698), .ZN(new_n466));
  OAI221_X1 g0266(.A(new_n466), .B1(new_n214), .B2(G1698), .C1(new_n318), .C2(new_n319), .ZN(new_n467));
  INV_X1    g0267(.A(G303), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n320), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n467), .A2(new_n469), .A3(new_n274), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT77), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT77), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n467), .A2(new_n469), .A3(new_n472), .A4(new_n274), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  OR2_X1    g0274(.A1(new_n443), .A2(new_n444), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n475), .A2(G270), .A3(new_n281), .ZN(new_n476));
  AND2_X1   g0276(.A1(new_n476), .A2(new_n448), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT78), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n474), .A2(new_n477), .A3(KEYINPUT78), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G190), .ZN(new_n483));
  NAND2_X1  g0283(.A1(G33), .A2(G283), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n484), .B(new_n262), .C1(G33), .C2(new_n205), .ZN(new_n485));
  INV_X1    g0285(.A(G116), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G20), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n485), .A2(new_n260), .A3(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT20), .ZN(new_n489));
  OR2_X1    g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(new_n489), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n490), .A2(new_n491), .B1(new_n486), .B2(new_n265), .ZN(new_n492));
  INV_X1    g0292(.A(new_n412), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G116), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n483), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n482), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n496), .B1(G200), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n303), .B1(new_n492), .B2(new_n494), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n480), .A2(new_n481), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT21), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n480), .A2(KEYINPUT21), .A3(new_n481), .A4(new_n499), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n474), .A2(new_n477), .A3(G179), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n495), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n505), .A2(KEYINPUT79), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT79), .ZN(new_n507));
  NOR3_X1   g0307(.A1(new_n495), .A2(new_n504), .A3(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n502), .B(new_n503), .C1(new_n506), .C2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n313), .A2(G77), .ZN(new_n510));
  XNOR2_X1  g0310(.A(KEYINPUT75), .B(KEYINPUT6), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G97), .A2(G107), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n511), .A2(new_n207), .A3(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n205), .A2(G107), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n513), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n510), .B1(new_n515), .B2(new_n262), .ZN(new_n516));
  NOR3_X1   g0316(.A1(new_n285), .A2(new_n316), .A3(G20), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT7), .B1(new_n320), .B2(new_n262), .ZN(new_n518));
  OAI21_X1  g0318(.A(G107), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n260), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n258), .A2(G97), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n412), .B2(new_n205), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n521), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n285), .A2(KEYINPUT4), .A3(G244), .A4(new_n290), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n320), .A2(new_n228), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n527), .B(new_n484), .C1(new_n528), .C2(KEYINPUT4), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n285), .A2(G250), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n290), .B1(new_n530), .B2(KEYINPUT4), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n274), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n475), .A2(G257), .A3(new_n281), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n533), .A2(new_n448), .ZN(new_n534));
  AND3_X1   g0334(.A1(new_n532), .A2(G179), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n303), .B1(new_n532), .B2(new_n534), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n526), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n532), .A2(new_n534), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G200), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n519), .B(new_n510), .C1(new_n262), .C2(new_n515), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n524), .B1(new_n540), .B2(new_n260), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n532), .A2(G190), .A3(new_n534), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n539), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n537), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n285), .A2(G244), .A3(G1698), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT76), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n285), .A2(KEYINPUT76), .A3(G244), .A4(G1698), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n353), .A2(G238), .B1(G33), .B2(G116), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n281), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(G45), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n209), .B1(new_n552), .B2(G1), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n253), .A2(new_n275), .A3(G45), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n281), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(G200), .B1(new_n551), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G33), .A2(G116), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n291), .B2(new_n227), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n559), .B1(new_n547), .B2(new_n548), .ZN(new_n560));
  OAI211_X1 g0360(.A(G190), .B(new_n555), .C1(new_n560), .C2(new_n281), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n285), .A2(new_n262), .A3(G68), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n270), .A2(new_n205), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n562), .B1(KEYINPUT19), .B2(new_n563), .ZN(new_n564));
  NOR3_X1   g0364(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n387), .A2(KEYINPUT19), .A3(new_n388), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n565), .B1(new_n566), .B2(new_n262), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n260), .B1(new_n564), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n265), .A2(new_n269), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n412), .A2(new_n330), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n557), .A2(new_n561), .A3(new_n571), .A4(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n301), .B(new_n555), .C1(new_n560), .C2(new_n281), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n568), .B(new_n569), .C1(new_n269), .C2(new_n412), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n549), .A2(new_n550), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n556), .B1(new_n577), .B2(new_n274), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n575), .B(new_n576), .C1(new_n578), .C2(G169), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  NOR4_X1   g0380(.A1(new_n498), .A2(new_n509), .A3(new_n544), .A4(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n404), .A2(new_n465), .A3(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(G372));
  NAND4_X1  g0383(.A1(new_n402), .A2(new_n304), .A3(new_n302), .A4(new_n273), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n399), .A2(new_n584), .ZN(new_n585));
  OR2_X1    g0385(.A1(new_n585), .A2(KEYINPUT92), .ZN(new_n586));
  XOR2_X1   g0386(.A(new_n340), .B(KEYINPUT17), .Z(new_n587));
  AOI21_X1  g0387(.A(new_n587), .B1(new_n585), .B2(KEYINPUT92), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n349), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n369), .A2(new_n370), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n373), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n509), .A2(new_n452), .ZN(new_n593));
  XNOR2_X1  g0393(.A(new_n555), .B(KEYINPUT87), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n560), .B2(new_n281), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n303), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n596), .A2(new_n575), .A3(new_n576), .ZN(new_n597));
  INV_X1    g0397(.A(new_n594), .ZN(new_n598));
  OAI21_X1  g0398(.A(G200), .B1(new_n551), .B2(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n599), .A2(new_n561), .A3(new_n571), .A4(new_n573), .ZN(new_n600));
  AND4_X1   g0400(.A1(new_n537), .A2(new_n597), .A3(new_n543), .A4(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n459), .B2(new_n460), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n593), .B1(new_n602), .B2(KEYINPUT88), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT88), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n601), .B(new_n604), .C1(new_n459), .C2(new_n460), .ZN(new_n605));
  AOI21_X1  g0405(.A(KEYINPUT89), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n602), .A2(KEYINPUT88), .ZN(new_n607));
  OR2_X1    g0407(.A1(new_n509), .A2(new_n452), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n607), .A2(KEYINPUT89), .A3(new_n605), .A4(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n597), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n538), .A2(G169), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n532), .A2(G179), .A3(new_n534), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n579), .A2(new_n574), .A3(new_n613), .A4(new_n526), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n610), .B1(new_n614), .B2(KEYINPUT26), .ZN(new_n615));
  OAI21_X1  g0415(.A(KEYINPUT90), .B1(new_n535), .B2(new_n536), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT90), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n611), .A2(new_n617), .A3(new_n612), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n541), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n575), .A2(new_n576), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n572), .B1(new_n595), .B2(G200), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n570), .B1(new_n578), .B2(G190), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n620), .A2(new_n596), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT26), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n619), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n615), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(KEYINPUT91), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT91), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n615), .A2(new_n625), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n609), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n404), .B1(new_n606), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n592), .A2(new_n632), .ZN(G369));
  NOR2_X1   g0433(.A1(new_n498), .A2(new_n509), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n253), .A2(new_n262), .A3(G13), .ZN(new_n635));
  OR2_X1    g0435(.A1(new_n635), .A2(KEYINPUT27), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(KEYINPUT27), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n636), .A2(G213), .A3(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(G343), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n495), .A2(new_n641), .ZN(new_n642));
  MUX2_X1   g0442(.A(new_n634), .B(new_n509), .S(new_n642), .Z(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(G330), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n465), .B1(new_n434), .B2(new_n641), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n452), .A2(new_n640), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n453), .A2(new_n640), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n509), .A2(new_n641), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n650), .B1(new_n465), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n649), .A2(new_n652), .ZN(G399));
  NOR2_X1   g0453(.A1(new_n213), .A2(G41), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n565), .A2(new_n486), .ZN(new_n655));
  NOR3_X1   g0455(.A1(new_n654), .A2(new_n253), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n224), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n656), .B1(new_n657), .B2(new_n654), .ZN(new_n658));
  XOR2_X1   g0458(.A(new_n658), .B(KEYINPUT28), .Z(new_n659));
  AOI21_X1  g0459(.A(new_n624), .B1(new_n619), .B2(new_n623), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n597), .B1(new_n614), .B2(KEYINPUT26), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n602), .B2(new_n593), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n641), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT29), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n641), .B1(new_n631), .B2(new_n606), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n666), .B1(new_n667), .B2(new_n665), .ZN(new_n668));
  INV_X1    g0468(.A(G330), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n595), .A2(new_n538), .A3(new_n301), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n497), .A2(new_n449), .A3(new_n670), .ZN(new_n671));
  NOR3_X1   g0471(.A1(new_n478), .A2(new_n551), .A3(new_n556), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n442), .A2(new_n446), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n672), .A2(KEYINPUT30), .A3(new_n673), .A4(new_n535), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT30), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n673), .A2(new_n578), .A3(new_n474), .A4(new_n477), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n675), .B1(new_n676), .B2(new_n612), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n671), .A2(new_n674), .A3(new_n677), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n678), .A2(KEYINPUT31), .A3(new_n640), .ZN(new_n679));
  AOI21_X1  g0479(.A(KEYINPUT31), .B1(new_n678), .B2(new_n640), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT93), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n678), .A2(new_n640), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT31), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT93), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n678), .A2(KEYINPUT31), .A3(new_n640), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n681), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n465), .A2(new_n581), .A3(new_n641), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n669), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n668), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n659), .B1(new_n691), .B2(G1), .ZN(G364));
  AND2_X1   g0492(.A1(new_n262), .A2(G13), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n253), .B1(new_n693), .B2(G45), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n654), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n645), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(G330), .B2(new_n643), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n218), .B1(G20), .B2(new_n303), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n699), .A2(KEYINPUT95), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(KEYINPUT95), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(G13), .A2(G33), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(G20), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n212), .A2(new_n285), .ZN(new_n708));
  XOR2_X1   g0508(.A(new_n708), .B(KEYINPUT94), .Z(new_n709));
  AOI22_X1  g0509(.A1(new_n709), .A2(G355), .B1(new_n486), .B2(new_n213), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n212), .A2(new_n320), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n711), .B1(new_n552), .B2(new_n657), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n248), .B2(new_n552), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n707), .B1(new_n710), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n702), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n262), .A2(G179), .ZN(new_n716));
  NOR2_X1   g0516(.A1(G190), .A2(G200), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  OR2_X1    g0519(.A1(new_n719), .A2(KEYINPUT97), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(KEYINPUT97), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G329), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n401), .A2(G179), .A3(G200), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(new_n262), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G294), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n262), .A2(new_n301), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n401), .A2(new_n299), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(G326), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n299), .A2(G190), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n716), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(G283), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n320), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n729), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n738), .A2(new_n401), .A3(G200), .ZN(new_n739));
  AOI211_X1 g0539(.A(new_n733), .B(new_n737), .C1(G322), .C2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n730), .A2(new_n716), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n468), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n729), .A2(new_n734), .ZN(new_n743));
  INV_X1    g0543(.A(G317), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n744), .A2(KEYINPUT33), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(KEYINPUT33), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n743), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n729), .A2(new_n717), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI211_X1 g0549(.A(new_n742), .B(new_n747), .C1(G311), .C2(new_n749), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n724), .A2(new_n728), .A3(new_n740), .A4(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n735), .A2(new_n206), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n731), .A2(new_n364), .ZN(new_n753));
  AOI211_X1 g0553(.A(new_n752), .B(new_n753), .C1(G97), .C2(new_n727), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n285), .B1(new_n741), .B2(new_n330), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT96), .ZN(new_n756));
  INV_X1    g0556(.A(G159), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n718), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT32), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n222), .A2(new_n743), .B1(new_n748), .B2(new_n202), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n760), .B1(G58), .B2(new_n739), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n754), .A2(new_n756), .A3(new_n759), .A4(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n715), .B1(new_n751), .B2(new_n762), .ZN(new_n763));
  NOR4_X1   g0563(.A1(new_n714), .A2(new_n654), .A3(new_n695), .A4(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n705), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n764), .B1(new_n643), .B2(new_n765), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n698), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(G396));
  OAI211_X1 g0568(.A(new_n306), .B(new_n641), .C1(new_n631), .C2(new_n606), .ZN(new_n769));
  INV_X1    g0569(.A(new_n667), .ZN(new_n770));
  INV_X1    g0570(.A(new_n273), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n300), .B1(new_n771), .B2(new_n641), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(new_n305), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n305), .A2(new_n640), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n769), .B1(new_n770), .B2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n690), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n696), .B1(new_n778), .B2(new_n779), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n735), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n320), .B1(new_n783), .B2(G68), .ZN(new_n784));
  OAI221_X1 g0584(.A(new_n784), .B1(new_n364), .B2(new_n741), .C1(new_n221), .C2(new_n726), .ZN(new_n785));
  INV_X1    g0585(.A(new_n743), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n739), .A2(G143), .B1(G150), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(G137), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n787), .B1(new_n788), .B2(new_n731), .C1(new_n757), .C2(new_n748), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n789), .B(KEYINPUT34), .Z(new_n790));
  AOI211_X1 g0590(.A(new_n785), .B(new_n790), .C1(G132), .C2(new_n723), .ZN(new_n791));
  INV_X1    g0591(.A(G311), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n722), .A2(new_n792), .B1(new_n330), .B2(new_n735), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT99), .ZN(new_n794));
  AOI22_X1  g0594(.A1(G116), .A2(new_n749), .B1(new_n786), .B2(G283), .ZN(new_n795));
  INV_X1    g0595(.A(G294), .ZN(new_n796));
  INV_X1    g0596(.A(new_n739), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n795), .B1(new_n206), .B2(new_n741), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n320), .B1(new_n731), .B2(new_n468), .C1(new_n726), .C2(new_n205), .ZN(new_n799));
  NOR3_X1   g0599(.A1(new_n794), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n702), .B1(new_n791), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n702), .A2(new_n703), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n696), .B1(new_n803), .B2(G77), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT98), .Z(new_n805));
  OAI211_X1 g0605(.A(new_n801), .B(new_n805), .C1(new_n777), .C2(new_n704), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT100), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n782), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(G384));
  NOR2_X1   g0609(.A1(new_n220), .A2(new_n486), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT35), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n810), .B1(new_n515), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(new_n811), .B2(new_n515), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT36), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n310), .A2(new_n657), .A3(G77), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n364), .A2(G68), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n253), .B(G13), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  OR3_X1    g0618(.A1(new_n399), .A2(KEYINPUT102), .A3(new_n640), .ZN(new_n819));
  OAI21_X1  g0619(.A(KEYINPUT102), .B1(new_n399), .B2(new_n640), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT38), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT37), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n345), .A2(new_n340), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n638), .B1(new_n326), .B2(new_n337), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n823), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n827), .A2(new_n345), .A3(new_n823), .A4(new_n340), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n827), .B1(new_n350), .B2(new_n341), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n822), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT101), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n826), .B(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n587), .B2(new_n349), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n823), .B1(new_n835), .B2(new_n825), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n837), .B(KEYINPUT38), .C1(new_n838), .C2(new_n830), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT39), .ZN(new_n840));
  AND3_X1   g0640(.A1(new_n833), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n835), .A2(new_n825), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n830), .B1(new_n842), .B2(KEYINPUT37), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n835), .B1(new_n350), .B2(new_n341), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n822), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n840), .B1(new_n845), .B2(new_n839), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n821), .B1(new_n841), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n349), .A2(new_n638), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n397), .A2(new_n398), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n385), .A2(new_n640), .ZN(new_n851));
  MUX2_X1   g0651(.A(new_n850), .B(new_n403), .S(new_n851), .Z(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(new_n769), .B2(new_n775), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n845), .A2(new_n839), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n849), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n591), .B1(new_n668), .B2(new_n404), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n856), .B(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n852), .A2(new_n776), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n679), .A2(new_n680), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n689), .A2(new_n860), .ZN(new_n861));
  AND2_X1   g0661(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT40), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(new_n833), .B2(new_n839), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n859), .A2(new_n861), .A3(new_n854), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n862), .A2(new_n864), .B1(new_n865), .B2(new_n863), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n404), .A2(new_n861), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n669), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n867), .B2(new_n866), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n858), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n253), .B2(new_n693), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n858), .A2(new_n869), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n818), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n873), .B(KEYINPUT103), .ZN(G367));
  NAND2_X1  g0674(.A1(new_n619), .A2(new_n640), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n537), .B(new_n543), .C1(new_n541), .C2(new_n641), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n465), .A2(new_n651), .A3(new_n877), .ZN(new_n878));
  OR2_X1    g0678(.A1(new_n878), .A2(KEYINPUT42), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n877), .A2(new_n452), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n640), .B1(new_n880), .B2(new_n537), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n881), .B1(new_n878), .B2(KEYINPUT42), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n641), .B1(new_n571), .B2(new_n573), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n623), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n610), .A2(new_n884), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT43), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n888), .A2(KEYINPUT43), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n883), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n879), .A2(new_n882), .A3(new_n890), .A4(new_n889), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n877), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n649), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n895), .B(new_n897), .ZN(new_n898));
  XOR2_X1   g0698(.A(new_n654), .B(KEYINPUT41), .Z(new_n899));
  INV_X1    g0699(.A(new_n649), .ZN(new_n900));
  AND3_X1   g0700(.A1(new_n652), .A2(KEYINPUT45), .A3(new_n877), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT45), .B1(new_n652), .B2(new_n877), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n465), .A2(new_n651), .ZN(new_n904));
  INV_X1    g0704(.A(new_n650), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT44), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n906), .A2(new_n907), .A3(new_n896), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT44), .B1(new_n652), .B2(new_n877), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n900), .B1(new_n903), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n904), .B1(new_n648), .B2(new_n651), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n645), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n644), .B(new_n904), .C1(new_n648), .C2(new_n651), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n904), .A2(new_n905), .A3(new_n877), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT45), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n652), .A2(KEYINPUT45), .A3(new_n877), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n920), .A2(new_n649), .A3(new_n909), .A4(new_n908), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n911), .A2(new_n915), .A3(new_n921), .A4(new_n691), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n899), .B1(new_n922), .B2(new_n691), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n898), .B1(new_n923), .B2(new_n695), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(KEYINPUT104), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT104), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n898), .B(new_n926), .C1(new_n923), .C2(new_n695), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n889), .A2(new_n705), .ZN(new_n929));
  INV_X1    g0729(.A(new_n243), .ZN(new_n930));
  OAI221_X1 g0730(.A(new_n706), .B1(new_n212), .B2(new_n269), .C1(new_n930), .C2(new_n711), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n696), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n735), .A2(new_n202), .ZN(new_n933));
  INV_X1    g0733(.A(G150), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n285), .B1(new_n797), .B2(new_n934), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n933), .B(new_n935), .C1(G137), .C2(new_n719), .ZN(new_n936));
  INV_X1    g0736(.A(new_n741), .ZN(new_n937));
  AOI22_X1  g0737(.A1(G50), .A2(new_n749), .B1(new_n937), .B2(G58), .ZN(new_n938));
  INV_X1    g0738(.A(new_n731), .ZN(new_n939));
  AOI22_X1  g0739(.A1(G143), .A2(new_n939), .B1(new_n786), .B2(G159), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n727), .A2(G68), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n936), .A2(new_n938), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  OAI221_X1 g0742(.A(new_n320), .B1(new_n718), .B2(new_n744), .C1(new_n205), .C2(new_n735), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT106), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n937), .A2(KEYINPUT46), .A3(G116), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT105), .Z(new_n946));
  AOI22_X1  g0746(.A1(G311), .A2(new_n939), .B1(new_n749), .B2(G283), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n739), .A2(G303), .B1(G294), .B2(new_n786), .ZN(new_n948));
  AOI21_X1  g0748(.A(KEYINPUT46), .B1(new_n937), .B2(G116), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(G107), .B2(new_n727), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n946), .A2(new_n947), .A3(new_n948), .A4(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n942), .B1(new_n944), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT47), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n715), .B1(new_n952), .B2(new_n953), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n932), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n929), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n928), .A2(new_n957), .ZN(G387));
  AOI22_X1  g0758(.A1(G322), .A2(new_n939), .B1(new_n749), .B2(G303), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n959), .B1(new_n792), .B2(new_n743), .C1(new_n744), .C2(new_n797), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT48), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n960), .A2(new_n961), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n727), .A2(G283), .B1(new_n937), .B2(G294), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT49), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(new_n966), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n320), .B1(new_n718), .B2(new_n732), .C1(new_n486), .C2(new_n735), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT107), .Z(new_n970));
  NAND3_X1  g0770(.A1(new_n967), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n741), .A2(new_n202), .B1(new_n718), .B2(new_n934), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n726), .A2(new_n269), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n285), .B1(new_n735), .B2(new_n205), .ZN(new_n974));
  NOR3_X1   g0774(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n739), .A2(G50), .B1(G68), .B2(new_n749), .ZN(new_n976));
  AOI22_X1  g0776(.A1(G159), .A2(new_n939), .B1(new_n786), .B2(new_n336), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n715), .B1(new_n971), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n709), .A2(new_n655), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(G107), .B2(new_n212), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n240), .A2(G45), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n267), .A2(G50), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT50), .ZN(new_n984));
  AOI211_X1 g0784(.A(G45), .B(new_n655), .C1(G68), .C2(G77), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n711), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n981), .B1(new_n982), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n696), .B1(new_n987), .B2(new_n707), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n979), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n648), .B2(new_n765), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n990), .B(KEYINPUT108), .Z(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(new_n695), .B2(new_n915), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n915), .A2(new_n691), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n915), .A2(new_n691), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n654), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n992), .B1(new_n993), .B2(new_n995), .ZN(G393));
  NAND2_X1  g0796(.A1(new_n911), .A2(new_n921), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n997), .A2(new_n694), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n896), .A2(new_n705), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n706), .B1(new_n205), .B2(new_n212), .C1(new_n251), .C2(new_n711), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n696), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n726), .A2(new_n202), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n320), .B(new_n1002), .C1(G87), .C2(new_n783), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(G50), .A2(new_n786), .B1(new_n937), .B2(G68), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n336), .A2(new_n749), .B1(new_n719), .B2(G143), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n739), .A2(G159), .B1(new_n939), .B2(G150), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT51), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n739), .A2(G311), .B1(new_n939), .B2(G317), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT52), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n285), .B(new_n752), .C1(G116), .C2(new_n727), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(G283), .A2(new_n937), .B1(new_n719), .B2(G322), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(G294), .A2(new_n749), .B1(new_n786), .B2(G303), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n1006), .A2(new_n1008), .B1(new_n1010), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1001), .B1(new_n1015), .B2(new_n702), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n998), .B1(new_n999), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n997), .A2(new_n994), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1018), .A2(new_n654), .A3(new_n922), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1019), .ZN(G390));
  NAND2_X1  g0820(.A1(new_n667), .A2(new_n665), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n666), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1021), .A2(new_n404), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n669), .B1(new_n689), .B2(new_n860), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n404), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1023), .A2(new_n592), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT111), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1024), .A2(new_n777), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n852), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n852), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n690), .A2(new_n777), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n664), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n774), .B1(new_n1033), .B2(new_n773), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1030), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n688), .A2(new_n689), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1036), .A2(G330), .A3(new_n777), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n1037), .A2(new_n852), .B1(new_n859), .B2(new_n1024), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n769), .A2(new_n775), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1035), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n857), .A2(KEYINPUT111), .A3(new_n1025), .ZN(new_n1042));
  AND3_X1   g0842(.A1(new_n1028), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n841), .A2(new_n846), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n853), .B2(new_n821), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1024), .A2(new_n859), .A3(KEYINPUT110), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1046), .A2(new_n690), .A3(new_n777), .A4(new_n1031), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT109), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n821), .B(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n833), .A2(new_n839), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(new_n852), .C2(new_n1034), .ZN(new_n1051));
  AND3_X1   g0851(.A1(new_n1045), .A2(new_n1047), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1024), .A2(new_n859), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1053), .A2(KEYINPUT110), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n1045), .B2(new_n1051), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(KEYINPUT112), .B1(new_n1043), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n654), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n1043), .B2(new_n1056), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1045), .A2(new_n1047), .A3(new_n1051), .ZN(new_n1060));
  AND2_X1   g0860(.A1(new_n1045), .A2(new_n1051), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1060), .B1(new_n1061), .B2(new_n1054), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT112), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1028), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1057), .A2(new_n1059), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(G125), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT114), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n285), .B1(new_n735), .B2(new_n364), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n722), .A2(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT115), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n937), .A2(G150), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT53), .ZN(new_n1074));
  INV_X1    g0874(.A(G132), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n797), .A2(new_n1075), .B1(new_n743), .B2(new_n788), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n726), .A2(new_n757), .ZN(new_n1077));
  INV_X1    g0877(.A(G128), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(KEYINPUT54), .B(G143), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n731), .A2(new_n1078), .B1(new_n748), .B2(new_n1079), .ZN(new_n1080));
  OR3_X1    g0880(.A1(new_n1076), .A2(new_n1077), .A3(new_n1080), .ZN(new_n1081));
  NOR3_X1   g0881(.A1(new_n1072), .A2(new_n1074), .A3(new_n1081), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(G283), .A2(new_n939), .B1(new_n786), .B2(G107), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n1083), .B1(new_n205), .B2(new_n748), .C1(new_n722), .C2(new_n796), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n285), .B1(new_n937), .B2(G87), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1085), .B1(new_n222), .B2(new_n735), .C1(new_n797), .C2(new_n486), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n1084), .A2(new_n1002), .A3(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n702), .B1(new_n1082), .B2(new_n1087), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1088), .B(new_n696), .C1(new_n336), .C2(new_n803), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n1044), .B2(new_n703), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n695), .B(new_n1060), .C1(new_n1061), .C2(new_n1054), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(KEYINPUT113), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT113), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1056), .A2(new_n1093), .A3(new_n695), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1090), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1066), .A2(new_n1095), .ZN(G378));
  INV_X1    g0896(.A(KEYINPUT57), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1028), .A2(new_n1042), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n1056), .B2(new_n1041), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n374), .B(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n638), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n366), .A2(new_n1102), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1101), .B(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n866), .A2(G330), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n865), .A2(new_n863), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n859), .A2(new_n864), .A3(new_n861), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1106), .A2(G330), .A3(new_n1107), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1101), .B(new_n1103), .Z(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  AND3_X1   g0910(.A1(new_n856), .A2(new_n1105), .A3(new_n1110), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n1105), .A2(new_n1110), .B1(new_n855), .B2(new_n849), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1097), .B1(new_n1099), .B2(new_n1113), .ZN(new_n1114));
  OR2_X1    g0914(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1098), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1115), .A2(new_n1117), .A3(KEYINPUT57), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1114), .A2(new_n1118), .A3(new_n654), .ZN(new_n1119));
  AOI211_X1 g0919(.A(G41), .B(new_n285), .C1(new_n937), .C2(G77), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1120), .B1(new_n221), .B2(new_n735), .C1(new_n722), .C2(new_n736), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n1121), .B(KEYINPUT116), .Z(new_n1122));
  NOR2_X1   g0922(.A1(new_n743), .A2(new_n205), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n731), .A2(new_n486), .B1(new_n748), .B2(new_n269), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n1123), .B(new_n1124), .C1(G107), .C2(new_n739), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1122), .A2(new_n941), .A3(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT58), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n364), .B1(new_n318), .B2(G41), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n797), .A2(new_n1078), .B1(new_n741), .B2(new_n1079), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(G125), .A2(new_n939), .B1(new_n749), .B2(G137), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n1075), .B2(new_n743), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n1129), .B(new_n1131), .C1(G150), .C2(new_n727), .ZN(new_n1132));
  XOR2_X1   g0932(.A(new_n1132), .B(KEYINPUT117), .Z(new_n1133));
  NOR2_X1   g0933(.A1(new_n1133), .A2(KEYINPUT59), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(KEYINPUT59), .ZN(new_n1135));
  AOI211_X1 g0935(.A(G33), .B(G41), .C1(new_n783), .C2(G159), .ZN(new_n1136));
  INV_X1    g0936(.A(G124), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1136), .B1(new_n1137), .B2(new_n718), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT118), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1135), .A2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1127), .B(new_n1128), .C1(new_n1134), .C2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT119), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n715), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(new_n1142), .B2(new_n1141), .ZN(new_n1144));
  XOR2_X1   g0944(.A(new_n1144), .B(KEYINPUT120), .Z(new_n1145));
  OAI21_X1  g0945(.A(new_n696), .B1(new_n803), .B2(G50), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1109), .A2(new_n703), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n1113), .B2(new_n694), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1119), .A2(new_n1151), .ZN(G375));
  NAND2_X1  g0952(.A1(new_n1037), .A2(new_n852), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n1053), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1034), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(new_n1029), .B2(new_n852), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n1154), .A2(new_n1039), .B1(new_n1156), .B2(new_n1032), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1158));
  AOI21_X1  g0958(.A(KEYINPUT111), .B1(new_n857), .B2(new_n1025), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1157), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT121), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n899), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1098), .A2(KEYINPUT121), .A3(new_n1157), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1162), .A2(new_n1163), .A3(new_n1064), .A4(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n285), .B1(new_n735), .B2(new_n221), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n731), .A2(new_n1075), .B1(new_n741), .B2(new_n757), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1166), .B(new_n1167), .C1(G50), .C2(new_n727), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n749), .A2(G150), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1169), .B1(new_n743), .B2(new_n1079), .C1(new_n797), .C2(new_n788), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(G128), .B2(new_n723), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n739), .A2(G283), .B1(new_n939), .B2(G294), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n206), .B2(new_n748), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(G303), .B2(new_n723), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n205), .A2(new_n741), .B1(new_n743), .B2(new_n486), .ZN(new_n1175));
  NOR4_X1   g0975(.A1(new_n1175), .A2(new_n973), .A3(new_n285), .A4(new_n933), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n1168), .A2(new_n1171), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n696), .B1(G68), .B2(new_n803), .C1(new_n1177), .C2(new_n715), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n852), .B2(new_n703), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n1041), .B2(new_n695), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1165), .A2(new_n1180), .ZN(G381));
  OR4_X1    g0981(.A1(G396), .A2(G381), .A3(G384), .A4(G393), .ZN(new_n1182));
  INV_X1    g0982(.A(G390), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n928), .A2(new_n957), .A3(new_n1183), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n1182), .A2(G375), .A3(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT122), .ZN(new_n1186));
  AND3_X1   g0986(.A1(new_n1066), .A2(new_n1095), .A3(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1186), .B1(new_n1066), .B2(new_n1095), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1185), .A2(new_n1189), .ZN(G407));
  NAND2_X1  g0990(.A1(new_n639), .A2(G213), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT123), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1189), .A2(new_n1151), .A3(new_n1119), .A4(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(G407), .A2(G213), .A3(new_n1193), .ZN(G409));
  XNOR2_X1  g0994(.A(G393), .B(new_n767), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n928), .A2(new_n957), .A3(new_n1183), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1183), .B1(new_n928), .B2(new_n957), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1195), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(G387), .A2(G390), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1195), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1199), .A2(new_n1184), .A3(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1198), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1064), .A2(KEYINPUT60), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1162), .A2(new_n1164), .A3(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT124), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1041), .B1(new_n1028), .B2(new_n1042), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1058), .B1(new_n1206), .B2(KEYINPUT60), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n1204), .A2(new_n1205), .A3(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1205), .B1(new_n1204), .B2(new_n1207), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1180), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n808), .ZN(new_n1211));
  OAI211_X1 g1011(.A(G384), .B(new_n1180), .C1(new_n1208), .C2(new_n1209), .ZN(new_n1212));
  AND3_X1   g1012(.A1(new_n1211), .A2(KEYINPUT63), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(G378), .A2(KEYINPUT122), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1066), .A2(new_n1095), .A3(new_n1186), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1099), .A2(new_n1113), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n1163), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n1151), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1214), .A2(new_n1215), .A3(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1119), .A2(G378), .A3(new_n1151), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1192), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1202), .B1(new_n1213), .B2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT63), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1192), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1150), .B1(new_n1216), .B2(new_n1163), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1187), .A2(new_n1188), .A3(new_n1225), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n1119), .A2(G378), .A3(new_n1151), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1224), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1223), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1192), .A2(G2897), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1204), .A2(new_n1207), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(KEYINPUT124), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1204), .A2(new_n1205), .A3(new_n1207), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(G384), .B1(new_n1236), .B2(new_n1180), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1212), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1232), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1211), .A2(new_n1212), .A3(new_n1231), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1239), .A2(new_n1228), .A3(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT61), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1222), .A2(new_n1230), .A3(new_n1241), .A4(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT125), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(KEYINPUT62), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT62), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1247), .A2(new_n1221), .A3(new_n1248), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1246), .A2(new_n1241), .A3(new_n1242), .A4(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n1202), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n1198), .A2(new_n1201), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1211), .A2(KEYINPUT63), .A3(new_n1212), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1252), .B1(new_n1228), .B2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(KEYINPUT63), .B1(new_n1247), .B2(new_n1221), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1231), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1257), .A2(new_n1221), .ZN(new_n1258));
  AOI21_X1  g1058(.A(KEYINPUT61), .B1(new_n1258), .B2(new_n1240), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1256), .A2(new_n1259), .A3(KEYINPUT125), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1245), .A2(new_n1251), .A3(new_n1260), .ZN(G405));
  INV_X1    g1061(.A(KEYINPUT127), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1229), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1189), .A2(G375), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1227), .B1(new_n1264), .B2(KEYINPUT126), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1265), .B1(KEYINPUT126), .B2(new_n1264), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1247), .A2(KEYINPUT127), .A3(new_n1202), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1252), .B1(new_n1262), .B2(new_n1229), .ZN(new_n1268));
  AND4_X1   g1068(.A1(new_n1263), .A2(new_n1266), .A3(new_n1267), .A4(new_n1268), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n1266), .A2(new_n1263), .B1(new_n1268), .B2(new_n1267), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1269), .A2(new_n1270), .ZN(G402));
endmodule


