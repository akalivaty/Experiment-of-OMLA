

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584;

  NOR2_X1 U323 ( .A1(n479), .A2(n578), .ZN(n480) );
  XNOR2_X1 U324 ( .A(n347), .B(n346), .ZN(n352) );
  XNOR2_X1 U325 ( .A(n345), .B(n344), .ZN(n346) );
  INV_X1 U326 ( .A(G71GAT), .ZN(n447) );
  XNOR2_X1 U327 ( .A(KEYINPUT106), .B(KEYINPUT38), .ZN(n481) );
  XOR2_X1 U328 ( .A(KEYINPUT37), .B(KEYINPUT105), .Z(n291) );
  INV_X1 U329 ( .A(KEYINPUT46), .ZN(n358) );
  AND2_X1 U330 ( .A1(n379), .A2(n378), .ZN(n380) );
  XNOR2_X1 U331 ( .A(n382), .B(KEYINPUT113), .ZN(n383) );
  NOR2_X1 U332 ( .A1(n470), .A2(n469), .ZN(n471) );
  XNOR2_X1 U333 ( .A(n293), .B(KEYINPUT33), .ZN(n294) );
  XNOR2_X1 U334 ( .A(n367), .B(n294), .ZN(n298) );
  XNOR2_X1 U335 ( .A(KEYINPUT26), .B(KEYINPUT98), .ZN(n461) );
  XNOR2_X1 U336 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U337 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U338 ( .A(n462), .B(n461), .ZN(n570) );
  XNOR2_X1 U339 ( .A(n304), .B(n303), .ZN(n388) );
  XNOR2_X1 U340 ( .A(n450), .B(n449), .ZN(n453) );
  XNOR2_X1 U341 ( .A(n357), .B(n356), .ZN(n572) );
  XNOR2_X1 U342 ( .A(n482), .B(n481), .ZN(n507) );
  XNOR2_X1 U343 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U344 ( .A(n483), .B(G43GAT), .ZN(n484) );
  XNOR2_X1 U345 ( .A(n489), .B(n488), .ZN(G1351GAT) );
  XNOR2_X1 U346 ( .A(n485), .B(n484), .ZN(G1330GAT) );
  XNOR2_X1 U347 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n292) );
  XNOR2_X1 U348 ( .A(n292), .B(KEYINPUT72), .ZN(n367) );
  AND2_X1 U349 ( .A1(G230GAT), .A2(G233GAT), .ZN(n293) );
  XOR2_X1 U350 ( .A(KEYINPUT73), .B(KEYINPUT31), .Z(n296) );
  XNOR2_X1 U351 ( .A(G204GAT), .B(KEYINPUT32), .ZN(n295) );
  XOR2_X1 U352 ( .A(n296), .B(n295), .Z(n297) );
  XNOR2_X1 U353 ( .A(n298), .B(n297), .ZN(n304) );
  XNOR2_X1 U354 ( .A(G120GAT), .B(G148GAT), .ZN(n299) );
  XNOR2_X1 U355 ( .A(n299), .B(G57GAT), .ZN(n424) );
  XNOR2_X1 U356 ( .A(G176GAT), .B(G92GAT), .ZN(n300) );
  XNOR2_X1 U357 ( .A(n300), .B(G64GAT), .ZN(n311) );
  XNOR2_X1 U358 ( .A(n424), .B(n311), .ZN(n302) );
  XOR2_X1 U359 ( .A(G106GAT), .B(G78GAT), .Z(n398) );
  XOR2_X1 U360 ( .A(G99GAT), .B(G85GAT), .Z(n329) );
  XNOR2_X1 U361 ( .A(n398), .B(n329), .ZN(n301) );
  XOR2_X1 U362 ( .A(KEYINPUT41), .B(n388), .Z(n554) );
  XNOR2_X1 U363 ( .A(G211GAT), .B(G218GAT), .ZN(n305) );
  XNOR2_X1 U364 ( .A(n305), .B(KEYINPUT21), .ZN(n306) );
  XOR2_X1 U365 ( .A(n306), .B(KEYINPUT87), .Z(n308) );
  XNOR2_X1 U366 ( .A(G197GAT), .B(G204GAT), .ZN(n307) );
  XNOR2_X1 U367 ( .A(n308), .B(n307), .ZN(n402) );
  XOR2_X1 U368 ( .A(G169GAT), .B(G8GAT), .Z(n343) );
  XOR2_X1 U369 ( .A(KEYINPUT97), .B(n343), .Z(n310) );
  NAND2_X1 U370 ( .A1(G226GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U371 ( .A(n310), .B(n309), .ZN(n312) );
  XOR2_X1 U372 ( .A(n312), .B(n311), .Z(n317) );
  XOR2_X1 U373 ( .A(G183GAT), .B(KEYINPUT17), .Z(n314) );
  XNOR2_X1 U374 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n313) );
  XNOR2_X1 U375 ( .A(n314), .B(n313), .ZN(n439) );
  XNOR2_X1 U376 ( .A(G36GAT), .B(G190GAT), .ZN(n315) );
  XNOR2_X1 U377 ( .A(n315), .B(KEYINPUT78), .ZN(n323) );
  XNOR2_X1 U378 ( .A(n439), .B(n323), .ZN(n316) );
  XNOR2_X1 U379 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U380 ( .A(n402), .B(n318), .ZN(n505) );
  XOR2_X1 U381 ( .A(KEYINPUT75), .B(KEYINPUT76), .Z(n320) );
  NAND2_X1 U382 ( .A1(G232GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U383 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U384 ( .A(n321), .B(KEYINPUT64), .Z(n325) );
  XNOR2_X1 U385 ( .A(G29GAT), .B(G134GAT), .ZN(n322) );
  XNOR2_X1 U386 ( .A(n322), .B(KEYINPUT77), .ZN(n429) );
  XNOR2_X1 U387 ( .A(n429), .B(n323), .ZN(n324) );
  XNOR2_X1 U388 ( .A(n325), .B(n324), .ZN(n333) );
  XOR2_X1 U389 ( .A(G92GAT), .B(KEYINPUT11), .Z(n327) );
  XNOR2_X1 U390 ( .A(G106GAT), .B(KEYINPUT9), .ZN(n326) );
  XNOR2_X1 U391 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U392 ( .A(n328), .B(KEYINPUT10), .Z(n331) );
  XNOR2_X1 U393 ( .A(G218GAT), .B(n329), .ZN(n330) );
  XNOR2_X1 U394 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U395 ( .A(n333), .B(n332), .Z(n337) );
  XNOR2_X1 U396 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n334) );
  XNOR2_X1 U397 ( .A(n334), .B(KEYINPUT7), .ZN(n350) );
  XNOR2_X1 U398 ( .A(G50GAT), .B(KEYINPUT74), .ZN(n335) );
  XNOR2_X1 U399 ( .A(n335), .B(G162GAT), .ZN(n408) );
  XNOR2_X1 U400 ( .A(n350), .B(n408), .ZN(n336) );
  XNOR2_X1 U401 ( .A(n337), .B(n336), .ZN(n561) );
  XOR2_X1 U402 ( .A(G113GAT), .B(G197GAT), .Z(n339) );
  XNOR2_X1 U403 ( .A(G50GAT), .B(G141GAT), .ZN(n338) );
  XNOR2_X1 U404 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U405 ( .A(n340), .B(G36GAT), .Z(n347) );
  XOR2_X1 U406 ( .A(KEYINPUT67), .B(KEYINPUT68), .Z(n342) );
  XNOR2_X1 U407 ( .A(KEYINPUT71), .B(KEYINPUT69), .ZN(n341) );
  XOR2_X1 U408 ( .A(n342), .B(n341), .Z(n345) );
  XNOR2_X1 U409 ( .A(n343), .B(G29GAT), .ZN(n344) );
  XOR2_X1 U410 ( .A(G1GAT), .B(KEYINPUT70), .Z(n349) );
  XNOR2_X1 U411 ( .A(G22GAT), .B(G15GAT), .ZN(n348) );
  XNOR2_X1 U412 ( .A(n349), .B(n348), .ZN(n369) );
  XNOR2_X1 U413 ( .A(n350), .B(n369), .ZN(n351) );
  XNOR2_X1 U414 ( .A(n352), .B(n351), .ZN(n357) );
  XOR2_X1 U415 ( .A(KEYINPUT66), .B(KEYINPUT29), .Z(n354) );
  NAND2_X1 U416 ( .A1(G229GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U417 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U418 ( .A(KEYINPUT30), .B(n355), .Z(n356) );
  AND2_X1 U419 ( .A1(n572), .A2(n554), .ZN(n359) );
  XNOR2_X1 U420 ( .A(n359), .B(n358), .ZN(n379) );
  XOR2_X1 U421 ( .A(KEYINPUT15), .B(KEYINPUT80), .Z(n361) );
  XNOR2_X1 U422 ( .A(KEYINPUT81), .B(KEYINPUT12), .ZN(n360) );
  XNOR2_X1 U423 ( .A(n361), .B(n360), .ZN(n377) );
  XOR2_X1 U424 ( .A(G64GAT), .B(G211GAT), .Z(n363) );
  XNOR2_X1 U425 ( .A(G127GAT), .B(G183GAT), .ZN(n362) );
  XNOR2_X1 U426 ( .A(n363), .B(n362), .ZN(n365) );
  XOR2_X1 U427 ( .A(G155GAT), .B(G78GAT), .Z(n364) );
  XNOR2_X1 U428 ( .A(n365), .B(n364), .ZN(n373) );
  XNOR2_X1 U429 ( .A(G57GAT), .B(KEYINPUT14), .ZN(n366) );
  XNOR2_X1 U430 ( .A(n366), .B(KEYINPUT79), .ZN(n368) );
  XOR2_X1 U431 ( .A(n368), .B(n367), .Z(n371) );
  XNOR2_X1 U432 ( .A(n369), .B(G8GAT), .ZN(n370) );
  XNOR2_X1 U433 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U434 ( .A(n373), .B(n372), .ZN(n375) );
  NAND2_X1 U435 ( .A1(G231GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U436 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U437 ( .A(n377), .B(n376), .ZN(n578) );
  INV_X1 U438 ( .A(n578), .ZN(n378) );
  XOR2_X1 U439 ( .A(KEYINPUT112), .B(n380), .Z(n381) );
  NOR2_X1 U440 ( .A1(n561), .A2(n381), .ZN(n384) );
  INV_X1 U441 ( .A(KEYINPUT47), .ZN(n382) );
  XNOR2_X1 U442 ( .A(n384), .B(n383), .ZN(n392) );
  XNOR2_X1 U443 ( .A(KEYINPUT36), .B(KEYINPUT104), .ZN(n385) );
  XNOR2_X1 U444 ( .A(n561), .B(n385), .ZN(n581) );
  NAND2_X1 U445 ( .A1(n581), .A2(n578), .ZN(n387) );
  XOR2_X1 U446 ( .A(KEYINPUT45), .B(KEYINPUT114), .Z(n386) );
  XNOR2_X1 U447 ( .A(n387), .B(n386), .ZN(n389) );
  INV_X1 U448 ( .A(n388), .ZN(n460) );
  NAND2_X1 U449 ( .A1(n389), .A2(n460), .ZN(n390) );
  OR2_X1 U450 ( .A1(n572), .A2(n390), .ZN(n391) );
  AND2_X1 U451 ( .A1(n392), .A2(n391), .ZN(n393) );
  XNOR2_X1 U452 ( .A(n393), .B(KEYINPUT48), .ZN(n534) );
  NOR2_X1 U453 ( .A1(n505), .A2(n534), .ZN(n394) );
  XNOR2_X1 U454 ( .A(n394), .B(KEYINPUT54), .ZN(n568) );
  XOR2_X1 U455 ( .A(KEYINPUT86), .B(KEYINPUT22), .Z(n396) );
  XNOR2_X1 U456 ( .A(KEYINPUT24), .B(G148GAT), .ZN(n395) );
  XNOR2_X1 U457 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U458 ( .A(n397), .B(KEYINPUT88), .Z(n400) );
  XNOR2_X1 U459 ( .A(G22GAT), .B(n398), .ZN(n399) );
  XNOR2_X1 U460 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U461 ( .A(n402), .B(n401), .ZN(n412) );
  XOR2_X1 U462 ( .A(KEYINPUT85), .B(KEYINPUT89), .Z(n404) );
  NAND2_X1 U463 ( .A1(G228GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U464 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U465 ( .A(n405), .B(KEYINPUT23), .Z(n410) );
  XOR2_X1 U466 ( .A(G155GAT), .B(KEYINPUT2), .Z(n407) );
  XNOR2_X1 U467 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n406) );
  XNOR2_X1 U468 ( .A(n407), .B(n406), .ZN(n421) );
  XNOR2_X1 U469 ( .A(n408), .B(n421), .ZN(n409) );
  XNOR2_X1 U470 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U471 ( .A(n412), .B(n411), .ZN(n472) );
  XOR2_X1 U472 ( .A(KEYINPUT90), .B(KEYINPUT94), .Z(n414) );
  XNOR2_X1 U473 ( .A(KEYINPUT1), .B(KEYINPUT5), .ZN(n413) );
  XNOR2_X1 U474 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U475 ( .A(KEYINPUT91), .B(KEYINPUT6), .Z(n416) );
  XNOR2_X1 U476 ( .A(KEYINPUT92), .B(KEYINPUT4), .ZN(n415) );
  XNOR2_X1 U477 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U478 ( .A(n418), .B(n417), .Z(n423) );
  XOR2_X1 U479 ( .A(G127GAT), .B(KEYINPUT82), .Z(n420) );
  XNOR2_X1 U480 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n419) );
  XNOR2_X1 U481 ( .A(n420), .B(n419), .ZN(n451) );
  XNOR2_X1 U482 ( .A(n451), .B(n421), .ZN(n422) );
  XNOR2_X1 U483 ( .A(n423), .B(n422), .ZN(n428) );
  XOR2_X1 U484 ( .A(G85GAT), .B(KEYINPUT95), .Z(n426) );
  XNOR2_X1 U485 ( .A(G162GAT), .B(n424), .ZN(n425) );
  XNOR2_X1 U486 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U487 ( .A(n428), .B(n427), .Z(n434) );
  XOR2_X1 U488 ( .A(n429), .B(KEYINPUT93), .Z(n431) );
  NAND2_X1 U489 ( .A1(G225GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U490 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U491 ( .A(G1GAT), .B(n432), .ZN(n433) );
  XNOR2_X1 U492 ( .A(n434), .B(n433), .ZN(n470) );
  XOR2_X1 U493 ( .A(KEYINPUT96), .B(n470), .Z(n569) );
  INV_X1 U494 ( .A(n569), .ZN(n523) );
  NOR2_X1 U495 ( .A1(n472), .A2(n523), .ZN(n435) );
  AND2_X1 U496 ( .A1(n568), .A2(n435), .ZN(n436) );
  XNOR2_X1 U497 ( .A(n436), .B(KEYINPUT55), .ZN(n454) );
  XOR2_X1 U498 ( .A(G190GAT), .B(G134GAT), .Z(n438) );
  NAND2_X1 U499 ( .A1(G227GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U500 ( .A(n438), .B(n437), .ZN(n440) );
  XOR2_X1 U501 ( .A(n440), .B(n439), .Z(n450) );
  XOR2_X1 U502 ( .A(KEYINPUT84), .B(KEYINPUT83), .Z(n442) );
  XNOR2_X1 U503 ( .A(G43GAT), .B(G99GAT), .ZN(n441) );
  XNOR2_X1 U504 ( .A(n442), .B(n441), .ZN(n446) );
  XOR2_X1 U505 ( .A(KEYINPUT20), .B(G176GAT), .Z(n444) );
  XNOR2_X1 U506 ( .A(G169GAT), .B(G15GAT), .ZN(n443) );
  XNOR2_X1 U507 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U508 ( .A(n446), .B(n445), .ZN(n448) );
  XNOR2_X1 U509 ( .A(n451), .B(G120GAT), .ZN(n452) );
  XNOR2_X1 U510 ( .A(n453), .B(n452), .ZN(n497) );
  NOR2_X1 U511 ( .A1(n454), .A2(n497), .ZN(n455) );
  XNOR2_X1 U512 ( .A(KEYINPUT122), .B(n455), .ZN(n566) );
  NAND2_X1 U513 ( .A1(n554), .A2(n566), .ZN(n459) );
  XOR2_X1 U514 ( .A(G176GAT), .B(KEYINPUT56), .Z(n457) );
  XNOR2_X1 U515 ( .A(KEYINPUT124), .B(KEYINPUT57), .ZN(n456) );
  XNOR2_X1 U516 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U517 ( .A(n459), .B(n458), .ZN(G1349GAT) );
  NAND2_X1 U518 ( .A1(n572), .A2(n460), .ZN(n493) );
  NAND2_X1 U519 ( .A1(n472), .A2(n497), .ZN(n462) );
  INV_X1 U520 ( .A(n570), .ZN(n550) );
  XOR2_X1 U521 ( .A(KEYINPUT27), .B(n505), .Z(n474) );
  NAND2_X1 U522 ( .A1(n550), .A2(n474), .ZN(n463) );
  XNOR2_X1 U523 ( .A(KEYINPUT99), .B(n463), .ZN(n468) );
  NOR2_X1 U524 ( .A1(n497), .A2(n505), .ZN(n464) );
  NOR2_X1 U525 ( .A1(n472), .A2(n464), .ZN(n465) );
  XOR2_X1 U526 ( .A(KEYINPUT100), .B(n465), .Z(n466) );
  XNOR2_X1 U527 ( .A(KEYINPUT25), .B(n466), .ZN(n467) );
  NOR2_X1 U528 ( .A1(n468), .A2(n467), .ZN(n469) );
  XNOR2_X1 U529 ( .A(n471), .B(KEYINPUT101), .ZN(n477) );
  XOR2_X1 U530 ( .A(n472), .B(KEYINPUT65), .Z(n473) );
  XNOR2_X1 U531 ( .A(KEYINPUT28), .B(n473), .ZN(n538) );
  NAND2_X1 U532 ( .A1(n523), .A2(n474), .ZN(n533) );
  NOR2_X1 U533 ( .A1(n538), .A2(n533), .ZN(n475) );
  NAND2_X1 U534 ( .A1(n475), .A2(n497), .ZN(n476) );
  NAND2_X1 U535 ( .A1(n477), .A2(n476), .ZN(n478) );
  XNOR2_X1 U536 ( .A(KEYINPUT102), .B(n478), .ZN(n491) );
  NAND2_X1 U537 ( .A1(n581), .A2(n491), .ZN(n479) );
  XNOR2_X1 U538 ( .A(n480), .B(n291), .ZN(n522) );
  OR2_X1 U539 ( .A1(n493), .A2(n522), .ZN(n482) );
  NOR2_X1 U540 ( .A1(n497), .A2(n507), .ZN(n485) );
  XNOR2_X1 U541 ( .A(KEYINPUT40), .B(KEYINPUT107), .ZN(n483) );
  NAND2_X1 U542 ( .A1(n561), .A2(n566), .ZN(n489) );
  XOR2_X1 U543 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n487) );
  XNOR2_X1 U544 ( .A(G190GAT), .B(KEYINPUT125), .ZN(n486) );
  NOR2_X1 U545 ( .A1(n561), .A2(n378), .ZN(n490) );
  XNOR2_X1 U546 ( .A(KEYINPUT16), .B(n490), .ZN(n492) );
  NAND2_X1 U547 ( .A1(n492), .A2(n491), .ZN(n511) );
  NOR2_X1 U548 ( .A1(n493), .A2(n511), .ZN(n500) );
  NAND2_X1 U549 ( .A1(n500), .A2(n523), .ZN(n494) );
  XNOR2_X1 U550 ( .A(KEYINPUT34), .B(n494), .ZN(n495) );
  XNOR2_X1 U551 ( .A(G1GAT), .B(n495), .ZN(G1324GAT) );
  INV_X1 U552 ( .A(n505), .ZN(n525) );
  NAND2_X1 U553 ( .A1(n500), .A2(n525), .ZN(n496) );
  XNOR2_X1 U554 ( .A(n496), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U555 ( .A(G15GAT), .B(KEYINPUT35), .Z(n499) );
  INV_X1 U556 ( .A(n497), .ZN(n535) );
  NAND2_X1 U557 ( .A1(n500), .A2(n535), .ZN(n498) );
  XNOR2_X1 U558 ( .A(n499), .B(n498), .ZN(G1326GAT) );
  XOR2_X1 U559 ( .A(G22GAT), .B(KEYINPUT103), .Z(n502) );
  NAND2_X1 U560 ( .A1(n500), .A2(n538), .ZN(n501) );
  XNOR2_X1 U561 ( .A(n502), .B(n501), .ZN(G1327GAT) );
  NOR2_X1 U562 ( .A1(n569), .A2(n507), .ZN(n504) );
  XNOR2_X1 U563 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n503) );
  XNOR2_X1 U564 ( .A(n504), .B(n503), .ZN(G1328GAT) );
  NOR2_X1 U565 ( .A1(n505), .A2(n507), .ZN(n506) );
  XOR2_X1 U566 ( .A(G36GAT), .B(n506), .Z(G1329GAT) );
  INV_X1 U567 ( .A(n538), .ZN(n508) );
  NOR2_X1 U568 ( .A1(n508), .A2(n507), .ZN(n509) );
  XOR2_X1 U569 ( .A(G50GAT), .B(n509), .Z(G1331GAT) );
  INV_X1 U570 ( .A(n572), .ZN(n510) );
  NAND2_X1 U571 ( .A1(n510), .A2(n554), .ZN(n521) );
  NOR2_X1 U572 ( .A1(n511), .A2(n521), .ZN(n512) );
  XNOR2_X1 U573 ( .A(n512), .B(KEYINPUT108), .ZN(n518) );
  NAND2_X1 U574 ( .A1(n518), .A2(n523), .ZN(n513) );
  XNOR2_X1 U575 ( .A(n513), .B(KEYINPUT42), .ZN(n514) );
  XNOR2_X1 U576 ( .A(G57GAT), .B(n514), .ZN(G1332GAT) );
  XOR2_X1 U577 ( .A(G64GAT), .B(KEYINPUT109), .Z(n516) );
  NAND2_X1 U578 ( .A1(n525), .A2(n518), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n516), .B(n515), .ZN(G1333GAT) );
  NAND2_X1 U580 ( .A1(n518), .A2(n535), .ZN(n517) );
  XNOR2_X1 U581 ( .A(n517), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U582 ( .A(G78GAT), .B(KEYINPUT43), .Z(n520) );
  NAND2_X1 U583 ( .A1(n518), .A2(n538), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  NOR2_X1 U585 ( .A1(n522), .A2(n521), .ZN(n530) );
  NAND2_X1 U586 ( .A1(n530), .A2(n523), .ZN(n524) );
  XNOR2_X1 U587 ( .A(G85GAT), .B(n524), .ZN(G1336GAT) );
  NAND2_X1 U588 ( .A1(n530), .A2(n525), .ZN(n526) );
  XNOR2_X1 U589 ( .A(n526), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n528) );
  NAND2_X1 U591 ( .A1(n530), .A2(n535), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U593 ( .A(G99GAT), .B(n529), .ZN(G1338GAT) );
  NAND2_X1 U594 ( .A1(n538), .A2(n530), .ZN(n531) );
  XNOR2_X1 U595 ( .A(n531), .B(KEYINPUT44), .ZN(n532) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(n532), .ZN(G1339GAT) );
  NOR2_X1 U597 ( .A1(n534), .A2(n533), .ZN(n549) );
  NAND2_X1 U598 ( .A1(n549), .A2(n535), .ZN(n536) );
  XOR2_X1 U599 ( .A(KEYINPUT115), .B(n536), .Z(n537) );
  NOR2_X1 U600 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U601 ( .A(KEYINPUT116), .B(n539), .ZN(n546) );
  NAND2_X1 U602 ( .A1(n546), .A2(n572), .ZN(n540) );
  XNOR2_X1 U603 ( .A(n540), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U604 ( .A(G120GAT), .B(KEYINPUT49), .Z(n542) );
  NAND2_X1 U605 ( .A1(n554), .A2(n546), .ZN(n541) );
  XNOR2_X1 U606 ( .A(n542), .B(n541), .ZN(G1341GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n544) );
  NAND2_X1 U608 ( .A1(n546), .A2(n578), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U610 ( .A(G127GAT), .B(n545), .ZN(G1342GAT) );
  XOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT51), .Z(n548) );
  NAND2_X1 U612 ( .A1(n561), .A2(n546), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(G1343GAT) );
  XOR2_X1 U614 ( .A(G141GAT), .B(KEYINPUT119), .Z(n553) );
  NAND2_X1 U615 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U616 ( .A(KEYINPUT118), .B(n551), .Z(n562) );
  NAND2_X1 U617 ( .A1(n562), .A2(n572), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n553), .B(n552), .ZN(G1344GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n556) );
  NAND2_X1 U620 ( .A1(n554), .A2(n562), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(n557), .ZN(G1345GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n559) );
  NAND2_X1 U624 ( .A1(n562), .A2(n578), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G155GAT), .B(n560), .ZN(G1346GAT) );
  NAND2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U628 ( .A(n563), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U629 ( .A(G169GAT), .B(KEYINPUT123), .Z(n565) );
  NAND2_X1 U630 ( .A1(n566), .A2(n572), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1348GAT) );
  NAND2_X1 U632 ( .A1(n566), .A2(n578), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n574) );
  NAND2_X1 U635 ( .A1(n568), .A2(n569), .ZN(n571) );
  NOR2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n582) );
  NAND2_X1 U637 ( .A1(n582), .A2(n572), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT61), .Z(n577) );
  NAND2_X1 U641 ( .A1(n582), .A2(n388), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  XOR2_X1 U643 ( .A(G211GAT), .B(KEYINPUT127), .Z(n580) );
  NAND2_X1 U644 ( .A1(n582), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1354GAT) );
  NAND2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(n583), .B(KEYINPUT62), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

