//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 0 1 1 1 0 0 0 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n824, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n954, new_n955, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n978, new_n979, new_n980, new_n981, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n990, new_n991, new_n992,
    new_n993, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT99), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G1gat), .ZN(new_n205));
  AOI21_X1  g004(.A(new_n204), .B1(KEYINPUT16), .B2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n202), .B(KEYINPUT99), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(G1gat), .ZN(new_n208));
  OAI21_X1  g007(.A(G8gat), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT16), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n207), .B1(new_n210), .B2(G1gat), .ZN(new_n211));
  INV_X1    g010(.A(G8gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n204), .A2(new_n205), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n209), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G43gat), .B(G50gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT15), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n217), .B(KEYINPUT96), .ZN(new_n218));
  NAND2_X1  g017(.A1(G29gat), .A2(G36gat), .ZN(new_n219));
  XOR2_X1   g018(.A(new_n219), .B(KEYINPUT97), .Z(new_n220));
  NOR2_X1   g019(.A1(new_n216), .A2(KEYINPUT15), .ZN(new_n221));
  INV_X1    g020(.A(G29gat), .ZN(new_n222));
  INV_X1    g021(.A(G36gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(new_n223), .A3(KEYINPUT14), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT14), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(G29gat), .B2(G36gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NOR3_X1   g026(.A1(new_n220), .A2(new_n221), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n218), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(KEYINPUT95), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(new_n219), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n227), .A2(KEYINPUT95), .ZN(new_n232));
  OAI211_X1 g031(.A(KEYINPUT15), .B(new_n216), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n229), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT100), .B1(new_n215), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n214), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n212), .B1(new_n211), .B2(new_n213), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n234), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n234), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT100), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n239), .A2(new_n240), .A3(new_n209), .A4(new_n214), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n235), .A2(new_n238), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(G229gat), .A2(G233gat), .ZN(new_n243));
  XOR2_X1   g042(.A(new_n243), .B(KEYINPUT13), .Z(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  XOR2_X1   g044(.A(KEYINPUT98), .B(KEYINPUT17), .Z(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n234), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n229), .A2(new_n233), .A3(KEYINPUT17), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n238), .B(new_n243), .C1(new_n250), .C2(new_n215), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT18), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n236), .A2(new_n237), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n254), .A2(new_n249), .A3(new_n248), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n255), .A2(KEYINPUT18), .A3(new_n243), .A4(new_n238), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n245), .A2(new_n253), .A3(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G113gat), .B(G141gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(G197gat), .ZN(new_n259));
  XOR2_X1   g058(.A(KEYINPUT11), .B(G169gat), .Z(new_n260));
  XNOR2_X1  g059(.A(new_n259), .B(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n261), .B(KEYINPUT12), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n245), .A2(new_n253), .A3(new_n256), .A4(new_n262), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT21), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT9), .ZN(new_n268));
  INV_X1    g067(.A(G71gat), .ZN(new_n269));
  INV_X1    g068(.A(G78gat), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT101), .ZN(new_n272));
  XOR2_X1   g071(.A(G57gat), .B(G64gat), .Z(new_n273));
  INV_X1    g072(.A(KEYINPUT101), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n274), .B(new_n268), .C1(new_n269), .C2(new_n270), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n272), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G71gat), .B(G78gat), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT102), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n276), .A2(KEYINPUT102), .A3(new_n278), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n272), .A2(new_n273), .A3(new_n277), .A4(new_n275), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n254), .B1(new_n267), .B2(new_n285), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n286), .A2(KEYINPUT104), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(KEYINPUT104), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n289), .B(KEYINPUT103), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n290), .B(G155gat), .ZN(new_n291));
  OR3_X1    g090(.A1(new_n287), .A2(new_n288), .A3(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n291), .B1(new_n287), .B2(new_n288), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n285), .A2(new_n267), .ZN(new_n295));
  NAND2_X1  g094(.A1(G231gat), .A2(G233gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G127gat), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G183gat), .B(G211gat), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n297), .A2(new_n298), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n299), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n301), .B1(new_n299), .B2(new_n302), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n294), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n297), .B(new_n298), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(new_n300), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n308), .A2(new_n303), .A3(new_n292), .A4(new_n293), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(G85gat), .A2(G92gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT105), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT105), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n314), .A2(G85gat), .A3(G92gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n313), .A2(new_n315), .A3(KEYINPUT7), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT7), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n312), .A2(KEYINPUT105), .A3(new_n317), .ZN(new_n318));
  NOR2_X1   g117(.A1(G85gat), .A2(G92gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(G99gat), .A2(G106gat), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n319), .B1(KEYINPUT8), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n316), .A2(new_n318), .A3(new_n321), .ZN(new_n322));
  OR2_X1    g121(.A1(G99gat), .A2(G106gat), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n322), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n320), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n316), .A2(new_n321), .A3(new_n325), .A4(new_n318), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  AND2_X1   g127(.A1(G232gat), .A2(G233gat), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n234), .A2(new_n328), .B1(KEYINPUT41), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n330), .B1(new_n250), .B2(new_n328), .ZN(new_n331));
  XNOR2_X1  g130(.A(G190gat), .B(G218gat), .ZN(new_n332));
  AND2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n331), .A2(new_n332), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT106), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n336), .B1(new_n331), .B2(new_n332), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n329), .A2(KEYINPUT41), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n338), .B(G134gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(G162gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n335), .A2(new_n341), .ZN(new_n342));
  OAI22_X1  g141(.A1(new_n333), .A2(new_n334), .B1(new_n337), .B2(new_n340), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n311), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n285), .A2(new_n327), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n284), .A2(new_n326), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT107), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n347), .B1(new_n348), .B2(new_n324), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n349), .B(new_n283), .C1(new_n348), .C2(new_n324), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(G230gat), .A2(G233gat), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n352), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT10), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n346), .A2(new_n350), .A3(new_n355), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n283), .A2(new_n328), .A3(KEYINPUT10), .A4(new_n284), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n354), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G120gat), .B(G148gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(G176gat), .B(G204gat), .ZN(new_n360));
  XOR2_X1   g159(.A(new_n359), .B(new_n360), .Z(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NOR3_X1   g161(.A1(new_n353), .A2(new_n358), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n362), .B1(new_n353), .B2(new_n358), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n345), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT34), .ZN(new_n368));
  NAND2_X1  g167(.A1(G227gat), .A2(G233gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n369), .B(KEYINPUT64), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n368), .B1(new_n371), .B2(KEYINPUT75), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(G134gat), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n374), .A2(KEYINPUT71), .A3(G127gat), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT71), .ZN(new_n377));
  XNOR2_X1  g176(.A(G127gat), .B(G134gat), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(G120gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(G113gat), .ZN(new_n381));
  INV_X1    g180(.A(G113gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(G120gat), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT1), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n374), .A2(G127gat), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT72), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT1), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n298), .A2(G134gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(KEYINPUT72), .A2(KEYINPUT1), .ZN(new_n391));
  AND4_X1   g190(.A1(new_n386), .A2(new_n389), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n381), .A2(new_n383), .ZN(new_n393));
  AOI22_X1  g192(.A1(new_n379), .A2(new_n385), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G183gat), .A2(G190gat), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT24), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n398));
  INV_X1    g197(.A(G183gat), .ZN(new_n399));
  INV_X1    g198(.A(G190gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n397), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT23), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n403), .A2(G176gat), .ZN(new_n404));
  INV_X1    g203(.A(G169gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT65), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT65), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(G169gat), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n404), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(G169gat), .A2(G176gat), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT66), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n403), .B1(G169gat), .B2(G176gat), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n402), .A2(new_n409), .A3(new_n414), .A4(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT25), .ZN(new_n417));
  AND3_X1   g216(.A1(new_n416), .A2(KEYINPUT67), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT67), .B1(new_n416), .B2(new_n417), .ZN(new_n419));
  AND3_X1   g218(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n415), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(G176gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT23), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT25), .B1(new_n424), .B2(G169gat), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT68), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n395), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(KEYINPUT68), .A2(G183gat), .A3(G190gat), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n428), .A2(new_n396), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n399), .A2(KEYINPUT69), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT69), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(G183gat), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n431), .A2(new_n433), .A3(new_n400), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n430), .A2(new_n434), .A3(new_n398), .ZN(new_n435));
  AND2_X1   g234(.A1(new_n426), .A2(new_n435), .ZN(new_n436));
  NOR3_X1   g235(.A1(new_n418), .A2(new_n419), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n405), .A2(new_n423), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(KEYINPUT26), .ZN(new_n439));
  INV_X1    g238(.A(new_n414), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n395), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(KEYINPUT27), .B(G183gat), .ZN(new_n442));
  AND2_X1   g241(.A1(new_n400), .A2(KEYINPUT28), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(KEYINPUT70), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT70), .B1(new_n442), .B2(new_n443), .ZN(new_n446));
  OR2_X1    g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT27), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n399), .ZN(new_n449));
  XNOR2_X1  g248(.A(KEYINPUT69), .B(G183gat), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n449), .B1(new_n450), .B2(new_n448), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT28), .B1(new_n451), .B2(new_n400), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n441), .B1(new_n447), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n394), .B1(new_n437), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n416), .A2(new_n417), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT67), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n416), .A2(KEYINPUT67), .A3(new_n417), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n426), .A2(new_n435), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  OR2_X1    g260(.A1(new_n439), .A2(new_n440), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n445), .A2(new_n446), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n462), .B(new_n395), .C1(new_n463), .C2(new_n452), .ZN(new_n464));
  AND2_X1   g263(.A1(KEYINPUT72), .A2(KEYINPUT1), .ZN(new_n465));
  NOR2_X1   g264(.A1(KEYINPUT72), .A2(KEYINPUT1), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n393), .A2(new_n467), .A3(new_n378), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n386), .A2(new_n390), .A3(new_n377), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n375), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n468), .B1(new_n470), .B2(new_n384), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n461), .A2(new_n464), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n455), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n373), .B1(new_n473), .B2(new_n371), .ZN(new_n474));
  AOI211_X1 g273(.A(new_n370), .B(new_n372), .C1(new_n455), .C2(new_n472), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n455), .A2(new_n370), .A3(new_n472), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT32), .ZN(new_n478));
  XOR2_X1   g277(.A(KEYINPUT73), .B(KEYINPUT33), .Z(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  XOR2_X1   g279(.A(G15gat), .B(G43gat), .Z(new_n481));
  XNOR2_X1  g280(.A(G71gat), .B(G99gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n481), .B(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n478), .A2(new_n480), .A3(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n483), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n477), .B(KEYINPUT32), .C1(new_n479), .C2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n476), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n476), .B1(new_n484), .B2(new_n486), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT93), .ZN(new_n490));
  OR3_X1    g289(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n490), .B1(new_n488), .B2(new_n489), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(G228gat), .A2(G233gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n494), .B(KEYINPUT88), .ZN(new_n495));
  AND2_X1   g294(.A1(G155gat), .A2(G162gat), .ZN(new_n496));
  NOR2_X1   g295(.A1(G155gat), .A2(G162gat), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(G141gat), .B(G148gat), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT2), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n500), .B1(G155gat), .B2(G162gat), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n498), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(G141gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(G148gat), .ZN(new_n504));
  INV_X1    g303(.A(G148gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(G141gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G155gat), .B(G162gat), .ZN(new_n508));
  INV_X1    g307(.A(G155gat), .ZN(new_n509));
  INV_X1    g308(.A(G162gat), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT2), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n507), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n502), .A2(new_n512), .ZN(new_n513));
  XOR2_X1   g312(.A(G197gat), .B(G204gat), .Z(new_n514));
  INV_X1    g313(.A(KEYINPUT77), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n515), .A2(G211gat), .ZN(new_n516));
  INV_X1    g315(.A(G211gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n517), .A2(KEYINPUT77), .ZN(new_n518));
  OAI21_X1  g317(.A(G218gat), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT76), .B(KEYINPUT22), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n514), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(G211gat), .B(G218gat), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT90), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(KEYINPUT77), .B(G211gat), .ZN(new_n524));
  INV_X1    g323(.A(G218gat), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n520), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(G197gat), .B(G204gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT90), .ZN(new_n529));
  INV_X1    g328(.A(new_n522), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n517), .A2(KEYINPUT77), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n515), .A2(G211gat), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n525), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  XOR2_X1   g333(.A(KEYINPUT76), .B(KEYINPUT22), .Z(new_n535));
  OAI211_X1 g334(.A(new_n522), .B(new_n527), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT89), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT89), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n526), .A2(new_n538), .A3(new_n522), .A4(new_n527), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n523), .A2(new_n531), .A3(new_n537), .A4(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT29), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT3), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n513), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT79), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT78), .B1(new_n522), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n528), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT78), .ZN(new_n549));
  AOI21_X1  g348(.A(KEYINPUT79), .B1(new_n521), .B2(new_n549), .ZN(new_n550));
  OAI211_X1 g349(.A(KEYINPUT80), .B(new_n548), .C1(new_n550), .C2(new_n522), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT80), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n549), .B(new_n527), .C1(new_n534), .C2(new_n535), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n522), .B1(new_n553), .B2(new_n545), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n521), .A2(new_n546), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n552), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n502), .A2(new_n512), .A3(new_n543), .ZN(new_n557));
  AOI22_X1  g356(.A1(new_n551), .A2(new_n556), .B1(new_n541), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n495), .B1(new_n544), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n551), .A2(new_n556), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n557), .A2(new_n541), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT84), .ZN(new_n563));
  AND3_X1   g362(.A1(new_n507), .A2(new_n508), .A3(new_n511), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n508), .B1(new_n511), .B2(new_n507), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n502), .A2(new_n512), .A3(KEYINPUT84), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NOR3_X1   g367(.A1(new_n554), .A2(new_n555), .A3(KEYINPUT29), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n568), .B1(new_n569), .B2(KEYINPUT3), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n562), .A2(G228gat), .A3(G233gat), .A4(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G78gat), .B(G106gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(KEYINPUT31), .B(G50gat), .ZN(new_n573));
  XOR2_X1   g372(.A(new_n572), .B(new_n573), .Z(new_n574));
  NOR2_X1   g373(.A1(new_n574), .A2(KEYINPUT91), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n559), .A2(new_n571), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(G22gat), .ZN(new_n578));
  INV_X1    g377(.A(new_n574), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT91), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(G22gat), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n559), .A2(new_n571), .A3(new_n582), .A4(new_n576), .ZN(new_n583));
  AND3_X1   g382(.A1(new_n578), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n581), .B1(new_n578), .B2(new_n583), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT81), .ZN(new_n587));
  NAND2_X1  g386(.A1(G226gat), .A2(G233gat), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n588), .B1(new_n461), .B2(new_n464), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n541), .B1(new_n437), .B2(new_n454), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n589), .B1(new_n590), .B2(new_n588), .ZN(new_n591));
  INV_X1    g390(.A(new_n560), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n587), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n590), .A2(new_n588), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT82), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n589), .A2(new_n595), .ZN(new_n596));
  AOI211_X1 g395(.A(KEYINPUT82), .B(new_n588), .C1(new_n461), .C2(new_n464), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n594), .B(new_n592), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(KEYINPUT29), .B1(new_n461), .B2(new_n464), .ZN(new_n599));
  INV_X1    g398(.A(new_n588), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI211_X1 g400(.A(KEYINPUT81), .B(new_n560), .C1(new_n601), .C2(new_n589), .ZN(new_n602));
  XNOR2_X1  g401(.A(G8gat), .B(G36gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(G64gat), .B(G92gat), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n603), .B(new_n604), .Z(new_n605));
  NAND4_X1  g404(.A1(new_n593), .A2(new_n598), .A3(new_n602), .A4(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(KEYINPUT83), .B(KEYINPUT30), .Z(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AND2_X1   g407(.A1(new_n605), .A2(KEYINPUT30), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n593), .A2(new_n598), .A3(new_n602), .A4(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n593), .A2(new_n598), .A3(new_n602), .ZN(new_n611));
  INV_X1    g410(.A(new_n605), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n608), .A2(new_n610), .A3(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n394), .A2(KEYINPUT4), .A3(new_n513), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT4), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n502), .A2(new_n512), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n616), .B1(new_n471), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  AND3_X1   g419(.A1(new_n502), .A2(new_n512), .A3(KEYINPUT84), .ZN(new_n621));
  AOI21_X1  g420(.A(KEYINPUT84), .B1(new_n502), .B2(new_n512), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n471), .B(new_n557), .C1(new_n623), .C2(new_n543), .ZN(new_n624));
  NAND2_X1  g423(.A1(G225gat), .A2(G233gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT85), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n620), .A2(new_n624), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n394), .B1(new_n566), .B2(new_n567), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n471), .A2(new_n617), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n626), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(KEYINPUT86), .B1(new_n631), .B2(KEYINPUT5), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n471), .B1(new_n621), .B2(new_n622), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n394), .A2(new_n513), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n627), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT86), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT5), .ZN(new_n637));
  NOR3_X1   g436(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n628), .B1(new_n632), .B2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(G1gat), .B(G29gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT0), .ZN(new_n641));
  XNOR2_X1  g440(.A(G57gat), .B(G85gat), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n641), .B(new_n642), .Z(new_n643));
  NAND2_X1  g442(.A1(new_n471), .A2(new_n557), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n644), .B1(new_n568), .B2(KEYINPUT3), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n645), .A2(new_n619), .A3(new_n626), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(new_n637), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n639), .A2(new_n643), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n643), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n636), .B1(new_n635), .B2(new_n637), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n630), .B1(new_n568), .B2(new_n471), .ZN(new_n651));
  OAI211_X1 g450(.A(KEYINPUT86), .B(KEYINPUT5), .C1(new_n651), .C2(new_n627), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n646), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n628), .A2(KEYINPUT5), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n649), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT6), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n648), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  OAI211_X1 g456(.A(KEYINPUT6), .B(new_n649), .C1(new_n653), .C2(new_n654), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT35), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n586), .A2(new_n614), .A3(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n493), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT74), .ZN(new_n662));
  AND3_X1   g461(.A1(new_n484), .A2(new_n662), .A3(new_n486), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n662), .B1(new_n484), .B2(new_n486), .ZN(new_n664));
  OAI22_X1  g463(.A1(new_n663), .A2(new_n664), .B1(new_n475), .B2(new_n474), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n578), .A2(new_n581), .A3(new_n583), .ZN(new_n666));
  INV_X1    g465(.A(new_n581), .ZN(new_n667));
  AOI21_X1  g466(.A(KEYINPUT3), .B1(new_n540), .B2(new_n541), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n562), .B1(new_n513), .B2(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n575), .B1(new_n669), .B2(new_n495), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n582), .B1(new_n670), .B2(new_n571), .ZN(new_n671));
  INV_X1    g470(.A(new_n583), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n667), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n665), .A2(new_n666), .A3(new_n673), .A4(new_n487), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n657), .A2(KEYINPUT87), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT87), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n648), .A2(new_n655), .A3(new_n676), .A4(new_n656), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n675), .A2(new_n677), .A3(new_n658), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n614), .ZN(new_n679));
  OAI21_X1  g478(.A(KEYINPUT35), .B1(new_n674), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(KEYINPUT94), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n584), .A2(new_n585), .A3(new_n488), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n682), .A2(new_n678), .A3(new_n614), .A4(new_n665), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT94), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n683), .A2(new_n684), .A3(KEYINPUT35), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n661), .B1(new_n681), .B2(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n627), .B1(new_n620), .B2(new_n624), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT39), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n649), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n651), .A2(new_n627), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(KEYINPUT39), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n689), .B1(new_n687), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT40), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n655), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n692), .ZN(new_n695));
  OAI21_X1  g494(.A(KEYINPUT92), .B1(new_n695), .B2(KEYINPUT40), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT92), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n692), .A2(new_n697), .A3(new_n693), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n694), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n608), .A2(new_n610), .A3(new_n613), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT37), .ZN(new_n702));
  INV_X1    g501(.A(new_n589), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n594), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n702), .B1(new_n704), .B2(new_n592), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n594), .B(new_n560), .C1(new_n596), .C2(new_n597), .ZN(new_n706));
  AOI21_X1  g505(.A(KEYINPUT38), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  OAI211_X1 g506(.A(new_n707), .B(new_n612), .C1(new_n611), .C2(KEYINPUT37), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n708), .A2(new_n657), .A3(new_n658), .A4(new_n606), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT38), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n613), .B1(new_n702), .B2(new_n605), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n611), .A2(KEYINPUT37), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n586), .B(new_n701), .C1(new_n709), .C2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n586), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n679), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT36), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n717), .B1(new_n488), .B2(new_n489), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n484), .A2(new_n486), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(KEYINPUT74), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n484), .A2(new_n662), .A3(new_n486), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n476), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n487), .A2(KEYINPUT36), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n718), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n714), .A2(new_n716), .A3(new_n724), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n266), .B(new_n367), .C1(new_n686), .C2(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n726), .A2(new_n678), .ZN(new_n727));
  XNOR2_X1  g526(.A(KEYINPUT108), .B(G1gat), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1324gat));
  INV_X1    g528(.A(new_n726), .ZN(new_n730));
  XOR2_X1   g529(.A(KEYINPUT16), .B(G8gat), .Z(new_n731));
  NAND4_X1  g530(.A1(new_n730), .A2(KEYINPUT42), .A3(new_n700), .A4(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n730), .A2(KEYINPUT109), .A3(new_n700), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT109), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n734), .B1(new_n726), .B2(new_n614), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n733), .A2(G8gat), .A3(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n731), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n737), .B1(new_n733), .B2(new_n735), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n732), .B(new_n736), .C1(new_n738), .C2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g538(.A(KEYINPUT110), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n740), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n718), .B(KEYINPUT110), .C1(new_n722), .C2(new_n723), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(G15gat), .B1(new_n726), .B2(new_n743), .ZN(new_n744));
  OR2_X1    g543(.A1(new_n493), .A2(G15gat), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n726), .B2(new_n745), .ZN(G1326gat));
  NAND3_X1  g545(.A1(new_n730), .A2(KEYINPUT111), .A3(new_n715), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT111), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(new_n726), .B2(new_n586), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(KEYINPUT43), .B(G22gat), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1327gat));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n344), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n686), .B2(new_n725), .ZN(new_n755));
  INV_X1    g554(.A(new_n366), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n310), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n266), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n661), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT35), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n673), .A2(new_n666), .A3(new_n487), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n762), .A2(new_n722), .ZN(new_n763));
  INV_X1    g562(.A(new_n658), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n764), .B1(new_n657), .B2(KEYINPUT87), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n700), .B1(new_n677), .B2(new_n765), .ZN(new_n766));
  AOI211_X1 g565(.A(KEYINPUT94), .B(new_n761), .C1(new_n763), .C2(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n684), .B1(new_n683), .B2(KEYINPUT35), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n760), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n743), .A2(new_n716), .A3(new_n714), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n344), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n755), .B(new_n759), .C1(new_n771), .C2(KEYINPUT44), .ZN(new_n772));
  OAI21_X1  g571(.A(G29gat), .B1(new_n772), .B2(new_n678), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT45), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n757), .A2(new_n344), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n266), .B(new_n775), .C1(new_n686), .C2(new_n725), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n678), .A2(G29gat), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n774), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  OR3_X1    g578(.A1(new_n776), .A2(new_n774), .A3(new_n778), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n773), .A2(new_n779), .A3(new_n780), .ZN(G1328gat));
  INV_X1    g580(.A(KEYINPUT112), .ZN(new_n782));
  AOI211_X1 g581(.A(G36gat), .B(new_n614), .C1(new_n782), .C2(KEYINPUT46), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n776), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n782), .A2(KEYINPUT46), .ZN(new_n786));
  XOR2_X1   g585(.A(new_n785), .B(new_n786), .Z(new_n787));
  OAI21_X1  g586(.A(KEYINPUT113), .B1(new_n772), .B2(new_n614), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(G36gat), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n772), .A2(KEYINPUT113), .A3(new_n614), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n787), .B1(new_n789), .B2(new_n790), .ZN(G1329gat));
  OAI21_X1  g590(.A(G43gat), .B1(new_n772), .B2(new_n743), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT47), .ZN(new_n793));
  OR3_X1    g592(.A1(new_n776), .A2(G43gat), .A3(new_n493), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n793), .B1(new_n792), .B2(new_n794), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n795), .A2(new_n796), .ZN(G1330gat));
  NAND2_X1  g596(.A1(new_n715), .A2(G50gat), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n776), .A2(new_n586), .ZN(new_n799));
  OAI22_X1  g598(.A1(new_n772), .A2(new_n798), .B1(new_n799), .B2(G50gat), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(KEYINPUT48), .ZN(G1331gat));
  NOR3_X1   g600(.A1(new_n345), .A2(new_n266), .A3(new_n756), .ZN(new_n802));
  AND4_X1   g601(.A1(new_n716), .A2(new_n714), .A3(new_n741), .A4(new_n742), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n802), .B1(new_n686), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n804), .A2(new_n678), .ZN(new_n805));
  XOR2_X1   g604(.A(new_n805), .B(G57gat), .Z(G1332gat));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  OAI211_X1 g607(.A(KEYINPUT114), .B(new_n802), .C1(new_n686), .C2(new_n803), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT49), .ZN(new_n810));
  INV_X1    g609(.A(G64gat), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n700), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  XOR2_X1   g611(.A(new_n812), .B(KEYINPUT115), .Z(new_n813));
  NAND3_X1  g612(.A1(new_n808), .A2(new_n809), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n810), .A2(new_n811), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n814), .B(new_n815), .ZN(G1333gat));
  NOR3_X1   g615(.A1(new_n804), .A2(G71gat), .A3(new_n493), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n741), .A2(new_n742), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n808), .A2(new_n809), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n817), .B1(new_n819), .B2(G71gat), .ZN(new_n820));
  XNOR2_X1  g619(.A(KEYINPUT116), .B(KEYINPUT50), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n820), .B(new_n822), .ZN(G1334gat));
  NAND3_X1  g622(.A1(new_n808), .A2(new_n809), .A3(new_n715), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n824), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g624(.A1(new_n311), .A2(new_n266), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT51), .B1(new_n771), .B2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n344), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n828), .B(new_n826), .C1(new_n686), .C2(new_n803), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT51), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OR2_X1    g630(.A1(new_n827), .A2(new_n831), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n678), .A2(new_n756), .A3(G85gat), .ZN(new_n833));
  XOR2_X1   g632(.A(new_n833), .B(KEYINPUT117), .Z(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n311), .A2(new_n266), .A3(new_n756), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n755), .B(new_n836), .C1(new_n771), .C2(KEYINPUT44), .ZN(new_n837));
  OAI21_X1  g636(.A(G85gat), .B1(new_n837), .B2(new_n678), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n835), .A2(new_n838), .ZN(G1336gat));
  OAI21_X1  g638(.A(G92gat), .B1(new_n837), .B2(new_n614), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n614), .A2(new_n756), .A3(G92gat), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n841), .B1(new_n827), .B2(new_n831), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT52), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT52), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n840), .A2(new_n842), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n844), .A2(new_n846), .ZN(G1337gat));
  NOR3_X1   g646(.A1(new_n493), .A2(G99gat), .A3(new_n756), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(G99gat), .B1(new_n837), .B2(new_n743), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(G1338gat));
  NOR3_X1   g650(.A1(new_n586), .A2(new_n756), .A3(G106gat), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n852), .B1(new_n827), .B2(new_n831), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT118), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n828), .B1(new_n686), .B2(new_n803), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n753), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n857), .A2(new_n715), .A3(new_n755), .A4(new_n836), .ZN(new_n858));
  AOI21_X1  g657(.A(KEYINPUT53), .B1(new_n858), .B2(G106gat), .ZN(new_n859));
  OAI211_X1 g658(.A(KEYINPUT118), .B(new_n852), .C1(new_n827), .C2(new_n831), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n855), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(G106gat), .B1(new_n837), .B2(new_n586), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n853), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(KEYINPUT53), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n861), .A2(new_n864), .ZN(G1339gat));
  NAND3_X1  g664(.A1(new_n356), .A2(new_n357), .A3(new_n354), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT119), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n356), .A2(new_n357), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n352), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n356), .A2(new_n357), .A3(KEYINPUT119), .A4(new_n354), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n868), .A2(new_n870), .A3(KEYINPUT54), .A4(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT54), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n361), .B1(new_n358), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT55), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI211_X1 g676(.A(new_n876), .B(new_n361), .C1(new_n358), .C2(new_n873), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n363), .B1(new_n878), .B2(new_n872), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n877), .A2(new_n266), .A3(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n242), .A2(new_n244), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n243), .B1(new_n255), .B2(new_n238), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n261), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n366), .A2(new_n265), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n828), .B1(new_n880), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n877), .A2(new_n879), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n342), .A2(new_n883), .A3(new_n343), .A4(new_n265), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n310), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n311), .A2(new_n758), .A3(new_n344), .A4(new_n756), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n715), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n678), .A2(new_n700), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n891), .A2(new_n491), .A3(new_n492), .A4(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(G113gat), .B1(new_n893), .B2(new_n758), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n678), .B1(new_n889), .B2(new_n890), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n895), .A2(new_n763), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n614), .ZN(new_n897));
  XOR2_X1   g696(.A(new_n897), .B(KEYINPUT120), .Z(new_n898));
  NAND2_X1  g697(.A1(new_n266), .A2(new_n382), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n894), .B1(new_n898), .B2(new_n899), .ZN(G1340gat));
  OAI21_X1  g699(.A(G120gat), .B1(new_n893), .B2(new_n756), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n366), .A2(new_n380), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n901), .B1(new_n898), .B2(new_n902), .ZN(G1341gat));
  OAI21_X1  g702(.A(G127gat), .B1(new_n893), .B2(new_n310), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n311), .A2(new_n298), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n897), .B2(new_n905), .ZN(G1342gat));
  NAND2_X1  g705(.A1(new_n828), .A2(new_n614), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT121), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n896), .A2(new_n374), .A3(new_n909), .ZN(new_n910));
  OR2_X1    g709(.A1(new_n910), .A2(KEYINPUT56), .ZN(new_n911));
  OAI21_X1  g710(.A(G134gat), .B1(new_n893), .B2(new_n344), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(KEYINPUT56), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(G1343gat));
  NOR2_X1   g713(.A1(new_n818), .A2(new_n586), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n895), .A2(new_n915), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n916), .A2(new_n614), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n266), .A2(new_n503), .ZN(new_n918));
  XOR2_X1   g717(.A(new_n918), .B(KEYINPUT124), .Z(new_n919));
  AOI21_X1  g718(.A(KEYINPUT58), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n889), .A2(new_n890), .ZN(new_n921));
  AOI21_X1  g720(.A(KEYINPUT57), .B1(new_n921), .B2(new_n715), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT57), .ZN(new_n923));
  AOI211_X1 g722(.A(new_n923), .B(new_n586), .C1(new_n889), .C2(new_n890), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(new_n892), .ZN(new_n926));
  OR3_X1    g725(.A1(new_n818), .A2(KEYINPUT122), .A3(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(KEYINPUT122), .B1(new_n818), .B2(new_n926), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n925), .A2(new_n758), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n920), .B1(new_n503), .B2(new_n930), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n917), .A2(new_n919), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT123), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n933), .B1(new_n925), .B2(new_n929), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n927), .A2(new_n928), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n935), .B(KEYINPUT123), .C1(new_n922), .C2(new_n924), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n934), .A2(new_n266), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n932), .B1(new_n937), .B2(G141gat), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT58), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n931), .B1(new_n938), .B2(new_n939), .ZN(G1344gat));
  NAND3_X1  g739(.A1(new_n934), .A2(new_n366), .A3(new_n936), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(G148gat), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT59), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(new_n925), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n945), .A2(new_n366), .A3(new_n935), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n943), .A2(new_n505), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n756), .A2(G148gat), .ZN(new_n948));
  AOI22_X1  g747(.A1(new_n946), .A2(new_n947), .B1(new_n917), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n944), .A2(new_n949), .ZN(G1345gat));
  NAND3_X1  g749(.A1(new_n917), .A2(new_n509), .A3(new_n311), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n934), .A2(new_n311), .A3(new_n936), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n952), .B2(new_n509), .ZN(G1346gat));
  NAND3_X1  g752(.A1(new_n916), .A2(new_n510), .A3(new_n909), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n934), .A2(new_n828), .A3(new_n936), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n954), .B1(new_n955), .B2(new_n510), .ZN(G1347gat));
  INV_X1    g755(.A(new_n678), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n957), .B1(new_n889), .B2(new_n890), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n674), .A2(new_n614), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(KEYINPUT125), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT125), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n958), .A2(new_n962), .A3(new_n959), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n964), .A2(new_n406), .A3(new_n408), .A4(new_n266), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n678), .A2(new_n700), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n493), .A2(new_n966), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n891), .A2(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(new_n968), .ZN(new_n969));
  OAI21_X1  g768(.A(G169gat), .B1(new_n969), .B2(new_n758), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n970), .A2(new_n971), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n965), .B1(new_n972), .B2(new_n973), .ZN(G1348gat));
  NAND3_X1  g773(.A1(new_n964), .A2(new_n423), .A3(new_n366), .ZN(new_n975));
  OAI21_X1  g774(.A(G176gat), .B1(new_n969), .B2(new_n756), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(G1349gat));
  AOI21_X1  g776(.A(new_n450), .B1(new_n968), .B2(new_n311), .ZN(new_n978));
  INV_X1    g777(.A(new_n442), .ZN(new_n979));
  NOR3_X1   g778(.A1(new_n960), .A2(new_n979), .A3(new_n310), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  XOR2_X1   g780(.A(new_n981), .B(KEYINPUT60), .Z(G1350gat));
  NAND4_X1  g781(.A1(new_n961), .A2(new_n400), .A3(new_n828), .A4(new_n963), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT61), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n891), .A2(new_n828), .A3(new_n967), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n984), .B1(new_n985), .B2(G190gat), .ZN(new_n986));
  AND3_X1   g785(.A1(new_n985), .A2(new_n984), .A3(G190gat), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n983), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  XOR2_X1   g787(.A(new_n988), .B(KEYINPUT127), .Z(G1351gat));
  AND3_X1   g788(.A1(new_n958), .A2(new_n700), .A3(new_n915), .ZN(new_n990));
  AOI21_X1  g789(.A(G197gat), .B1(new_n990), .B2(new_n266), .ZN(new_n991));
  NOR3_X1   g790(.A1(new_n925), .A2(new_n818), .A3(new_n966), .ZN(new_n992));
  AND2_X1   g791(.A1(new_n266), .A2(G197gat), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n991), .B1(new_n992), .B2(new_n993), .ZN(G1352gat));
  INV_X1    g793(.A(G204gat), .ZN(new_n995));
  AOI21_X1  g794(.A(new_n995), .B1(new_n992), .B2(new_n366), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n990), .A2(new_n995), .A3(new_n366), .ZN(new_n997));
  AND2_X1   g796(.A1(new_n997), .A2(KEYINPUT62), .ZN(new_n998));
  NOR2_X1   g797(.A1(new_n997), .A2(KEYINPUT62), .ZN(new_n999));
  OR3_X1    g798(.A1(new_n996), .A2(new_n998), .A3(new_n999), .ZN(G1353gat));
  NAND3_X1  g799(.A1(new_n990), .A2(new_n524), .A3(new_n311), .ZN(new_n1001));
  NOR2_X1   g800(.A1(new_n818), .A2(new_n966), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n945), .A2(new_n311), .A3(new_n1002), .ZN(new_n1003));
  AND3_X1   g802(.A1(new_n1003), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1004));
  AOI21_X1  g803(.A(KEYINPUT63), .B1(new_n1003), .B2(G211gat), .ZN(new_n1005));
  OAI21_X1  g804(.A(new_n1001), .B1(new_n1004), .B2(new_n1005), .ZN(G1354gat));
  NAND3_X1  g805(.A1(new_n990), .A2(new_n525), .A3(new_n828), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n828), .ZN(new_n1008));
  INV_X1    g807(.A(new_n1008), .ZN(new_n1009));
  OAI21_X1  g808(.A(new_n1007), .B1(new_n1009), .B2(new_n525), .ZN(G1355gat));
endmodule


