

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X1 U555 ( .A(n721), .Z(n764) );
  NOR2_X1 U556 ( .A1(G651), .A2(G543), .ZN(n647) );
  XNOR2_X1 U557 ( .A(KEYINPUT26), .B(KEYINPUT64), .ZN(n722) );
  XNOR2_X1 U558 ( .A(n723), .B(n722), .ZN(n726) );
  NOR2_X1 U559 ( .A1(n727), .A2(n977), .ZN(n730) );
  NAND2_X1 U560 ( .A1(G160), .A2(G40), .ZN(n716) );
  NOR2_X2 U561 ( .A1(G651), .A2(n633), .ZN(n650) );
  AND2_X2 U562 ( .A1(n520), .A2(G2104), .ZN(n886) );
  XNOR2_X1 U563 ( .A(n524), .B(n523), .ZN(n889) );
  NOR2_X1 U564 ( .A1(n548), .A2(n547), .ZN(G160) );
  INV_X1 U565 ( .A(G2105), .ZN(n520) );
  NAND2_X1 U566 ( .A1(n886), .A2(G102), .ZN(n519) );
  XNOR2_X1 U567 ( .A(n519), .B(KEYINPUT92), .ZN(n522) );
  NOR2_X1 U568 ( .A1(G2104), .A2(n520), .ZN(n882) );
  NAND2_X1 U569 ( .A1(G126), .A2(n882), .ZN(n521) );
  NAND2_X1 U570 ( .A1(n522), .A2(n521), .ZN(n528) );
  XNOR2_X1 U571 ( .A(KEYINPUT17), .B(KEYINPUT65), .ZN(n524) );
  NOR2_X1 U572 ( .A1(G2105), .A2(G2104), .ZN(n523) );
  NAND2_X1 U573 ( .A1(n889), .A2(G138), .ZN(n526) );
  AND2_X1 U574 ( .A1(G2105), .A2(G2104), .ZN(n881) );
  NAND2_X1 U575 ( .A1(G114), .A2(n881), .ZN(n525) );
  NAND2_X1 U576 ( .A1(n526), .A2(n525), .ZN(n527) );
  NOR2_X1 U577 ( .A1(n528), .A2(n527), .ZN(G164) );
  NAND2_X1 U578 ( .A1(n647), .A2(G89), .ZN(n529) );
  XNOR2_X1 U579 ( .A(n529), .B(KEYINPUT4), .ZN(n531) );
  XOR2_X1 U580 ( .A(KEYINPUT0), .B(G543), .Z(n633) );
  INV_X1 U581 ( .A(G651), .ZN(n534) );
  NOR2_X1 U582 ( .A1(n633), .A2(n534), .ZN(n653) );
  NAND2_X1 U583 ( .A1(G76), .A2(n653), .ZN(n530) );
  NAND2_X1 U584 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U585 ( .A(n532), .B(KEYINPUT5), .ZN(n540) );
  NAND2_X1 U586 ( .A1(n650), .A2(G51), .ZN(n533) );
  XNOR2_X1 U587 ( .A(n533), .B(KEYINPUT76), .ZN(n537) );
  NOR2_X1 U588 ( .A1(G543), .A2(n534), .ZN(n535) );
  XOR2_X1 U589 ( .A(KEYINPUT1), .B(n535), .Z(n649) );
  NAND2_X1 U590 ( .A1(G63), .A2(n649), .ZN(n536) );
  NAND2_X1 U591 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U592 ( .A(KEYINPUT6), .B(n538), .Z(n539) );
  NAND2_X1 U593 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U594 ( .A(n541), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U595 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U596 ( .A1(n889), .A2(G137), .ZN(n544) );
  NAND2_X1 U597 ( .A1(G101), .A2(n886), .ZN(n542) );
  XOR2_X1 U598 ( .A(KEYINPUT23), .B(n542), .Z(n543) );
  NAND2_X1 U599 ( .A1(n544), .A2(n543), .ZN(n548) );
  NAND2_X1 U600 ( .A1(G113), .A2(n881), .ZN(n546) );
  NAND2_X1 U601 ( .A1(G125), .A2(n882), .ZN(n545) );
  NAND2_X1 U602 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U603 ( .A(G2435), .B(G2454), .Z(n550) );
  XNOR2_X1 U604 ( .A(G2430), .B(G2438), .ZN(n549) );
  XNOR2_X1 U605 ( .A(n550), .B(n549), .ZN(n557) );
  XOR2_X1 U606 ( .A(G2446), .B(KEYINPUT107), .Z(n552) );
  XNOR2_X1 U607 ( .A(G2451), .B(G2443), .ZN(n551) );
  XNOR2_X1 U608 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U609 ( .A(n553), .B(G2427), .Z(n555) );
  XNOR2_X1 U610 ( .A(G1348), .B(G1341), .ZN(n554) );
  XNOR2_X1 U611 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U612 ( .A(n557), .B(n556), .ZN(n558) );
  AND2_X1 U613 ( .A1(n558), .A2(G14), .ZN(G401) );
  NAND2_X1 U614 ( .A1(n649), .A2(G64), .ZN(n559) );
  XNOR2_X1 U615 ( .A(n559), .B(KEYINPUT68), .ZN(n561) );
  NAND2_X1 U616 ( .A1(G52), .A2(n650), .ZN(n560) );
  NAND2_X1 U617 ( .A1(n561), .A2(n560), .ZN(n567) );
  NAND2_X1 U618 ( .A1(n653), .A2(G77), .ZN(n562) );
  XOR2_X1 U619 ( .A(KEYINPUT69), .B(n562), .Z(n564) );
  NAND2_X1 U620 ( .A1(n647), .A2(G90), .ZN(n563) );
  NAND2_X1 U621 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U622 ( .A(KEYINPUT9), .B(n565), .Z(n566) );
  NOR2_X1 U623 ( .A1(n567), .A2(n566), .ZN(G171) );
  AND2_X1 U624 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U625 ( .A1(G99), .A2(n886), .ZN(n569) );
  NAND2_X1 U626 ( .A1(G111), .A2(n881), .ZN(n568) );
  NAND2_X1 U627 ( .A1(n569), .A2(n568), .ZN(n572) );
  NAND2_X1 U628 ( .A1(n882), .A2(G123), .ZN(n570) );
  XOR2_X1 U629 ( .A(KEYINPUT18), .B(n570), .Z(n571) );
  NOR2_X1 U630 ( .A1(n572), .A2(n571), .ZN(n574) );
  NAND2_X1 U631 ( .A1(n889), .A2(G135), .ZN(n573) );
  NAND2_X1 U632 ( .A1(n574), .A2(n573), .ZN(n930) );
  XNOR2_X1 U633 ( .A(G2096), .B(n930), .ZN(n575) );
  OR2_X1 U634 ( .A1(G2100), .A2(n575), .ZN(G156) );
  INV_X1 U635 ( .A(G132), .ZN(G219) );
  INV_X1 U636 ( .A(G57), .ZN(G237) );
  INV_X1 U637 ( .A(G69), .ZN(G235) );
  INV_X1 U638 ( .A(G108), .ZN(G238) );
  INV_X1 U639 ( .A(G120), .ZN(G236) );
  NAND2_X1 U640 ( .A1(G75), .A2(n653), .ZN(n577) );
  NAND2_X1 U641 ( .A1(G88), .A2(n647), .ZN(n576) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n581) );
  NAND2_X1 U643 ( .A1(G62), .A2(n649), .ZN(n579) );
  NAND2_X1 U644 ( .A1(G50), .A2(n650), .ZN(n578) );
  NAND2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U646 ( .A1(n581), .A2(n580), .ZN(G166) );
  NAND2_X1 U647 ( .A1(G7), .A2(G661), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n582), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U649 ( .A(G223), .ZN(n831) );
  NAND2_X1 U650 ( .A1(n831), .A2(G567), .ZN(n583) );
  XOR2_X1 U651 ( .A(KEYINPUT11), .B(n583), .Z(G234) );
  NAND2_X1 U652 ( .A1(n647), .A2(G81), .ZN(n584) );
  XNOR2_X1 U653 ( .A(n584), .B(KEYINPUT12), .ZN(n586) );
  NAND2_X1 U654 ( .A1(G68), .A2(n653), .ZN(n585) );
  NAND2_X1 U655 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U656 ( .A(n587), .B(KEYINPUT13), .ZN(n589) );
  NAND2_X1 U657 ( .A1(G43), .A2(n650), .ZN(n588) );
  NAND2_X1 U658 ( .A1(n589), .A2(n588), .ZN(n592) );
  NAND2_X1 U659 ( .A1(n649), .A2(G56), .ZN(n590) );
  XOR2_X1 U660 ( .A(KEYINPUT14), .B(n590), .Z(n591) );
  NOR2_X1 U661 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U662 ( .A(KEYINPUT73), .B(n593), .ZN(n977) );
  INV_X1 U663 ( .A(n977), .ZN(n594) );
  NAND2_X1 U664 ( .A1(n594), .A2(G860), .ZN(G153) );
  INV_X1 U665 ( .A(G171), .ZN(G301) );
  NAND2_X1 U666 ( .A1(G868), .A2(G301), .ZN(n605) );
  NAND2_X1 U667 ( .A1(G66), .A2(n649), .ZN(n601) );
  NAND2_X1 U668 ( .A1(G79), .A2(n653), .ZN(n596) );
  NAND2_X1 U669 ( .A1(G92), .A2(n647), .ZN(n595) );
  NAND2_X1 U670 ( .A1(n596), .A2(n595), .ZN(n599) );
  NAND2_X1 U671 ( .A1(n650), .A2(G54), .ZN(n597) );
  XOR2_X1 U672 ( .A(KEYINPUT74), .B(n597), .Z(n598) );
  NOR2_X1 U673 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U674 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U675 ( .A(n602), .B(KEYINPUT15), .ZN(n603) );
  XOR2_X2 U676 ( .A(KEYINPUT75), .B(n603), .Z(n974) );
  OR2_X1 U677 ( .A1(n974), .A2(G868), .ZN(n604) );
  NAND2_X1 U678 ( .A1(n605), .A2(n604), .ZN(G284) );
  NAND2_X1 U679 ( .A1(n649), .A2(G65), .ZN(n606) );
  XNOR2_X1 U680 ( .A(n606), .B(KEYINPUT70), .ZN(n608) );
  NAND2_X1 U681 ( .A1(G53), .A2(n650), .ZN(n607) );
  NAND2_X1 U682 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U683 ( .A(KEYINPUT71), .B(n609), .ZN(n613) );
  NAND2_X1 U684 ( .A1(n653), .A2(G78), .ZN(n611) );
  NAND2_X1 U685 ( .A1(G91), .A2(n647), .ZN(n610) );
  AND2_X1 U686 ( .A1(n611), .A2(n610), .ZN(n612) );
  NAND2_X1 U687 ( .A1(n613), .A2(n612), .ZN(G299) );
  INV_X1 U688 ( .A(G868), .ZN(n670) );
  NOR2_X1 U689 ( .A1(G286), .A2(n670), .ZN(n615) );
  NOR2_X1 U690 ( .A1(G868), .A2(G299), .ZN(n614) );
  NOR2_X1 U691 ( .A1(n615), .A2(n614), .ZN(G297) );
  INV_X1 U692 ( .A(G559), .ZN(n616) );
  NOR2_X1 U693 ( .A1(G860), .A2(n616), .ZN(n617) );
  XNOR2_X1 U694 ( .A(KEYINPUT77), .B(n617), .ZN(n618) );
  NAND2_X1 U695 ( .A1(n618), .A2(n974), .ZN(n619) );
  XNOR2_X1 U696 ( .A(n619), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U697 ( .A1(G868), .A2(n977), .ZN(n620) );
  XNOR2_X1 U698 ( .A(KEYINPUT78), .B(n620), .ZN(n623) );
  NAND2_X1 U699 ( .A1(G868), .A2(n974), .ZN(n621) );
  NOR2_X1 U700 ( .A1(G559), .A2(n621), .ZN(n622) );
  NOR2_X1 U701 ( .A1(n623), .A2(n622), .ZN(G282) );
  NAND2_X1 U702 ( .A1(G80), .A2(n653), .ZN(n625) );
  NAND2_X1 U703 ( .A1(G93), .A2(n647), .ZN(n624) );
  NAND2_X1 U704 ( .A1(n625), .A2(n624), .ZN(n628) );
  NAND2_X1 U705 ( .A1(G55), .A2(n650), .ZN(n626) );
  XNOR2_X1 U706 ( .A(KEYINPUT79), .B(n626), .ZN(n627) );
  NOR2_X1 U707 ( .A1(n628), .A2(n627), .ZN(n630) );
  NAND2_X1 U708 ( .A1(n649), .A2(G67), .ZN(n629) );
  NAND2_X1 U709 ( .A1(n630), .A2(n629), .ZN(n671) );
  NAND2_X1 U710 ( .A1(n974), .A2(G559), .ZN(n668) );
  XNOR2_X1 U711 ( .A(n977), .B(n668), .ZN(n631) );
  NOR2_X1 U712 ( .A1(G860), .A2(n631), .ZN(n632) );
  XOR2_X1 U713 ( .A(n671), .B(n632), .Z(G145) );
  NAND2_X1 U714 ( .A1(G74), .A2(G651), .ZN(n638) );
  NAND2_X1 U715 ( .A1(G49), .A2(n650), .ZN(n635) );
  NAND2_X1 U716 ( .A1(G87), .A2(n633), .ZN(n634) );
  NAND2_X1 U717 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U718 ( .A1(n649), .A2(n636), .ZN(n637) );
  NAND2_X1 U719 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U720 ( .A(n639), .B(KEYINPUT80), .ZN(G288) );
  NAND2_X1 U721 ( .A1(G86), .A2(n647), .ZN(n641) );
  NAND2_X1 U722 ( .A1(G48), .A2(n650), .ZN(n640) );
  NAND2_X1 U723 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U724 ( .A1(n653), .A2(G73), .ZN(n642) );
  XOR2_X1 U725 ( .A(KEYINPUT2), .B(n642), .Z(n643) );
  NOR2_X1 U726 ( .A1(n644), .A2(n643), .ZN(n646) );
  NAND2_X1 U727 ( .A1(n649), .A2(G61), .ZN(n645) );
  NAND2_X1 U728 ( .A1(n646), .A2(n645), .ZN(G305) );
  NAND2_X1 U729 ( .A1(G85), .A2(n647), .ZN(n648) );
  XNOR2_X1 U730 ( .A(n648), .B(KEYINPUT66), .ZN(n658) );
  NAND2_X1 U731 ( .A1(G60), .A2(n649), .ZN(n652) );
  NAND2_X1 U732 ( .A1(G47), .A2(n650), .ZN(n651) );
  NAND2_X1 U733 ( .A1(n652), .A2(n651), .ZN(n656) );
  NAND2_X1 U734 ( .A1(G72), .A2(n653), .ZN(n654) );
  XNOR2_X1 U735 ( .A(KEYINPUT67), .B(n654), .ZN(n655) );
  NOR2_X1 U736 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U737 ( .A1(n658), .A2(n657), .ZN(G290) );
  XOR2_X1 U738 ( .A(KEYINPUT82), .B(KEYINPUT83), .Z(n660) );
  XNOR2_X1 U739 ( .A(KEYINPUT19), .B(KEYINPUT81), .ZN(n659) );
  XNOR2_X1 U740 ( .A(n660), .B(n659), .ZN(n663) );
  XNOR2_X1 U741 ( .A(G166), .B(G305), .ZN(n661) );
  XNOR2_X1 U742 ( .A(n661), .B(G290), .ZN(n662) );
  XNOR2_X1 U743 ( .A(n663), .B(n662), .ZN(n665) );
  INV_X1 U744 ( .A(G299), .ZN(n966) );
  XNOR2_X1 U745 ( .A(n977), .B(n966), .ZN(n664) );
  XNOR2_X1 U746 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U747 ( .A(G288), .B(n666), .ZN(n667) );
  XNOR2_X1 U748 ( .A(n667), .B(n671), .ZN(n903) );
  XNOR2_X1 U749 ( .A(n903), .B(n668), .ZN(n669) );
  NOR2_X1 U750 ( .A1(n670), .A2(n669), .ZN(n673) );
  NOR2_X1 U751 ( .A1(G868), .A2(n671), .ZN(n672) );
  NOR2_X1 U752 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U753 ( .A(KEYINPUT84), .B(n674), .ZN(G295) );
  NAND2_X1 U754 ( .A1(G2084), .A2(G2078), .ZN(n675) );
  XNOR2_X1 U755 ( .A(n675), .B(KEYINPUT20), .ZN(n676) );
  XNOR2_X1 U756 ( .A(KEYINPUT85), .B(n676), .ZN(n677) );
  NAND2_X1 U757 ( .A1(n677), .A2(G2090), .ZN(n678) );
  XNOR2_X1 U758 ( .A(KEYINPUT21), .B(n678), .ZN(n679) );
  NAND2_X1 U759 ( .A1(n679), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U760 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U761 ( .A(KEYINPUT72), .B(G82), .Z(G220) );
  NOR2_X1 U762 ( .A1(G236), .A2(G238), .ZN(n681) );
  NOR2_X1 U763 ( .A1(G235), .A2(G237), .ZN(n680) );
  NAND2_X1 U764 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U765 ( .A(KEYINPUT88), .B(n682), .ZN(n913) );
  NAND2_X1 U766 ( .A1(n913), .A2(G567), .ZN(n683) );
  XOR2_X1 U767 ( .A(KEYINPUT89), .B(n683), .Z(n690) );
  NOR2_X1 U768 ( .A1(G220), .A2(G219), .ZN(n684) );
  XOR2_X1 U769 ( .A(KEYINPUT86), .B(n684), .Z(n685) );
  XNOR2_X1 U770 ( .A(n685), .B(KEYINPUT22), .ZN(n686) );
  NOR2_X1 U771 ( .A1(G218), .A2(n686), .ZN(n687) );
  NAND2_X1 U772 ( .A1(G96), .A2(n687), .ZN(n912) );
  NAND2_X1 U773 ( .A1(G2106), .A2(n912), .ZN(n688) );
  XOR2_X1 U774 ( .A(KEYINPUT87), .B(n688), .Z(n689) );
  NAND2_X1 U775 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U776 ( .A(n691), .B(KEYINPUT90), .ZN(n906) );
  NAND2_X1 U777 ( .A1(G661), .A2(G483), .ZN(n692) );
  NOR2_X1 U778 ( .A1(n906), .A2(n692), .ZN(n834) );
  NAND2_X1 U779 ( .A1(G36), .A2(n834), .ZN(n693) );
  XOR2_X1 U780 ( .A(KEYINPUT91), .B(n693), .Z(G176) );
  INV_X1 U781 ( .A(G166), .ZN(G303) );
  XOR2_X1 U782 ( .A(KEYINPUT93), .B(G1986), .Z(n694) );
  XNOR2_X1 U783 ( .A(G290), .B(n694), .ZN(n976) );
  NOR2_X2 U784 ( .A1(G164), .A2(G1384), .ZN(n717) );
  NOR2_X1 U785 ( .A1(n717), .A2(n716), .ZN(n826) );
  NAND2_X1 U786 ( .A1(n976), .A2(n826), .ZN(n695) );
  XNOR2_X1 U787 ( .A(n695), .B(KEYINPUT94), .ZN(n715) );
  NAND2_X1 U788 ( .A1(G95), .A2(n886), .ZN(n697) );
  NAND2_X1 U789 ( .A1(G131), .A2(n889), .ZN(n696) );
  NAND2_X1 U790 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U791 ( .A(KEYINPUT95), .B(n698), .ZN(n702) );
  NAND2_X1 U792 ( .A1(n881), .A2(G107), .ZN(n700) );
  NAND2_X1 U793 ( .A1(G119), .A2(n882), .ZN(n699) );
  AND2_X1 U794 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U795 ( .A1(n702), .A2(n701), .ZN(n875) );
  NAND2_X1 U796 ( .A1(G1991), .A2(n875), .ZN(n713) );
  NAND2_X1 U797 ( .A1(G105), .A2(n886), .ZN(n703) );
  XNOR2_X1 U798 ( .A(n703), .B(KEYINPUT38), .ZN(n711) );
  NAND2_X1 U799 ( .A1(G129), .A2(n882), .ZN(n704) );
  XNOR2_X1 U800 ( .A(n704), .B(KEYINPUT96), .ZN(n706) );
  NAND2_X1 U801 ( .A1(n881), .A2(G117), .ZN(n705) );
  NAND2_X1 U802 ( .A1(n706), .A2(n705), .ZN(n709) );
  NAND2_X1 U803 ( .A1(G141), .A2(n889), .ZN(n707) );
  XNOR2_X1 U804 ( .A(KEYINPUT97), .B(n707), .ZN(n708) );
  NOR2_X1 U805 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U806 ( .A1(n711), .A2(n710), .ZN(n873) );
  NAND2_X1 U807 ( .A1(G1996), .A2(n873), .ZN(n712) );
  NAND2_X1 U808 ( .A1(n713), .A2(n712), .ZN(n933) );
  NAND2_X1 U809 ( .A1(n933), .A2(n826), .ZN(n714) );
  NAND2_X1 U810 ( .A1(n715), .A2(n714), .ZN(n806) );
  INV_X1 U811 ( .A(n716), .ZN(n718) );
  NAND2_X1 U812 ( .A1(n718), .A2(n717), .ZN(n721) );
  NAND2_X1 U813 ( .A1(G8), .A2(n764), .ZN(n799) );
  NOR2_X1 U814 ( .A1(G1981), .A2(G305), .ZN(n719) );
  XOR2_X1 U815 ( .A(n719), .B(KEYINPUT24), .Z(n720) );
  NOR2_X1 U816 ( .A1(n799), .A2(n720), .ZN(n804) );
  NOR2_X1 U817 ( .A1(G1976), .A2(G288), .ZN(n971) );
  INV_X1 U818 ( .A(n721), .ZN(n748) );
  NAND2_X1 U819 ( .A1(G1996), .A2(n748), .ZN(n723) );
  NAND2_X1 U820 ( .A1(G1341), .A2(n764), .ZN(n724) );
  XOR2_X1 U821 ( .A(KEYINPUT101), .B(n724), .Z(n725) );
  NAND2_X1 U822 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U823 ( .A1(n730), .A2(n974), .ZN(n729) );
  INV_X1 U824 ( .A(KEYINPUT102), .ZN(n728) );
  XNOR2_X1 U825 ( .A(n729), .B(n728), .ZN(n736) );
  NAND2_X1 U826 ( .A1(n974), .A2(n730), .ZN(n734) );
  NAND2_X1 U827 ( .A1(G1348), .A2(n764), .ZN(n732) );
  XNOR2_X1 U828 ( .A(n748), .B(KEYINPUT100), .ZN(n750) );
  NAND2_X1 U829 ( .A1(G2067), .A2(n750), .ZN(n731) );
  NAND2_X1 U830 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U831 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U832 ( .A1(n736), .A2(n735), .ZN(n741) );
  NAND2_X1 U833 ( .A1(G2072), .A2(n750), .ZN(n737) );
  XNOR2_X1 U834 ( .A(n737), .B(KEYINPUT27), .ZN(n739) );
  INV_X1 U835 ( .A(G1956), .ZN(n995) );
  NOR2_X1 U836 ( .A1(n750), .A2(n995), .ZN(n738) );
  NOR2_X1 U837 ( .A1(n739), .A2(n738), .ZN(n743) );
  NAND2_X1 U838 ( .A1(n966), .A2(n743), .ZN(n740) );
  NAND2_X1 U839 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U840 ( .A(KEYINPUT103), .B(n742), .ZN(n746) );
  OR2_X1 U841 ( .A1(n966), .A2(n743), .ZN(n744) );
  XOR2_X1 U842 ( .A(KEYINPUT28), .B(n744), .Z(n745) );
  NOR2_X1 U843 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U844 ( .A(KEYINPUT29), .B(n747), .ZN(n754) );
  XNOR2_X1 U845 ( .A(G1961), .B(KEYINPUT98), .ZN(n993) );
  NOR2_X1 U846 ( .A1(n748), .A2(n993), .ZN(n749) );
  XNOR2_X1 U847 ( .A(n749), .B(KEYINPUT99), .ZN(n752) );
  XNOR2_X1 U848 ( .A(G2078), .B(KEYINPUT25), .ZN(n946) );
  NAND2_X1 U849 ( .A1(n750), .A2(n946), .ZN(n751) );
  NAND2_X1 U850 ( .A1(n752), .A2(n751), .ZN(n755) );
  NAND2_X1 U851 ( .A1(n755), .A2(G171), .ZN(n753) );
  NAND2_X1 U852 ( .A1(n754), .A2(n753), .ZN(n763) );
  NOR2_X1 U853 ( .A1(G171), .A2(n755), .ZN(n760) );
  NOR2_X1 U854 ( .A1(G1966), .A2(n799), .ZN(n775) );
  NOR2_X1 U855 ( .A1(G2084), .A2(n764), .ZN(n772) );
  NOR2_X1 U856 ( .A1(n775), .A2(n772), .ZN(n756) );
  NAND2_X1 U857 ( .A1(G8), .A2(n756), .ZN(n757) );
  XNOR2_X1 U858 ( .A(KEYINPUT30), .B(n757), .ZN(n758) );
  NOR2_X1 U859 ( .A1(G168), .A2(n758), .ZN(n759) );
  NOR2_X1 U860 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U861 ( .A(KEYINPUT31), .B(n761), .Z(n762) );
  NAND2_X1 U862 ( .A1(n763), .A2(n762), .ZN(n773) );
  NAND2_X1 U863 ( .A1(n773), .A2(G286), .ZN(n769) );
  NOR2_X1 U864 ( .A1(G1971), .A2(n799), .ZN(n766) );
  NOR2_X1 U865 ( .A1(G2090), .A2(n764), .ZN(n765) );
  NOR2_X1 U866 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U867 ( .A1(n767), .A2(G303), .ZN(n768) );
  NAND2_X1 U868 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U869 ( .A1(n770), .A2(G8), .ZN(n771) );
  XNOR2_X1 U870 ( .A(n771), .B(KEYINPUT32), .ZN(n779) );
  NAND2_X1 U871 ( .A1(G8), .A2(n772), .ZN(n777) );
  INV_X1 U872 ( .A(n773), .ZN(n774) );
  NOR2_X1 U873 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U874 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U875 ( .A1(n779), .A2(n778), .ZN(n798) );
  NOR2_X1 U876 ( .A1(G1971), .A2(G303), .ZN(n780) );
  XOR2_X1 U877 ( .A(n780), .B(KEYINPUT104), .Z(n781) );
  NAND2_X1 U878 ( .A1(n798), .A2(n781), .ZN(n782) );
  NOR2_X1 U879 ( .A1(n782), .A2(KEYINPUT33), .ZN(n783) );
  NOR2_X1 U880 ( .A1(KEYINPUT105), .A2(n783), .ZN(n784) );
  NOR2_X1 U881 ( .A1(n971), .A2(n784), .ZN(n792) );
  NAND2_X1 U882 ( .A1(G1976), .A2(G288), .ZN(n972) );
  NOR2_X1 U883 ( .A1(KEYINPUT105), .A2(n799), .ZN(n787) );
  NAND2_X1 U884 ( .A1(n972), .A2(n787), .ZN(n786) );
  INV_X1 U885 ( .A(KEYINPUT33), .ZN(n785) );
  NAND2_X1 U886 ( .A1(n786), .A2(n785), .ZN(n790) );
  AND2_X1 U887 ( .A1(n971), .A2(KEYINPUT33), .ZN(n788) );
  NAND2_X1 U888 ( .A1(n788), .A2(n787), .ZN(n789) );
  NAND2_X1 U889 ( .A1(n790), .A2(n789), .ZN(n791) );
  NOR2_X1 U890 ( .A1(n792), .A2(n791), .ZN(n795) );
  XNOR2_X1 U891 ( .A(G1981), .B(G305), .ZN(n964) );
  AND2_X1 U892 ( .A1(n799), .A2(KEYINPUT105), .ZN(n793) );
  NOR2_X1 U893 ( .A1(n964), .A2(n793), .ZN(n794) );
  NAND2_X1 U894 ( .A1(n795), .A2(n794), .ZN(n802) );
  NOR2_X1 U895 ( .A1(G2090), .A2(G303), .ZN(n796) );
  NAND2_X1 U896 ( .A1(G8), .A2(n796), .ZN(n797) );
  NAND2_X1 U897 ( .A1(n798), .A2(n797), .ZN(n800) );
  NAND2_X1 U898 ( .A1(n800), .A2(n799), .ZN(n801) );
  NAND2_X1 U899 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR2_X1 U900 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U901 ( .A1(n806), .A2(n805), .ZN(n816) );
  NAND2_X1 U902 ( .A1(G104), .A2(n886), .ZN(n808) );
  NAND2_X1 U903 ( .A1(G140), .A2(n889), .ZN(n807) );
  NAND2_X1 U904 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U905 ( .A(KEYINPUT34), .B(n809), .ZN(n814) );
  NAND2_X1 U906 ( .A1(G116), .A2(n881), .ZN(n811) );
  NAND2_X1 U907 ( .A1(G128), .A2(n882), .ZN(n810) );
  NAND2_X1 U908 ( .A1(n811), .A2(n810), .ZN(n812) );
  XOR2_X1 U909 ( .A(KEYINPUT35), .B(n812), .Z(n813) );
  NOR2_X1 U910 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U911 ( .A(KEYINPUT36), .B(n815), .ZN(n897) );
  XNOR2_X1 U912 ( .A(G2067), .B(KEYINPUT37), .ZN(n823) );
  NOR2_X1 U913 ( .A1(n897), .A2(n823), .ZN(n914) );
  NAND2_X1 U914 ( .A1(n826), .A2(n914), .ZN(n821) );
  NAND2_X1 U915 ( .A1(n816), .A2(n821), .ZN(n829) );
  NOR2_X1 U916 ( .A1(G1996), .A2(n873), .ZN(n922) );
  NOR2_X1 U917 ( .A1(G1986), .A2(G290), .ZN(n817) );
  NOR2_X1 U918 ( .A1(G1991), .A2(n875), .ZN(n929) );
  NOR2_X1 U919 ( .A1(n817), .A2(n929), .ZN(n818) );
  NOR2_X1 U920 ( .A1(n933), .A2(n818), .ZN(n819) );
  NOR2_X1 U921 ( .A1(n922), .A2(n819), .ZN(n820) );
  XNOR2_X1 U922 ( .A(KEYINPUT39), .B(n820), .ZN(n822) );
  NAND2_X1 U923 ( .A1(n822), .A2(n821), .ZN(n824) );
  NAND2_X1 U924 ( .A1(n897), .A2(n823), .ZN(n915) );
  NAND2_X1 U925 ( .A1(n824), .A2(n915), .ZN(n825) );
  XNOR2_X1 U926 ( .A(KEYINPUT106), .B(n825), .ZN(n827) );
  NAND2_X1 U927 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U928 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U929 ( .A(n830), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U930 ( .A1(G2106), .A2(n831), .ZN(G217) );
  AND2_X1 U931 ( .A1(G15), .A2(G2), .ZN(n832) );
  NAND2_X1 U932 ( .A1(G661), .A2(n832), .ZN(G259) );
  NAND2_X1 U933 ( .A1(G3), .A2(G1), .ZN(n833) );
  NAND2_X1 U934 ( .A1(n834), .A2(n833), .ZN(G188) );
  XOR2_X1 U935 ( .A(G96), .B(KEYINPUT108), .Z(G221) );
  XOR2_X1 U936 ( .A(KEYINPUT112), .B(G2678), .Z(n836) );
  XNOR2_X1 U937 ( .A(KEYINPUT43), .B(G2100), .ZN(n835) );
  XNOR2_X1 U938 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U939 ( .A(n837), .B(KEYINPUT111), .Z(n839) );
  XNOR2_X1 U940 ( .A(G2067), .B(G2090), .ZN(n838) );
  XNOR2_X1 U941 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U942 ( .A(G2096), .B(G2084), .Z(n841) );
  XNOR2_X1 U943 ( .A(G2078), .B(G2072), .ZN(n840) );
  XNOR2_X1 U944 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U945 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U946 ( .A(KEYINPUT110), .B(KEYINPUT42), .ZN(n844) );
  XNOR2_X1 U947 ( .A(n845), .B(n844), .ZN(G227) );
  XOR2_X1 U948 ( .A(G1991), .B(G1976), .Z(n847) );
  XNOR2_X1 U949 ( .A(G1996), .B(G1956), .ZN(n846) );
  XNOR2_X1 U950 ( .A(n847), .B(n846), .ZN(n857) );
  XOR2_X1 U951 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n849) );
  XNOR2_X1 U952 ( .A(G1971), .B(KEYINPUT41), .ZN(n848) );
  XNOR2_X1 U953 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U954 ( .A(G1986), .B(G1981), .Z(n851) );
  XNOR2_X1 U955 ( .A(G1966), .B(G1961), .ZN(n850) );
  XNOR2_X1 U956 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U957 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U958 ( .A(KEYINPUT115), .B(G2474), .ZN(n854) );
  XNOR2_X1 U959 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U960 ( .A(n857), .B(n856), .Z(G229) );
  NAND2_X1 U961 ( .A1(G100), .A2(n886), .ZN(n859) );
  NAND2_X1 U962 ( .A1(G112), .A2(n881), .ZN(n858) );
  NAND2_X1 U963 ( .A1(n859), .A2(n858), .ZN(n865) );
  NAND2_X1 U964 ( .A1(G124), .A2(n882), .ZN(n860) );
  XNOR2_X1 U965 ( .A(n860), .B(KEYINPUT44), .ZN(n863) );
  NAND2_X1 U966 ( .A1(G136), .A2(n889), .ZN(n861) );
  XNOR2_X1 U967 ( .A(n861), .B(KEYINPUT116), .ZN(n862) );
  NAND2_X1 U968 ( .A1(n863), .A2(n862), .ZN(n864) );
  NOR2_X1 U969 ( .A1(n865), .A2(n864), .ZN(G162) );
  NAND2_X1 U970 ( .A1(G118), .A2(n881), .ZN(n867) );
  NAND2_X1 U971 ( .A1(G130), .A2(n882), .ZN(n866) );
  NAND2_X1 U972 ( .A1(n867), .A2(n866), .ZN(n872) );
  NAND2_X1 U973 ( .A1(G106), .A2(n886), .ZN(n869) );
  NAND2_X1 U974 ( .A1(G142), .A2(n889), .ZN(n868) );
  NAND2_X1 U975 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U976 ( .A(n870), .B(KEYINPUT45), .Z(n871) );
  NOR2_X1 U977 ( .A1(n872), .A2(n871), .ZN(n874) );
  XNOR2_X1 U978 ( .A(n874), .B(n873), .ZN(n896) );
  XNOR2_X1 U979 ( .A(G160), .B(n875), .ZN(n876) );
  XNOR2_X1 U980 ( .A(n876), .B(n930), .ZN(n880) );
  XOR2_X1 U981 ( .A(KEYINPUT48), .B(KEYINPUT119), .Z(n878) );
  XNOR2_X1 U982 ( .A(KEYINPUT46), .B(KEYINPUT118), .ZN(n877) );
  XNOR2_X1 U983 ( .A(n878), .B(n877), .ZN(n879) );
  XOR2_X1 U984 ( .A(n880), .B(n879), .Z(n894) );
  NAND2_X1 U985 ( .A1(G115), .A2(n881), .ZN(n884) );
  NAND2_X1 U986 ( .A1(G127), .A2(n882), .ZN(n883) );
  NAND2_X1 U987 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U988 ( .A(n885), .B(KEYINPUT47), .ZN(n888) );
  NAND2_X1 U989 ( .A1(G103), .A2(n886), .ZN(n887) );
  NAND2_X1 U990 ( .A1(n888), .A2(n887), .ZN(n892) );
  NAND2_X1 U991 ( .A1(G139), .A2(n889), .ZN(n890) );
  XNOR2_X1 U992 ( .A(KEYINPUT117), .B(n890), .ZN(n891) );
  NOR2_X1 U993 ( .A1(n892), .A2(n891), .ZN(n917) );
  XNOR2_X1 U994 ( .A(G164), .B(n917), .ZN(n893) );
  XNOR2_X1 U995 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U996 ( .A(n896), .B(n895), .ZN(n899) );
  XNOR2_X1 U997 ( .A(n897), .B(G162), .ZN(n898) );
  XNOR2_X1 U998 ( .A(n899), .B(n898), .ZN(n900) );
  NOR2_X1 U999 ( .A1(G37), .A2(n900), .ZN(G395) );
  XOR2_X1 U1000 ( .A(KEYINPUT120), .B(G286), .Z(n902) );
  XNOR2_X1 U1001 ( .A(G171), .B(n974), .ZN(n901) );
  XNOR2_X1 U1002 ( .A(n902), .B(n901), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n905), .ZN(G397) );
  XNOR2_X1 U1005 ( .A(KEYINPUT109), .B(n906), .ZN(G319) );
  NOR2_X1 U1006 ( .A1(G227), .A2(G229), .ZN(n907) );
  XNOR2_X1 U1007 ( .A(KEYINPUT49), .B(n907), .ZN(n908) );
  NOR2_X1 U1008 ( .A1(G401), .A2(n908), .ZN(n910) );
  NOR2_X1 U1009 ( .A1(G395), .A2(G397), .ZN(n909) );
  AND2_X1 U1010 ( .A1(n910), .A2(n909), .ZN(n911) );
  NAND2_X1 U1011 ( .A1(n911), .A2(G319), .ZN(G225) );
  XNOR2_X1 U1012 ( .A(KEYINPUT121), .B(G225), .ZN(G308) );
  NOR2_X1 U1014 ( .A1(n913), .A2(n912), .ZN(G325) );
  INV_X1 U1015 ( .A(G325), .ZN(G261) );
  INV_X1 U1016 ( .A(KEYINPUT55), .ZN(n959) );
  INV_X1 U1017 ( .A(n914), .ZN(n916) );
  NAND2_X1 U1018 ( .A1(n916), .A2(n915), .ZN(n927) );
  XOR2_X1 U1019 ( .A(G2072), .B(n917), .Z(n919) );
  XOR2_X1 U1020 ( .A(G164), .B(G2078), .Z(n918) );
  NOR2_X1 U1021 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1022 ( .A(KEYINPUT50), .B(n920), .ZN(n925) );
  XOR2_X1 U1023 ( .A(G2090), .B(G162), .Z(n921) );
  NOR2_X1 U1024 ( .A1(n922), .A2(n921), .ZN(n923) );
  XOR2_X1 U1025 ( .A(KEYINPUT51), .B(n923), .Z(n924) );
  NAND2_X1 U1026 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1027 ( .A1(n927), .A2(n926), .ZN(n935) );
  XOR2_X1 U1028 ( .A(G2084), .B(G160), .Z(n928) );
  NOR2_X1 U1029 ( .A1(n929), .A2(n928), .ZN(n931) );
  NAND2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1033 ( .A(KEYINPUT122), .B(n936), .ZN(n937) );
  XOR2_X1 U1034 ( .A(KEYINPUT52), .B(n937), .Z(n938) );
  NAND2_X1 U1035 ( .A1(n959), .A2(n938), .ZN(n939) );
  NAND2_X1 U1036 ( .A1(n939), .A2(G29), .ZN(n1019) );
  XNOR2_X1 U1037 ( .A(KEYINPUT123), .B(G2090), .ZN(n940) );
  XNOR2_X1 U1038 ( .A(n940), .B(G35), .ZN(n957) );
  XNOR2_X1 U1039 ( .A(KEYINPUT54), .B(G34), .ZN(n941) );
  XNOR2_X1 U1040 ( .A(n941), .B(KEYINPUT124), .ZN(n942) );
  XNOR2_X1 U1041 ( .A(G2084), .B(n942), .ZN(n955) );
  XOR2_X1 U1042 ( .A(G1991), .B(G25), .Z(n943) );
  NAND2_X1 U1043 ( .A1(n943), .A2(G28), .ZN(n952) );
  XNOR2_X1 U1044 ( .A(G2067), .B(G26), .ZN(n945) );
  XNOR2_X1 U1045 ( .A(G33), .B(G2072), .ZN(n944) );
  NOR2_X1 U1046 ( .A1(n945), .A2(n944), .ZN(n950) );
  XOR2_X1 U1047 ( .A(n946), .B(G27), .Z(n948) );
  XNOR2_X1 U1048 ( .A(G1996), .B(G32), .ZN(n947) );
  NOR2_X1 U1049 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1050 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1051 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1052 ( .A(KEYINPUT53), .B(n953), .ZN(n954) );
  NOR2_X1 U1053 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1054 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1055 ( .A(n959), .B(n958), .ZN(n961) );
  INV_X1 U1056 ( .A(G29), .ZN(n960) );
  NAND2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1058 ( .A1(G11), .A2(n962), .ZN(n1017) );
  XNOR2_X1 U1059 ( .A(G16), .B(KEYINPUT56), .ZN(n987) );
  XOR2_X1 U1060 ( .A(G168), .B(G1966), .Z(n963) );
  NOR2_X1 U1061 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1062 ( .A(KEYINPUT57), .B(n965), .Z(n985) );
  XNOR2_X1 U1063 ( .A(G166), .B(G1971), .ZN(n969) );
  XNOR2_X1 U1064 ( .A(n966), .B(KEYINPUT125), .ZN(n967) );
  XNOR2_X1 U1065 ( .A(n967), .B(n995), .ZN(n968) );
  NAND2_X1 U1066 ( .A1(n969), .A2(n968), .ZN(n970) );
  NOR2_X1 U1067 ( .A1(n971), .A2(n970), .ZN(n973) );
  NAND2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n983) );
  XOR2_X1 U1069 ( .A(G1348), .B(n974), .Z(n975) );
  NOR2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n981) );
  XNOR2_X1 U1071 ( .A(G301), .B(G1961), .ZN(n979) );
  XNOR2_X1 U1072 ( .A(n977), .B(G1341), .ZN(n978) );
  NOR2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n1015) );
  INV_X1 U1078 ( .A(G16), .ZN(n1013) );
  XOR2_X1 U1079 ( .A(G1976), .B(G23), .Z(n989) );
  XOR2_X1 U1080 ( .A(G1971), .B(G22), .Z(n988) );
  NAND2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n991) );
  XNOR2_X1 U1082 ( .A(G24), .B(G1986), .ZN(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n992) );
  XOR2_X1 U1084 ( .A(KEYINPUT58), .B(n992), .Z(n1010) );
  XOR2_X1 U1085 ( .A(n993), .B(G5), .Z(n1005) );
  XOR2_X1 U1086 ( .A(G1348), .B(KEYINPUT59), .Z(n994) );
  XNOR2_X1 U1087 ( .A(G4), .B(n994), .ZN(n1002) );
  XOR2_X1 U1088 ( .A(G1341), .B(G19), .Z(n997) );
  XNOR2_X1 U1089 ( .A(n995), .B(G20), .ZN(n996) );
  NAND2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n999) );
  XNOR2_X1 U1091 ( .A(G6), .B(G1981), .ZN(n998) );
  NOR2_X1 U1092 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1093 ( .A(KEYINPUT126), .B(n1000), .Z(n1001) );
  NOR2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1095 ( .A(KEYINPUT60), .B(n1003), .ZN(n1004) );
  NAND2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(G21), .B(G1966), .ZN(n1006) );
  NOR2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1099 ( .A(KEYINPUT127), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1101 ( .A(KEYINPUT61), .B(n1011), .ZN(n1012) );
  NAND2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XOR2_X1 U1106 ( .A(KEYINPUT62), .B(n1020), .Z(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

