//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 1 0 1 1 0 1 0 0 1 0 1 0 0 1 0 1 1 0 1 0 0 0 0 1 1 0 1 1 0 1 0 0 0 1 0 0 1 1 1 0 1 1 1 0 1 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n821, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1055, new_n1056, new_n1057, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101;
  INV_X1    g000(.A(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G125), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G140), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT16), .ZN(new_n191));
  OR3_X1    g005(.A1(new_n189), .A2(KEYINPUT16), .A3(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT76), .ZN(new_n194));
  NOR3_X1   g008(.A1(new_n189), .A2(KEYINPUT16), .A3(G140), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(KEYINPUT76), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(G146), .A3(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT78), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  AND3_X1   g014(.A1(new_n188), .A2(new_n190), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G119), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G128), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G119), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT24), .B(G110), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT23), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n209), .B1(new_n202), .B2(G128), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n204), .A2(KEYINPUT23), .A3(G119), .ZN(new_n211));
  INV_X1    g025(.A(G110), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n210), .A2(new_n211), .A3(new_n212), .A4(new_n203), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n208), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT77), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT77), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n208), .A2(new_n213), .A3(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n201), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT76), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n219), .B1(new_n191), .B2(new_n192), .ZN(new_n220));
  NOR3_X1   g034(.A1(new_n220), .A2(new_n200), .A3(new_n196), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT78), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n199), .A2(new_n218), .A3(new_n223), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n206), .A2(new_n207), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n210), .A2(new_n203), .A3(new_n211), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n225), .B1(G110), .B2(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(G146), .B1(new_n194), .B2(new_n197), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n227), .B1(new_n228), .B2(new_n221), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n224), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT80), .ZN(new_n231));
  INV_X1    g045(.A(G137), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT22), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT22), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G137), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT79), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n233), .A2(new_n235), .A3(KEYINPUT79), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n231), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  AND2_X1   g055(.A1(KEYINPUT69), .A2(G953), .ZN(new_n242));
  NOR2_X1   g056(.A1(KEYINPUT69), .A2(G953), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G221), .ZN(new_n246));
  INV_X1    g060(.A(G234), .ZN(new_n247));
  NOR3_X1   g061(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n238), .A2(new_n239), .A3(new_n231), .ZN(new_n249));
  AND3_X1   g063(.A1(new_n241), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n248), .B1(new_n241), .B2(new_n249), .ZN(new_n251));
  OR2_X1    g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n230), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT72), .B(G902), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n250), .A2(new_n251), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n255), .A2(new_n224), .A3(new_n229), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n253), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n258), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n253), .A2(new_n254), .A3(new_n256), .A4(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G217), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n263), .B1(new_n254), .B2(G234), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n264), .B(KEYINPUT75), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n262), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n253), .A2(new_n256), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n264), .A2(G902), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n272), .B(KEYINPUT82), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT65), .ZN(new_n274));
  AND3_X1   g088(.A1(new_n200), .A2(KEYINPUT64), .A3(G143), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n200), .A2(G143), .ZN(new_n276));
  OAI21_X1  g090(.A(KEYINPUT64), .B1(new_n200), .B2(G143), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(KEYINPUT0), .B(G128), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n274), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT11), .ZN(new_n281));
  INV_X1    g095(.A(G134), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n281), .B1(new_n282), .B2(G137), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n232), .A2(KEYINPUT11), .A3(G134), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(G137), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(G131), .ZN(new_n287));
  XNOR2_X1  g101(.A(KEYINPUT66), .B(G131), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n288), .A2(new_n283), .A3(new_n284), .A4(new_n285), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n277), .A2(new_n276), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n200), .A2(KEYINPUT64), .A3(G143), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n279), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n293), .A2(KEYINPUT65), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G143), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G146), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n276), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n298), .A2(KEYINPUT0), .A3(G128), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n280), .A2(new_n290), .A3(new_n295), .A4(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n202), .A2(G116), .ZN(new_n301));
  INV_X1    g115(.A(G116), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G119), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT2), .B(G113), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G113), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT2), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT2), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G113), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(G116), .B(G119), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT67), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n313), .B1(new_n311), .B2(new_n312), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n306), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT68), .ZN(new_n317));
  INV_X1    g131(.A(new_n285), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n282), .A2(G137), .ZN(new_n319));
  OAI21_X1  g133(.A(G131), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n204), .B1(new_n276), .B2(KEYINPUT1), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n321), .B1(new_n292), .B2(new_n291), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT1), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n276), .A2(new_n297), .A3(new_n323), .A4(G128), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n289), .B(new_n320), .C1(new_n322), .C2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(KEYINPUT67), .B1(new_n304), .B2(new_n305), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT68), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(new_n330), .A3(new_n306), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n300), .A2(new_n317), .A3(new_n326), .A4(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  AOI22_X1  g147(.A1(new_n300), .A2(new_n326), .B1(new_n317), .B2(new_n331), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT28), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT28), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT70), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT70), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n332), .A2(new_n339), .A3(new_n336), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n335), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G237), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n244), .A2(G210), .A3(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n343), .B(KEYINPUT27), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT26), .B(G101), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n344), .B(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT31), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n317), .A2(new_n331), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n300), .A2(new_n326), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT30), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT30), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n300), .A2(new_n354), .A3(new_n326), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n351), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n346), .A2(new_n332), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n349), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n300), .A2(new_n354), .A3(new_n326), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n354), .B1(new_n300), .B2(new_n326), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n350), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n361), .A2(KEYINPUT31), .A3(new_n346), .A4(new_n332), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT71), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n348), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n364), .B1(new_n348), .B2(new_n363), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT32), .ZN(new_n368));
  NOR3_X1   g182(.A1(new_n368), .A2(G472), .A3(G902), .ZN(new_n369));
  AOI21_X1  g183(.A(KEYINPUT74), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n348), .A2(new_n363), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(KEYINPUT71), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n348), .A2(new_n363), .A3(new_n364), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n372), .A2(KEYINPUT74), .A3(new_n373), .A4(new_n369), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n370), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g190(.A1(G472), .A2(G902), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n372), .A2(new_n377), .A3(new_n373), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n346), .A2(KEYINPUT29), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n254), .B1(new_n341), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT73), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI211_X1 g196(.A(KEYINPUT73), .B(new_n254), .C1(new_n341), .C2(new_n379), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT29), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n347), .B1(new_n356), .B2(new_n333), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n384), .B(new_n385), .C1(new_n341), .C2(new_n347), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n382), .A2(new_n383), .A3(new_n386), .ZN(new_n387));
  AOI22_X1  g201(.A1(new_n378), .A2(new_n368), .B1(new_n387), .B2(G472), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n273), .B1(new_n376), .B2(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n322), .A2(new_n325), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT10), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT85), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT84), .ZN(new_n394));
  INV_X1    g208(.A(G104), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(KEYINPUT84), .A2(G104), .ZN(new_n397));
  AOI21_X1  g211(.A(G107), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G107), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n399), .A2(G104), .ZN(new_n400));
  OAI21_X1  g214(.A(G101), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  NOR3_X1   g215(.A1(new_n395), .A2(KEYINPUT3), .A3(G107), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT3), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n403), .B1(new_n398), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n396), .A2(G107), .A3(new_n397), .ZN(new_n406));
  INV_X1    g220(.A(G101), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n393), .B(new_n401), .C1(new_n405), .C2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  AND2_X1   g224(.A1(KEYINPUT84), .A2(G104), .ZN(new_n411));
  NOR2_X1   g225(.A1(KEYINPUT84), .A2(G104), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n399), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n402), .B1(new_n413), .B2(KEYINPUT3), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n411), .A2(new_n412), .ZN(new_n415));
  AOI21_X1  g229(.A(G101), .B1(new_n415), .B2(G107), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n393), .B1(new_n417), .B2(new_n401), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n392), .B1(new_n410), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n279), .B1(new_n291), .B2(new_n292), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n299), .B1(new_n420), .B2(KEYINPUT65), .ZN(new_n421));
  NOR3_X1   g235(.A1(new_n278), .A2(new_n274), .A3(new_n279), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n403), .B(new_n406), .C1(new_n398), .C2(new_n404), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT4), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(new_n425), .A3(G101), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n425), .B1(new_n414), .B2(new_n416), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n424), .A2(G101), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n423), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n290), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n324), .B1(new_n298), .B2(new_n321), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n417), .A2(new_n401), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n391), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n419), .A2(new_n430), .A3(new_n431), .A4(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n244), .A2(G227), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n436), .B(KEYINPUT83), .ZN(new_n437));
  XNOR2_X1  g251(.A(G110), .B(G140), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n437), .B(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n435), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n419), .A2(new_n430), .A3(new_n434), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n290), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n435), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n401), .B1(new_n405), .B2(new_n408), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT85), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(new_n390), .A3(new_n409), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n433), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n290), .ZN(new_n450));
  AOI21_X1  g264(.A(KEYINPUT12), .B1(new_n290), .B2(KEYINPUT86), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n451), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n449), .A2(new_n290), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n445), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n444), .B1(new_n455), .B2(new_n440), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT87), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n453), .B1(new_n449), .B2(new_n290), .ZN(new_n458));
  AOI211_X1 g272(.A(new_n431), .B(new_n451), .C1(new_n448), .C2(new_n433), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n435), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AOI22_X1  g274(.A1(new_n460), .A2(new_n439), .B1(new_n443), .B2(new_n441), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT87), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n457), .A2(G469), .A3(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(G469), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n458), .A2(new_n459), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n435), .A2(KEYINPUT88), .A3(new_n440), .ZN(new_n467));
  AOI21_X1  g281(.A(KEYINPUT88), .B1(new_n435), .B2(new_n440), .ZN(new_n468));
  NOR3_X1   g282(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n440), .B1(new_n443), .B2(new_n435), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n465), .B(new_n254), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(G902), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n465), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n464), .A2(new_n471), .A3(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(KEYINPUT9), .B(G234), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n246), .B1(new_n477), .B2(new_n472), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(G113), .B(G122), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(new_n395), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n228), .A2(new_n221), .ZN(new_n483));
  OR2_X1    g297(.A1(KEYINPUT69), .A2(G953), .ZN(new_n484));
  NAND2_X1  g298(.A1(KEYINPUT69), .A2(G953), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n484), .A2(G214), .A3(new_n342), .A4(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n296), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n244), .A2(G143), .A3(G214), .A4(new_n342), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n288), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n489), .A2(KEYINPUT17), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n490), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n487), .A2(new_n488), .A3(new_n288), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n483), .B(new_n491), .C1(KEYINPUT17), .C2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(KEYINPUT18), .A2(G131), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n487), .A2(new_n488), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT93), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n487), .A2(new_n488), .A3(KEYINPUT93), .A4(new_n496), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n496), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n200), .B1(new_n188), .B2(new_n190), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(G125), .B(G140), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n200), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT92), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n504), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(KEYINPUT92), .B1(new_n201), .B2(new_n503), .ZN(new_n509));
  AOI22_X1  g323(.A1(new_n489), .A2(new_n502), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n501), .A2(KEYINPUT94), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(KEYINPUT94), .B1(new_n501), .B2(new_n510), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n482), .B(new_n495), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT96), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n501), .A2(new_n510), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT94), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n501), .A2(KEYINPUT94), .A3(new_n510), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n520), .A2(KEYINPUT96), .A3(new_n482), .A4(new_n495), .ZN(new_n521));
  INV_X1    g335(.A(new_n482), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT19), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n505), .B1(KEYINPUT95), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n524), .B1(new_n505), .B2(new_n525), .ZN(new_n526));
  OR2_X1    g340(.A1(new_n526), .A2(G146), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n494), .A2(new_n199), .A3(new_n223), .A4(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n520), .A2(new_n528), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n515), .A2(new_n521), .B1(new_n522), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(G475), .A2(G902), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(KEYINPUT20), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n529), .A2(new_n522), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT17), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n492), .A2(new_n535), .A3(new_n493), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n200), .B1(new_n220), .B2(new_n196), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n491), .A2(new_n537), .A3(new_n198), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n539), .B1(new_n518), .B2(new_n519), .ZN(new_n540));
  AOI21_X1  g354(.A(KEYINPUT96), .B1(new_n540), .B2(new_n482), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n513), .A2(new_n514), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n534), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OR2_X1    g357(.A1(new_n532), .A2(KEYINPUT97), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT20), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n532), .A2(KEYINPUT97), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n520), .A2(new_n495), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n522), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n550), .B1(new_n541), .B2(new_n542), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n472), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n533), .A2(new_n548), .B1(new_n552), .B2(G475), .ZN(new_n553));
  OAI21_X1  g367(.A(G214), .B1(G237), .B2(G902), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n311), .A2(new_n312), .ZN(new_n556));
  AOI211_X1 g370(.A(KEYINPUT68), .B(new_n556), .C1(new_n328), .C2(new_n327), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n330), .B1(new_n329), .B2(new_n306), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n426), .B(new_n429), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(G113), .B1(new_n301), .B2(KEYINPUT5), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n312), .A2(KEYINPUT5), .ZN(new_n562));
  AOI22_X1  g376(.A1(new_n327), .A2(new_n328), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n563), .B1(new_n410), .B2(new_n418), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(G110), .B(G122), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n559), .A2(new_n564), .A3(new_n566), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(KEYINPUT6), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT6), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n565), .A2(new_n571), .A3(new_n567), .ZN(new_n572));
  OAI21_X1  g386(.A(G125), .B1(new_n421), .B2(new_n422), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n390), .A2(new_n189), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  XOR2_X1   g389(.A(KEYINPUT89), .B(G224), .Z(new_n576));
  NOR2_X1   g390(.A1(new_n576), .A2(G953), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n575), .B(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n570), .A2(new_n572), .A3(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n566), .B(KEYINPUT8), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT90), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n562), .B1(new_n561), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n560), .A2(KEYINPUT90), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n329), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n584), .B1(new_n447), .B2(new_n409), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n563), .B1(new_n417), .B2(new_n401), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n580), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n587), .A2(new_n569), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n573), .A2(KEYINPUT91), .ZN(new_n589));
  OAI21_X1  g403(.A(KEYINPUT7), .B1(new_n576), .B2(G953), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n575), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n590), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n573), .B(new_n574), .C1(KEYINPUT91), .C2(new_n592), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(G902), .B1(new_n588), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n579), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(G210), .B1(G237), .B2(G902), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n579), .A2(new_n595), .A3(new_n597), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n555), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(G952), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n602), .A2(G953), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n603), .B1(new_n247), .B2(new_n342), .ZN(new_n604));
  AOI211_X1 g418(.A(new_n254), .B(new_n244), .C1(G234), .C2(G237), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT21), .B(G898), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n604), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n302), .A2(G122), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT98), .ZN(new_n611));
  INV_X1    g425(.A(G122), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n611), .B1(G116), .B2(new_n612), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n302), .A2(KEYINPUT98), .A3(G122), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n610), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(KEYINPUT14), .B1(new_n613), .B2(new_n614), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n615), .A2(new_n616), .A3(G107), .ZN(new_n617));
  OAI221_X1 g431(.A(new_n610), .B1(KEYINPUT14), .B2(new_n399), .C1(new_n613), .C2(new_n614), .ZN(new_n618));
  XNOR2_X1  g432(.A(G128), .B(G143), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT99), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n619), .A2(new_n620), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n622), .A2(new_n623), .A3(new_n282), .ZN(new_n624));
  OR2_X1    g438(.A1(new_n619), .A2(new_n620), .ZN(new_n625));
  AOI21_X1  g439(.A(G134), .B1(new_n625), .B2(new_n621), .ZN(new_n626));
  OAI211_X1 g440(.A(new_n617), .B(new_n618), .C1(new_n624), .C2(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n282), .B1(new_n622), .B2(new_n623), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n619), .A2(KEYINPUT13), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n296), .A2(G128), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n629), .B(G134), .C1(KEYINPUT13), .C2(new_n630), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n615), .A2(G107), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n615), .A2(G107), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n628), .B(new_n631), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n627), .A2(new_n634), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n476), .A2(new_n263), .A3(G953), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n627), .A2(new_n634), .A3(new_n636), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n638), .A2(KEYINPUT100), .A3(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT100), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n635), .A2(new_n641), .A3(new_n637), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n640), .A2(new_n254), .A3(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(G478), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n644), .A2(KEYINPUT15), .ZN(new_n645));
  OR2_X1    g459(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n643), .A2(new_n645), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n553), .A2(new_n601), .A3(new_n609), .A4(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n480), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n389), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G101), .ZN(G3));
  NAND3_X1  g467(.A1(new_n372), .A2(new_n373), .A3(new_n254), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT101), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT102), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n372), .A2(KEYINPUT101), .A3(new_n373), .A4(new_n254), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n656), .A2(new_n657), .A3(G472), .A4(new_n658), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n659), .A2(new_n378), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n656), .A2(G472), .A3(new_n658), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(KEYINPUT102), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n480), .A2(new_n273), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n660), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(new_n664), .B(KEYINPUT103), .Z(new_n665));
  INV_X1    g479(.A(KEYINPUT33), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n640), .A2(new_n666), .A3(new_n642), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n638), .A2(KEYINPUT33), .A3(new_n639), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n667), .A2(G478), .A3(new_n254), .A4(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n643), .A2(new_n644), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n515), .A2(new_n521), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n532), .B1(new_n672), .B2(new_n534), .ZN(new_n673));
  INV_X1    g487(.A(new_n547), .ZN(new_n674));
  OAI22_X1  g488(.A1(new_n673), .A2(new_n545), .B1(new_n530), .B2(new_n674), .ZN(new_n675));
  AOI22_X1  g489(.A1(new_n515), .A2(new_n521), .B1(new_n522), .B2(new_n549), .ZN(new_n676));
  OAI21_X1  g490(.A(G475), .B1(new_n676), .B2(G902), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n671), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n579), .A2(new_n595), .A3(new_n597), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n597), .B1(new_n579), .B2(new_n595), .ZN(new_n680));
  OAI211_X1 g494(.A(new_n609), .B(new_n554), .C1(new_n679), .C2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n665), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT34), .B(G104), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G6));
  NAND3_X1  g501(.A1(new_n543), .A2(new_n545), .A3(new_n531), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n533), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n689), .A2(new_n609), .A3(new_n677), .A4(new_n648), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT104), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n554), .B1(new_n679), .B2(new_n680), .ZN(new_n693));
  AND4_X1   g507(.A1(new_n609), .A2(new_n689), .A3(new_n677), .A4(new_n648), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n693), .B1(new_n694), .B2(KEYINPUT104), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n665), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT35), .B(G107), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G9));
  AOI21_X1  g512(.A(new_n265), .B1(new_n259), .B2(new_n261), .ZN(new_n699));
  INV_X1    g513(.A(new_n270), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n701), .B1(new_n224), .B2(new_n229), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  OR3_X1    g517(.A1(new_n250), .A2(new_n251), .A3(KEYINPUT36), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n224), .A2(new_n229), .A3(new_n701), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n703), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n224), .A2(new_n701), .A3(new_n229), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n704), .B1(new_n708), .B2(new_n702), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n700), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n699), .A2(new_n710), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n480), .A2(new_n650), .A3(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(new_n660), .A3(new_n662), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(KEYINPUT106), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT37), .B(G110), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G12));
  AOI221_X4 g530(.A(KEYINPUT87), .B1(new_n441), .B2(new_n443), .C1(new_n460), .C2(new_n439), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n460), .A2(new_n439), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n462), .B1(new_n718), .B2(new_n444), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n473), .B1(new_n720), .B2(G469), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n478), .B1(new_n721), .B2(new_n471), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n378), .A2(new_n368), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n372), .A2(new_n373), .A3(new_n369), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT74), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n387), .A2(G472), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n723), .A2(new_n726), .A3(new_n727), .A4(new_n374), .ZN(new_n728));
  AOI22_X1  g542(.A1(new_n688), .A2(new_n533), .B1(new_n552), .B2(G475), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n604), .B1(new_n606), .B2(G900), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(KEYINPUT107), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n729), .A2(new_n648), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  OR2_X1    g547(.A1(new_n699), .A2(new_n710), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n601), .A2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n722), .A2(new_n728), .A3(new_n733), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G128), .ZN(G30));
  NOR2_X1   g552(.A1(new_n356), .A2(new_n333), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n739), .A2(new_n347), .ZN(new_n740));
  OR2_X1    g554(.A1(new_n333), .A2(new_n334), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n472), .B1(new_n741), .B2(new_n346), .ZN(new_n742));
  OAI21_X1  g556(.A(G472), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(KEYINPUT108), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT108), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n745), .B(G472), .C1(new_n740), .C2(new_n742), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n723), .A2(new_n726), .A3(new_n748), .A4(new_n374), .ZN(new_n749));
  NOR4_X1   g563(.A1(new_n553), .A2(new_n555), .A3(new_n649), .A4(new_n734), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n679), .A2(new_n680), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(KEYINPUT38), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT38), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n753), .B1(new_n679), .B2(new_n680), .ZN(new_n754));
  AND4_X1   g568(.A1(new_n749), .A2(new_n750), .A3(new_n752), .A4(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n731), .B(KEYINPUT39), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n475), .A2(new_n479), .A3(new_n756), .ZN(new_n757));
  OR2_X1    g571(.A1(new_n757), .A2(KEYINPUT40), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(KEYINPUT40), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n755), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G143), .ZN(G45));
  INV_X1    g575(.A(new_n731), .ZN(new_n762));
  AOI211_X1 g576(.A(new_n671), .B(new_n762), .C1(new_n675), .C2(new_n677), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n722), .A2(new_n728), .A3(new_n736), .A4(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G146), .ZN(G48));
  NAND2_X1  g579(.A1(new_n435), .A2(new_n440), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT88), .ZN(new_n767));
  AOI22_X1  g581(.A1(new_n454), .A2(new_n452), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n435), .A2(KEYINPUT88), .A3(new_n440), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n470), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n254), .ZN(new_n771));
  OAI21_X1  g585(.A(G469), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(new_n479), .A3(new_n471), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT109), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n772), .A2(KEYINPUT109), .A3(new_n479), .A4(new_n471), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n389), .A2(new_n684), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(KEYINPUT41), .B(G113), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n778), .B(new_n779), .ZN(G15));
  INV_X1    g594(.A(KEYINPUT82), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n272), .B(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n728), .A2(new_n782), .A3(new_n775), .A4(new_n776), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n729), .A2(KEYINPUT104), .A3(new_n609), .A4(new_n648), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n692), .A2(new_n601), .A3(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(new_n302), .ZN(G18));
  NAND4_X1  g601(.A1(new_n675), .A2(new_n609), .A3(new_n677), .A4(new_n649), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(new_n773), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n728), .A2(new_n789), .A3(new_n736), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G119), .ZN(G21));
  NAND2_X1  g605(.A1(new_n452), .A2(new_n454), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n766), .A2(new_n767), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(new_n769), .A3(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n470), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n465), .B1(new_n796), .B2(new_n254), .ZN(new_n797));
  AOI211_X1 g611(.A(G469), .B(new_n771), .C1(new_n794), .C2(new_n795), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT109), .B1(new_n799), .B2(new_n479), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n545), .B1(new_n543), .B2(new_n531), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n530), .A2(new_n674), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n677), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n803), .A2(new_n601), .A3(new_n609), .A4(new_n648), .ZN(new_n804));
  INV_X1    g618(.A(new_n776), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n800), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n272), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n371), .A2(new_n377), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n365), .A2(new_n366), .A3(new_n771), .ZN(new_n809));
  INV_X1    g623(.A(G472), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n807), .B(new_n808), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT110), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n654), .A2(G472), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n814), .A2(KEYINPUT110), .A3(new_n807), .A4(new_n808), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n806), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G122), .ZN(G24));
  AND3_X1   g632(.A1(new_n814), .A2(new_n734), .A3(new_n808), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n773), .A2(new_n693), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n819), .A2(new_n763), .A3(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(G125), .ZN(G27));
  NOR3_X1   g636(.A1(new_n679), .A2(new_n680), .A3(new_n555), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n473), .B1(new_n461), .B2(G469), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n471), .A2(new_n824), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n823), .A2(new_n825), .A3(new_n479), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n728), .A2(new_n782), .A3(new_n763), .A4(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT42), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT111), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n826), .A2(new_n763), .A3(KEYINPUT42), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n723), .A2(new_n727), .A3(new_n724), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(new_n807), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n830), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n272), .B1(new_n388), .B2(new_n724), .ZN(new_n835));
  NOR4_X1   g649(.A1(new_n553), .A2(new_n828), .A3(new_n671), .A4(new_n762), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n835), .A2(KEYINPUT111), .A3(new_n836), .A4(new_n826), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n829), .A2(new_n834), .A3(new_n837), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(G131), .ZN(G33));
  NAND4_X1  g653(.A1(new_n728), .A2(new_n733), .A3(new_n782), .A4(new_n826), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(G134), .ZN(G36));
  NAND3_X1  g655(.A1(new_n662), .A2(new_n378), .A3(new_n659), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT43), .B1(new_n803), .B2(new_n671), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT43), .ZN(new_n844));
  INV_X1    g658(.A(new_n671), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n553), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n843), .A2(new_n846), .A3(new_n734), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n842), .A2(KEYINPUT44), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(new_n823), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT113), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n848), .A2(KEYINPUT113), .A3(new_n823), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n465), .B1(new_n461), .B2(KEYINPUT45), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n853), .B1(new_n720), .B2(KEYINPUT45), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n474), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT46), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT45), .B1(new_n457), .B2(new_n463), .ZN(new_n858));
  INV_X1    g672(.A(new_n853), .ZN(new_n859));
  OAI211_X1 g673(.A(KEYINPUT46), .B(new_n474), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT112), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n854), .A2(KEYINPUT112), .A3(KEYINPUT46), .A4(new_n474), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n857), .A2(new_n862), .A3(new_n471), .A4(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n864), .A2(new_n479), .A3(new_n756), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT44), .B1(new_n842), .B2(new_n847), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n851), .A2(new_n852), .A3(new_n867), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(G137), .ZN(G39));
  NAND2_X1  g683(.A1(new_n864), .A2(new_n479), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT47), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n864), .A2(KEYINPUT47), .A3(new_n479), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n763), .ZN(new_n875));
  INV_X1    g689(.A(new_n823), .ZN(new_n876));
  NOR4_X1   g690(.A1(new_n875), .A2(new_n728), .A3(new_n782), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(G140), .ZN(G42));
  INV_X1    g693(.A(KEYINPUT51), .ZN(new_n880));
  INV_X1    g694(.A(new_n604), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n843), .A2(new_n846), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n882), .B1(new_n813), .B2(new_n815), .ZN(new_n883));
  AOI211_X1 g697(.A(new_n554), .B(new_n773), .C1(new_n752), .C2(new_n754), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT50), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n882), .ZN(new_n886));
  AND4_X1   g700(.A1(KEYINPUT50), .A2(new_n886), .A3(new_n816), .A4(new_n884), .ZN(new_n887));
  OR2_X1    g701(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n747), .B1(new_n368), .B2(new_n378), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n376), .A2(new_n782), .A3(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n799), .A2(new_n479), .A3(new_n881), .A4(new_n823), .ZN(new_n891));
  OAI21_X1  g705(.A(KEYINPUT118), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n749), .ZN(new_n893));
  INV_X1    g707(.A(new_n891), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT118), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n893), .A2(new_n894), .A3(new_n895), .A4(new_n782), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n803), .A2(new_n845), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n892), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n843), .A2(new_n846), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n899), .A2(new_n819), .A3(new_n894), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n888), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n880), .B1(new_n902), .B2(KEYINPUT120), .ZN(new_n903));
  INV_X1    g717(.A(new_n799), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n904), .A2(new_n479), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT121), .B1(new_n874), .B2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT121), .ZN(new_n907));
  INV_X1    g721(.A(new_n905), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n872), .A2(new_n907), .A3(new_n873), .A4(new_n908), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n883), .A2(new_n823), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n906), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n903), .B(new_n911), .C1(KEYINPUT120), .C2(new_n902), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n899), .A2(new_n835), .A3(new_n894), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT48), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n883), .A2(new_n820), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n915), .A2(new_n603), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n892), .A2(new_n896), .A3(new_n678), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT122), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AND4_X1   g732(.A1(KEYINPUT122), .A2(new_n917), .A3(new_n603), .A4(new_n915), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n914), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n888), .A2(new_n901), .A3(KEYINPUT119), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n905), .B(KEYINPUT117), .Z(new_n922));
  OAI21_X1  g736(.A(new_n910), .B1(new_n874), .B2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT119), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n885), .A2(new_n887), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n898), .A2(new_n900), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n921), .A2(new_n923), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n920), .B1(new_n928), .B2(new_n880), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n912), .A2(new_n929), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n711), .A2(new_n648), .A3(new_n762), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n931), .A2(new_n729), .A3(new_n823), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n722), .A2(new_n728), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n819), .A2(new_n763), .A3(new_n826), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n840), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n838), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n553), .A2(new_n649), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n803), .A2(new_n671), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n937), .A2(new_n938), .A3(new_n682), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n660), .A2(new_n662), .A3(new_n663), .A4(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n940), .A2(new_n713), .A3(new_n652), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n389), .A2(new_n692), .A3(new_n695), .A4(new_n777), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n942), .A2(new_n778), .A3(new_n817), .A4(new_n790), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n936), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n478), .B1(new_n471), .B2(new_n824), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n553), .A2(new_n693), .A3(new_n649), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT115), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n947), .B1(new_n734), .B2(new_n762), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n711), .A2(KEYINPUT115), .A3(new_n731), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n749), .A2(new_n945), .A3(new_n946), .A4(new_n950), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n737), .A2(new_n764), .A3(new_n821), .A4(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(KEYINPUT52), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n735), .B1(new_n376), .B2(new_n388), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n480), .A2(new_n732), .ZN(new_n955));
  AND4_X1   g769(.A1(new_n479), .A2(new_n475), .A3(new_n678), .A4(new_n731), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT52), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n957), .A2(new_n958), .A3(new_n821), .A4(new_n951), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n953), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(KEYINPUT53), .B1(new_n944), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n840), .A2(new_n933), .A3(new_n934), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n835), .A2(new_n826), .A3(new_n836), .ZN(new_n963));
  AOI22_X1  g777(.A1(new_n830), .A2(new_n963), .B1(new_n827), .B2(new_n828), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n962), .B1(new_n964), .B2(new_n837), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n940), .A2(new_n713), .A3(new_n652), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n790), .B1(new_n783), .B2(new_n683), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n649), .B1(new_n675), .B2(new_n677), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n775), .A2(new_n682), .A3(new_n776), .A4(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n813), .B2(new_n815), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n967), .A2(new_n786), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n965), .A2(new_n966), .A3(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT53), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n953), .A2(new_n959), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(KEYINPUT54), .B1(new_n961), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n973), .B1(new_n972), .B2(new_n974), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n940), .A2(new_n713), .A3(KEYINPUT53), .A4(new_n652), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n936), .A2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n967), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT116), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n980), .A2(new_n981), .A3(new_n942), .A4(new_n817), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n943), .A2(KEYINPUT116), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n979), .A2(new_n960), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT54), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n977), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n976), .A2(new_n986), .ZN(new_n987));
  OAI22_X1  g801(.A1(new_n930), .A2(new_n987), .B1(G952), .B2(G953), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n807), .A2(new_n479), .A3(new_n554), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n989), .B(KEYINPUT114), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n990), .B1(new_n752), .B2(new_n754), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n803), .A2(new_n671), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n799), .B(KEYINPUT49), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n991), .A2(new_n893), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n988), .A2(new_n994), .ZN(G75));
  NAND2_X1  g809(.A1(new_n977), .A2(new_n984), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n996), .A2(new_n771), .A3(new_n598), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT56), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n570), .A2(new_n572), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(new_n578), .ZN(new_n1000));
  XOR2_X1   g814(.A(KEYINPUT123), .B(KEYINPUT55), .Z(new_n1001));
  XNOR2_X1  g815(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  AND3_X1   g816(.A1(new_n997), .A2(new_n998), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1002), .B1(new_n997), .B2(new_n998), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n244), .A2(G952), .ZN(new_n1005));
  NOR3_X1   g819(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(G51));
  XNOR2_X1  g820(.A(new_n473), .B(KEYINPUT57), .ZN(new_n1007));
  AND3_X1   g821(.A1(new_n977), .A2(new_n984), .A3(new_n985), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n985), .B1(new_n977), .B2(new_n984), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1007), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(new_n796), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n996), .A2(new_n771), .ZN(new_n1012));
  OR2_X1    g826(.A1(new_n1012), .A2(new_n854), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1005), .B1(new_n1011), .B2(new_n1013), .ZN(G54));
  NAND2_X1  g828(.A1(KEYINPUT58), .A2(G475), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n530), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1005), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NOR3_X1   g832(.A1(new_n1012), .A2(new_n530), .A3(new_n1015), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n1018), .A2(new_n1019), .ZN(G60));
  NAND2_X1  g834(.A1(G478), .A2(G902), .ZN(new_n1021));
  XOR2_X1   g835(.A(new_n1021), .B(KEYINPUT59), .Z(new_n1022));
  INV_X1    g836(.A(new_n1022), .ZN(new_n1023));
  AOI22_X1  g837(.A1(new_n987), .A2(new_n1023), .B1(new_n667), .B2(new_n668), .ZN(new_n1024));
  AND3_X1   g838(.A1(new_n667), .A2(new_n668), .A3(new_n1023), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1025), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1026), .A2(new_n1017), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n1024), .A2(new_n1027), .ZN(G63));
  INV_X1    g842(.A(KEYINPUT124), .ZN(new_n1029));
  AND4_X1   g843(.A1(new_n953), .A2(new_n983), .A3(new_n982), .A4(new_n959), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n943), .A2(new_n941), .ZN(new_n1031));
  NAND4_X1  g845(.A1(new_n1031), .A2(new_n953), .A3(new_n959), .A4(new_n965), .ZN(new_n1032));
  AOI22_X1  g846(.A1(new_n1030), .A2(new_n979), .B1(new_n1032), .B2(new_n973), .ZN(new_n1033));
  NAND2_X1  g847(.A1(G217), .A2(G902), .ZN(new_n1034));
  XNOR2_X1  g848(.A(new_n1034), .B(KEYINPUT60), .ZN(new_n1035));
  OAI211_X1 g849(.A(new_n1029), .B(new_n268), .C1(new_n1033), .C2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n1035), .B1(new_n977), .B2(new_n984), .ZN(new_n1037));
  OAI21_X1  g851(.A(KEYINPUT124), .B1(new_n1037), .B2(new_n269), .ZN(new_n1038));
  INV_X1    g852(.A(new_n707), .ZN(new_n1039));
  INV_X1    g853(.A(new_n709), .ZN(new_n1040));
  NOR2_X1   g854(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g855(.A(new_n1041), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n1005), .B1(new_n1037), .B2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g857(.A1(new_n1036), .A2(new_n1038), .A3(new_n1043), .A4(KEYINPUT61), .ZN(new_n1044));
  INV_X1    g858(.A(KEYINPUT61), .ZN(new_n1045));
  INV_X1    g859(.A(new_n1035), .ZN(new_n1046));
  NAND4_X1  g860(.A1(new_n983), .A2(new_n982), .A3(new_n953), .A4(new_n959), .ZN(new_n1047));
  INV_X1    g861(.A(new_n979), .ZN(new_n1048));
  NOR2_X1   g862(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  OAI211_X1 g863(.A(new_n1042), .B(new_n1046), .C1(new_n1049), .C2(new_n961), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n1050), .A2(new_n1017), .ZN(new_n1051));
  NOR2_X1   g865(.A1(new_n1037), .A2(new_n269), .ZN(new_n1052));
  OAI21_X1  g866(.A(new_n1045), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n1044), .A2(new_n1053), .ZN(G66));
  OAI21_X1  g868(.A(G953), .B1(new_n576), .B2(new_n607), .ZN(new_n1055));
  OAI21_X1  g869(.A(new_n1055), .B1(new_n1031), .B2(new_n245), .ZN(new_n1056));
  OAI21_X1  g870(.A(new_n999), .B1(G898), .B2(new_n244), .ZN(new_n1057));
  XNOR2_X1  g871(.A(new_n1056), .B(new_n1057), .ZN(G69));
  INV_X1    g872(.A(new_n389), .ZN(new_n1059));
  NAND3_X1  g873(.A1(new_n937), .A2(new_n938), .A3(new_n823), .ZN(new_n1060));
  NOR3_X1   g874(.A1(new_n1059), .A2(new_n757), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g875(.A(new_n1061), .B1(new_n874), .B2(new_n877), .ZN(new_n1062));
  INV_X1    g876(.A(KEYINPUT62), .ZN(new_n1063));
  AND3_X1   g877(.A1(new_n755), .A2(new_n758), .A3(new_n759), .ZN(new_n1064));
  NAND2_X1  g878(.A1(new_n957), .A2(new_n821), .ZN(new_n1065));
  OAI21_X1  g879(.A(new_n1063), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND4_X1  g880(.A1(new_n760), .A2(KEYINPUT62), .A3(new_n821), .A4(new_n957), .ZN(new_n1067));
  NAND2_X1  g881(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g882(.A1(new_n1062), .A2(new_n1068), .A3(new_n868), .ZN(new_n1069));
  NAND2_X1  g883(.A1(new_n1069), .A2(new_n244), .ZN(new_n1070));
  NAND2_X1  g884(.A1(new_n353), .A2(new_n355), .ZN(new_n1071));
  XOR2_X1   g885(.A(new_n1071), .B(new_n526), .Z(new_n1072));
  INV_X1    g886(.A(new_n1072), .ZN(new_n1073));
  AND4_X1   g887(.A1(new_n737), .A2(new_n764), .A3(new_n840), .A4(new_n821), .ZN(new_n1074));
  AND2_X1   g888(.A1(new_n835), .A2(new_n946), .ZN(new_n1075));
  NAND4_X1  g889(.A1(new_n864), .A2(new_n1075), .A3(new_n479), .A4(new_n756), .ZN(new_n1076));
  AND3_X1   g890(.A1(new_n1074), .A2(new_n838), .A3(new_n1076), .ZN(new_n1077));
  NAND4_X1  g891(.A1(new_n868), .A2(new_n878), .A3(new_n244), .A4(new_n1077), .ZN(new_n1078));
  AOI21_X1  g892(.A(new_n1073), .B1(G900), .B2(new_n245), .ZN(new_n1079));
  AOI22_X1  g893(.A1(new_n1070), .A2(new_n1073), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g894(.A(new_n244), .B1(G227), .B2(G900), .ZN(new_n1081));
  INV_X1    g895(.A(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g896(.A(new_n1080), .B(new_n1082), .ZN(G72));
  NAND2_X1  g897(.A1(G472), .A2(G902), .ZN(new_n1084));
  XOR2_X1   g898(.A(new_n1084), .B(KEYINPUT63), .Z(new_n1085));
  NOR2_X1   g899(.A1(new_n356), .A2(new_n357), .ZN(new_n1086));
  AOI21_X1  g900(.A(new_n1086), .B1(new_n385), .B2(KEYINPUT127), .ZN(new_n1087));
  OAI21_X1  g901(.A(new_n1087), .B1(KEYINPUT127), .B2(new_n385), .ZN(new_n1088));
  OAI211_X1 g902(.A(new_n1085), .B(new_n1088), .C1(new_n961), .C2(new_n975), .ZN(new_n1089));
  INV_X1    g903(.A(new_n740), .ZN(new_n1090));
  NAND4_X1  g904(.A1(new_n1062), .A2(new_n1068), .A3(new_n868), .A4(new_n1031), .ZN(new_n1091));
  AOI21_X1  g905(.A(new_n1090), .B1(new_n1091), .B2(new_n1085), .ZN(new_n1092));
  INV_X1    g906(.A(KEYINPUT125), .ZN(new_n1093));
  OAI211_X1 g907(.A(new_n1089), .B(new_n1017), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g908(.A1(new_n868), .A2(new_n878), .A3(new_n1031), .A4(new_n1077), .ZN(new_n1095));
  INV_X1    g909(.A(KEYINPUT126), .ZN(new_n1096));
  AND3_X1   g910(.A1(new_n1095), .A2(new_n1096), .A3(new_n1085), .ZN(new_n1097));
  AOI21_X1  g911(.A(new_n1096), .B1(new_n1095), .B2(new_n1085), .ZN(new_n1098));
  NAND2_X1  g912(.A1(new_n739), .A2(new_n347), .ZN(new_n1099));
  NOR3_X1   g913(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  AND2_X1   g914(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1101));
  NOR3_X1   g915(.A1(new_n1094), .A2(new_n1100), .A3(new_n1101), .ZN(G57));
endmodule


