//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 0 1 1 1 0 0 0 0 0 0 1 1 0 0 0 1 0 1 0 1 0 0 0 1 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n743,
    new_n744, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n804, new_n806, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n877,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n978, new_n979, new_n980, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1010, new_n1011, new_n1012;
  INV_X1    g000(.A(G22gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G15gat), .ZN(new_n203));
  INV_X1    g002(.A(G15gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G22gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G1gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT88), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(KEYINPUT16), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n203), .A2(new_n205), .A3(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n208), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  AND2_X1   g011(.A1(new_n203), .A2(new_n205), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n213), .A2(KEYINPUT88), .A3(new_n210), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(G8gat), .A3(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT89), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n213), .A2(new_n216), .A3(new_n210), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n211), .A2(KEYINPUT89), .ZN(new_n218));
  AOI21_X1  g017(.A(G8gat), .B1(new_n206), .B2(new_n207), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  AND3_X1   g019(.A1(new_n215), .A2(KEYINPUT90), .A3(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(KEYINPUT90), .B1(new_n215), .B2(new_n220), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT14), .ZN(new_n223));
  INV_X1    g022(.A(G29gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G36gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NOR3_X1   g028(.A1(new_n223), .A2(new_n228), .A3(G29gat), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT15), .ZN(new_n232));
  INV_X1    g031(.A(G43gat), .ZN(new_n233));
  INV_X1    g032(.A(G50gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(G43gat), .A2(G50gat), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n232), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n229), .A2(new_n231), .A3(new_n237), .ZN(new_n238));
  AND2_X1   g037(.A1(G43gat), .A2(G50gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(G43gat), .A2(G50gat), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT15), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n235), .A2(new_n232), .A3(new_n236), .ZN(new_n242));
  AOI21_X1  g041(.A(G36gat), .B1(new_n225), .B2(new_n226), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n241), .B(new_n242), .C1(new_n243), .C2(new_n230), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT87), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n238), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n247));
  AND2_X1   g046(.A1(new_n241), .A2(new_n242), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT87), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  NOR3_X1   g049(.A1(new_n221), .A2(new_n222), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n215), .A2(new_n220), .ZN(new_n252));
  OAI21_X1  g051(.A(KEYINPUT17), .B1(new_n246), .B2(new_n249), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n247), .A2(new_n248), .A3(KEYINPUT87), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n244), .A2(new_n245), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT17), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n254), .A2(new_n255), .A3(new_n256), .A4(new_n238), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n252), .B1(new_n253), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(G229gat), .A2(G233gat), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NOR3_X1   g059(.A1(new_n251), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(KEYINPUT91), .B1(new_n261), .B2(KEYINPUT18), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(KEYINPUT18), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(new_n259), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT90), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n215), .A2(KEYINPUT90), .A3(new_n220), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n254), .A2(new_n255), .A3(new_n238), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n270), .B1(new_n268), .B2(new_n269), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT93), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AOI211_X1 g073(.A(KEYINPUT93), .B(new_n270), .C1(new_n268), .C2(new_n269), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n266), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n253), .A2(new_n257), .ZN(new_n277));
  INV_X1    g076(.A(new_n252), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n279), .A2(new_n259), .A3(new_n271), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT91), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT18), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n262), .A2(new_n263), .A3(new_n276), .A4(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(G113gat), .B(G141gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G169gat), .B(G197gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(new_n289), .B(KEYINPUT12), .Z(new_n290));
  XNOR2_X1  g089(.A(new_n290), .B(KEYINPUT86), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n284), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT94), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n276), .A2(new_n263), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n290), .B1(new_n282), .B2(new_n280), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AND3_X1   g095(.A1(new_n292), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n293), .B1(new_n292), .B2(new_n296), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G8gat), .B(G36gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(G64gat), .B(G92gat), .ZN(new_n301));
  XOR2_X1   g100(.A(new_n300), .B(new_n301), .Z(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G211gat), .B(G218gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT65), .B(G211gat), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT22), .B1(new_n306), .B2(G218gat), .ZN(new_n307));
  XOR2_X1   g106(.A(G197gat), .B(G204gat), .Z(new_n308));
  OAI21_X1  g107(.A(new_n305), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AND2_X1   g108(.A1(KEYINPUT65), .A2(G211gat), .ZN(new_n310));
  NOR2_X1   g109(.A1(KEYINPUT65), .A2(G211gat), .ZN(new_n311));
  OAI21_X1  g110(.A(G218gat), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT22), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n308), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n314), .A2(new_n315), .A3(new_n304), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n309), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G226gat), .ZN(new_n318));
  INV_X1    g117(.A(G233gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AND2_X1   g119(.A1(G183gat), .A2(G190gat), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT24), .ZN(new_n322));
  AOI22_X1  g121(.A1(new_n321), .A2(new_n322), .B1(G169gat), .B2(G176gat), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT23), .ZN(new_n324));
  INV_X1    g123(.A(G169gat), .ZN(new_n325));
  INV_X1    g124(.A(G176gat), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(G183gat), .ZN(new_n330));
  INV_X1    g129(.A(G190gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(G183gat), .A2(G190gat), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(KEYINPUT24), .A3(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n323), .A2(new_n329), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT25), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n323), .A2(new_n329), .A3(new_n334), .A4(KEYINPUT25), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n330), .A2(KEYINPUT27), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT27), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(G183gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n340), .A2(new_n342), .A3(new_n331), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT28), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(KEYINPUT27), .B(G183gat), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n346), .A2(KEYINPUT28), .A3(new_n331), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n325), .A2(new_n326), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT26), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n333), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n351), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT29), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n320), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI22_X1  g156(.A1(new_n337), .A2(new_n338), .B1(new_n348), .B2(new_n353), .ZN(new_n358));
  INV_X1    g157(.A(new_n320), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n317), .B1(new_n357), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT66), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n359), .B1(new_n358), .B2(KEYINPUT29), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n355), .A2(new_n320), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n366), .A2(KEYINPUT66), .A3(new_n317), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT67), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n364), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n369), .B1(new_n364), .B2(new_n365), .ZN(new_n372));
  NOR3_X1   g171(.A1(new_n371), .A2(new_n372), .A3(new_n317), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n303), .B1(new_n368), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n366), .A2(KEYINPUT67), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n309), .A2(new_n316), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(new_n370), .A3(new_n376), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n377), .A2(new_n367), .A3(new_n363), .A4(new_n302), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n374), .A2(KEYINPUT30), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n368), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT30), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n380), .A2(new_n381), .A3(new_n377), .A4(new_n302), .ZN(new_n382));
  INV_X1    g181(.A(G141gat), .ZN(new_n383));
  INV_X1    g182(.A(G148gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G141gat), .A2(G148gat), .ZN(new_n386));
  AND2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(G155gat), .ZN(new_n388));
  INV_X1    g187(.A(G162gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(G155gat), .A2(G162gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n388), .A2(KEYINPUT69), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT69), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(G155gat), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n389), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT2), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n387), .B(new_n392), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n391), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n385), .B(new_n386), .C1(new_n399), .C2(new_n397), .ZN(new_n400));
  NOR2_X1   g199(.A1(G155gat), .A2(G162gat), .ZN(new_n401));
  NOR3_X1   g200(.A1(new_n399), .A2(new_n401), .A3(KEYINPUT68), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT68), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n403), .B1(new_n390), .B2(new_n391), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n400), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n398), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT71), .ZN(new_n407));
  XOR2_X1   g206(.A(G127gat), .B(G134gat), .Z(new_n408));
  XNOR2_X1  g207(.A(G113gat), .B(G120gat), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n408), .B1(KEYINPUT1), .B2(new_n409), .ZN(new_n410));
  XOR2_X1   g209(.A(G113gat), .B(G120gat), .Z(new_n411));
  INV_X1    g210(.A(KEYINPUT1), .ZN(new_n412));
  XNOR2_X1  g211(.A(G127gat), .B(G134gat), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT71), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n398), .A2(new_n405), .A3(new_n417), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n407), .A2(KEYINPUT4), .A3(new_n416), .A4(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n406), .A2(KEYINPUT3), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT3), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n398), .A2(new_n405), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n410), .A2(new_n414), .A3(KEYINPUT70), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT70), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n415), .A2(new_n424), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n420), .A2(new_n422), .A3(new_n423), .A4(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(G225gat), .A2(G233gat), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT4), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n428), .B1(new_n406), .B2(new_n415), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n419), .A2(new_n426), .A3(new_n427), .A4(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT5), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n425), .A2(new_n406), .A3(new_n423), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n416), .A2(new_n405), .A3(new_n398), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n427), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n431), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n426), .A2(new_n431), .A3(new_n427), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n407), .A2(new_n428), .A3(new_n416), .A4(new_n418), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n433), .A2(KEYINPUT4), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AOI22_X1  g239(.A1(new_n430), .A2(new_n436), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  XOR2_X1   g240(.A(G1gat), .B(G29gat), .Z(new_n442));
  XNOR2_X1  g241(.A(KEYINPUT72), .B(KEYINPUT0), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n442), .B(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(G57gat), .B(G85gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n444), .B(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT6), .B1(new_n441), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n436), .A2(new_n430), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n440), .A2(new_n431), .A3(new_n427), .A4(new_n426), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n446), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n447), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n450), .A2(KEYINPUT6), .A3(new_n451), .ZN(new_n454));
  AOI22_X1  g253(.A1(new_n379), .A2(new_n382), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(G227gat), .A2(G233gat), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n339), .A2(new_n416), .A3(new_n354), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n358), .A2(new_n416), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n457), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT33), .ZN(new_n462));
  XOR2_X1   g261(.A(G71gat), .B(G99gat), .Z(new_n463));
  XNOR2_X1  g262(.A(G15gat), .B(G43gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n463), .B(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT64), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n467), .B1(new_n466), .B2(new_n465), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n461), .A2(KEYINPUT32), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n355), .A2(new_n415), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n456), .B1(new_n470), .B2(new_n458), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT32), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n465), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n471), .A2(KEYINPUT33), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n469), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n470), .A2(new_n456), .A3(new_n458), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n476), .B(KEYINPUT34), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n461), .A2(KEYINPUT32), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n461), .A2(new_n462), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n479), .A2(new_n480), .A3(new_n465), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT34), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n476), .B(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n481), .A2(new_n483), .A3(new_n469), .ZN(new_n484));
  AND2_X1   g283(.A1(new_n478), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G78gat), .B(G106gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(KEYINPUT31), .B(G50gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(G228gat), .A2(G233gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n422), .A2(new_n356), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n489), .B1(new_n490), .B2(new_n317), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT74), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT29), .B1(new_n309), .B2(new_n316), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n406), .B1(new_n493), .B2(KEYINPUT3), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n491), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n492), .B1(new_n491), .B2(new_n494), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n376), .B1(new_n356), .B2(new_n422), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n309), .A2(KEYINPUT73), .A3(new_n316), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n356), .B1(new_n309), .B2(KEYINPUT73), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n421), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n407), .A2(new_n418), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n497), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n489), .ZN(new_n503));
  OAI22_X1  g302(.A1(new_n495), .A2(new_n496), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n488), .B1(new_n504), .B2(G22gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n317), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n304), .B1(new_n314), .B2(new_n315), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT73), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT29), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n309), .A2(KEYINPUT73), .A3(new_n316), .ZN(new_n510));
  AOI21_X1  g309(.A(KEYINPUT3), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n398), .A2(new_n405), .A3(new_n417), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n417), .B1(new_n398), .B2(new_n405), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n506), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n489), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n516), .B(new_n202), .C1(new_n496), .C2(new_n495), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT75), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n491), .A2(new_n494), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT74), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n491), .A2(new_n492), .A3(new_n494), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT75), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n522), .A2(new_n523), .A3(new_n202), .A4(new_n516), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n505), .A2(new_n518), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT77), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n517), .A2(KEYINPUT76), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n202), .B1(new_n522), .B2(new_n516), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT76), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n504), .A2(new_n530), .A3(G22gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(new_n488), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n525), .B(new_n526), .C1(new_n529), .C2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n504), .A2(G22gat), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n535), .A2(KEYINPUT76), .A3(new_n517), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n536), .A2(new_n488), .A3(new_n531), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n526), .B1(new_n537), .B2(new_n525), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n455), .B(new_n485), .C1(new_n534), .C2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT35), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT84), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n534), .A2(new_n538), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT35), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n478), .A2(new_n484), .A3(new_n543), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n451), .B1(new_n441), .B2(KEYINPUT82), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT82), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n450), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n447), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n544), .B1(new_n548), .B2(new_n454), .ZN(new_n549));
  AND3_X1   g348(.A1(new_n379), .A2(KEYINPUT78), .A3(new_n382), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT78), .B1(new_n379), .B2(new_n382), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n541), .B1(new_n542), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n448), .A2(new_n449), .A3(new_n446), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT6), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n446), .B1(new_n450), .B2(new_n546), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n441), .A2(KEYINPUT82), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n454), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n485), .B(new_n543), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n379), .A2(KEYINPUT78), .A3(new_n382), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n379), .A2(new_n382), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT78), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n561), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n525), .B1(new_n529), .B2(new_n532), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT77), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(new_n533), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n566), .A2(KEYINPUT84), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n540), .A2(new_n553), .A3(new_n570), .ZN(new_n571));
  OR3_X1    g370(.A1(new_n534), .A2(new_n538), .A3(new_n455), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n485), .B(KEYINPUT36), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n548), .A2(new_n454), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n364), .A2(new_n365), .A3(new_n376), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(KEYINPUT83), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n376), .B1(new_n375), .B2(new_n370), .ZN(new_n577));
  OAI21_X1  g376(.A(KEYINPUT37), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT38), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n377), .A2(new_n367), .A3(new_n363), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n303), .B1(new_n581), .B2(KEYINPUT37), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT37), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n584), .B1(new_n380), .B2(new_n377), .ZN(new_n585));
  OAI21_X1  g384(.A(KEYINPUT38), .B1(new_n585), .B2(new_n582), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n583), .A2(new_n586), .A3(new_n378), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n569), .B1(new_n574), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n427), .B1(new_n440), .B2(new_n426), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT39), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(new_n446), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n432), .A2(new_n433), .A3(new_n427), .ZN(new_n593));
  AND3_X1   g392(.A1(new_n593), .A2(KEYINPUT79), .A3(KEYINPUT39), .ZN(new_n594));
  AOI21_X1  g393(.A(KEYINPUT79), .B1(new_n593), .B2(KEYINPUT39), .ZN(new_n595));
  NOR3_X1   g394(.A1(new_n589), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT80), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT81), .ZN(new_n598));
  OAI22_X1  g397(.A1(new_n592), .A2(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT40), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n557), .A2(new_n558), .ZN(new_n601));
  OAI22_X1  g400(.A1(new_n592), .A2(new_n596), .B1(new_n597), .B2(KEYINPUT40), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(new_n598), .ZN(new_n603));
  NOR3_X1   g402(.A1(new_n592), .A2(new_n596), .A3(new_n597), .ZN(new_n604));
  OAI211_X1 g403(.A(new_n600), .B(new_n601), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  NOR3_X1   g404(.A1(new_n605), .A2(new_n550), .A3(new_n551), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n572), .B(new_n573), .C1(new_n588), .C2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n299), .B1(new_n571), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT108), .ZN(new_n609));
  NAND2_X1  g408(.A1(G71gat), .A2(G78gat), .ZN(new_n610));
  INV_X1    g409(.A(G71gat), .ZN(new_n611));
  INV_X1    g410(.A(G78gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G57gat), .B(G64gat), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT95), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT9), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n610), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n618), .B1(new_n614), .B2(new_n615), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n610), .B(new_n613), .C1(new_n616), .C2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(G57gat), .ZN(new_n621));
  OR2_X1    g420(.A1(KEYINPUT96), .A2(G64gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(KEYINPUT96), .A2(G64gat), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT97), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n610), .B1(new_n613), .B2(new_n617), .ZN(new_n627));
  INV_X1    g426(.A(G64gat), .ZN(new_n628));
  OAI21_X1  g427(.A(KEYINPUT97), .B1(new_n628), .B2(G57gat), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n626), .B(new_n627), .C1(new_n624), .C2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n620), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT21), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(G231gat), .A2(G233gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G127gat), .B(G155gat), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n636), .B(KEYINPUT20), .Z(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n635), .B(new_n638), .ZN(new_n639));
  OAI22_X1  g438(.A1(new_n221), .A2(new_n222), .B1(new_n632), .B2(new_n631), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT99), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n635), .B(new_n637), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(new_n641), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G183gat), .B(G211gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(KEYINPUT98), .B(KEYINPUT19), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G134gat), .B(G162gat), .ZN(new_n652));
  AOI21_X1  g451(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G99gat), .B(G106gat), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT100), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT7), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n660), .A2(G85gat), .A3(G92gat), .A4(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(G99gat), .A2(G106gat), .ZN(new_n664));
  INV_X1    g463(.A(G85gat), .ZN(new_n665));
  INV_X1    g464(.A(G92gat), .ZN(new_n666));
  AOI22_X1  g465(.A1(KEYINPUT8), .A2(new_n664), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OAI211_X1 g466(.A(new_n658), .B(new_n659), .C1(new_n665), .C2(new_n666), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n657), .B1(new_n663), .B2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT101), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n662), .A2(new_n656), .A3(new_n668), .A4(new_n667), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  OAI211_X1 g472(.A(KEYINPUT101), .B(new_n657), .C1(new_n663), .C2(new_n669), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(KEYINPUT102), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT102), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n673), .A2(new_n677), .A3(new_n674), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(new_n277), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n676), .A2(new_n270), .A3(new_n678), .ZN(new_n681));
  NAND3_X1  g480(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(G190gat), .B(G218gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT103), .B(KEYINPUT104), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n684), .B(new_n685), .Z(new_n686));
  NAND2_X1  g485(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n683), .A2(new_n686), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n655), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  OR2_X1    g489(.A1(new_n683), .A2(new_n686), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n691), .A2(new_n654), .A3(new_n687), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n643), .A2(new_n645), .A3(new_n649), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n651), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT10), .ZN(new_n696));
  AOI22_X1  g495(.A1(new_n673), .A2(new_n674), .B1(new_n620), .B2(new_n630), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n670), .A2(new_n672), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n698), .A2(new_n620), .A3(new_n630), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n696), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n631), .A2(new_n696), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n676), .A2(new_n678), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(G230gat), .A2(G233gat), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n697), .A2(new_n699), .A3(new_n704), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(G120gat), .B(G148gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT106), .ZN(new_n710));
  XNOR2_X1  g509(.A(G176gat), .B(G204gat), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n712), .B1(new_n706), .B2(new_n707), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n705), .A2(new_n708), .A3(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n704), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n716), .B1(new_n700), .B2(new_n702), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n712), .B1(new_n717), .B2(new_n706), .ZN(new_n718));
  OR2_X1    g517(.A1(new_n718), .A2(KEYINPUT107), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(KEYINPUT107), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n715), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n609), .B1(new_n695), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n695), .A2(new_n722), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(KEYINPUT108), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n608), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n453), .A2(new_n454), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(new_n207), .ZN(G1324gat));
  NOR2_X1   g528(.A1(new_n550), .A2(new_n551), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n726), .A2(new_n731), .ZN(new_n732));
  XOR2_X1   g531(.A(KEYINPUT16), .B(G8gat), .Z(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT42), .ZN(new_n735));
  OAI21_X1  g534(.A(G8gat), .B1(new_n726), .B2(new_n731), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT109), .ZN(new_n737));
  OR2_X1    g536(.A1(new_n736), .A2(KEYINPUT109), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n735), .A2(new_n737), .A3(new_n738), .ZN(G1325gat));
  OAI21_X1  g538(.A(G15gat), .B1(new_n726), .B2(new_n573), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n485), .A2(new_n204), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n726), .B2(new_n741), .ZN(G1326gat));
  NOR2_X1   g541(.A1(new_n726), .A2(new_n569), .ZN(new_n743));
  XOR2_X1   g542(.A(KEYINPUT43), .B(G22gat), .Z(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(G1327gat));
  NAND2_X1  g544(.A1(new_n651), .A2(new_n694), .ZN(new_n746));
  INV_X1    g545(.A(new_n693), .ZN(new_n747));
  AND4_X1   g546(.A1(new_n608), .A2(new_n746), .A3(new_n747), .A4(new_n721), .ZN(new_n748));
  INV_X1    g547(.A(new_n727), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n748), .A2(new_n224), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT45), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n571), .A2(new_n607), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(new_n747), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT44), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n693), .B1(new_n571), .B2(new_n607), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT44), .ZN(new_n757));
  INV_X1    g556(.A(new_n746), .ZN(new_n758));
  AOI22_X1  g557(.A1(new_n284), .A2(new_n291), .B1(new_n294), .B2(new_n295), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n758), .A2(new_n759), .A3(new_n722), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n755), .A2(new_n757), .A3(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT110), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n755), .A2(KEYINPUT110), .A3(new_n757), .A4(new_n760), .ZN(new_n764));
  AND3_X1   g563(.A1(new_n763), .A2(new_n749), .A3(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n751), .B1(new_n765), .B2(new_n224), .ZN(G1328gat));
  NAND3_X1  g565(.A1(new_n748), .A2(new_n228), .A3(new_n730), .ZN(new_n767));
  XOR2_X1   g566(.A(new_n767), .B(KEYINPUT46), .Z(new_n768));
  AND3_X1   g567(.A1(new_n763), .A2(new_n730), .A3(new_n764), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n228), .B2(new_n769), .ZN(G1329gat));
  OAI21_X1  g569(.A(G43gat), .B1(new_n761), .B2(new_n573), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n748), .A2(new_n233), .A3(new_n485), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n771), .A2(KEYINPUT47), .A3(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n772), .ZN(new_n774));
  INV_X1    g573(.A(new_n573), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n763), .A2(new_n775), .A3(new_n764), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n774), .B1(new_n776), .B2(G43gat), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n773), .B1(new_n777), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g577(.A(G50gat), .B1(new_n761), .B2(new_n569), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n569), .A2(G50gat), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT111), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n748), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n779), .A2(KEYINPUT48), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n782), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n763), .A2(new_n542), .A3(new_n764), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n784), .B1(new_n785), .B2(G50gat), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n783), .B1(new_n786), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g586(.A1(new_n292), .A2(new_n296), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n695), .A2(new_n788), .A3(new_n721), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n752), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n790), .A2(new_n727), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(new_n621), .ZN(G1332gat));
  NAND2_X1  g591(.A1(new_n730), .A2(KEYINPUT112), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT112), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n794), .B1(new_n550), .B2(new_n551), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n790), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n798));
  AND2_X1   g597(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n800), .B1(new_n797), .B2(new_n798), .ZN(G1333gat));
  OAI21_X1  g600(.A(G71gat), .B1(new_n790), .B2(new_n573), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n485), .A2(new_n611), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n802), .B1(new_n790), .B2(new_n803), .ZN(new_n804));
  XOR2_X1   g603(.A(new_n804), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g604(.A1(new_n790), .A2(new_n569), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(new_n612), .ZN(G1335gat));
  NOR2_X1   g606(.A1(new_n758), .A2(new_n788), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n722), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(KEYINPUT113), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n755), .A2(new_n757), .A3(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(G85gat), .B1(new_n812), .B2(new_n727), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n756), .A2(new_n808), .ZN(new_n814));
  OR2_X1    g613(.A1(new_n814), .A2(KEYINPUT51), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(KEYINPUT51), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n815), .A2(new_n722), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n749), .A2(new_n665), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n813), .B1(new_n817), .B2(new_n818), .ZN(G1336gat));
  INV_X1    g618(.A(new_n812), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n730), .ZN(new_n821));
  NOR2_X1   g620(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n814), .B(new_n822), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n796), .A2(G92gat), .A3(new_n721), .ZN(new_n824));
  AOI22_X1  g623(.A1(new_n821), .A2(G92gat), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n826));
  INV_X1    g625(.A(new_n796), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n666), .B1(new_n820), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n815), .A2(new_n816), .A3(new_n824), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n826), .ZN(new_n830));
  OAI22_X1  g629(.A1(new_n825), .A2(new_n826), .B1(new_n828), .B2(new_n830), .ZN(G1337gat));
  OAI21_X1  g630(.A(G99gat), .B1(new_n812), .B2(new_n573), .ZN(new_n832));
  INV_X1    g631(.A(G99gat), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n485), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n832), .B1(new_n817), .B2(new_n834), .ZN(G1338gat));
  NAND2_X1  g634(.A1(new_n820), .A2(new_n542), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n569), .A2(G106gat), .A3(new_n721), .ZN(new_n837));
  AOI22_X1  g636(.A1(new_n836), .A2(G106gat), .B1(new_n823), .B2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT53), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n836), .A2(G106gat), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n815), .A2(new_n816), .A3(new_n837), .ZN(new_n841));
  XOR2_X1   g640(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI22_X1  g642(.A1(new_n838), .A2(new_n839), .B1(new_n840), .B2(new_n843), .ZN(G1339gat));
  NAND2_X1  g643(.A1(new_n724), .A2(new_n759), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n274), .A2(new_n275), .A3(new_n266), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n259), .B1(new_n279), .B2(new_n271), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n289), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n690), .A2(new_n296), .A3(new_n692), .A4(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n700), .A2(new_n702), .A3(new_n716), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n705), .A2(new_n850), .A3(KEYINPUT54), .ZN(new_n851));
  INV_X1    g650(.A(new_n712), .ZN(new_n852));
  XNOR2_X1  g651(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n852), .B1(new_n717), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT55), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n717), .A2(new_n853), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n851), .A2(KEYINPUT55), .A3(new_n712), .A4(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n857), .A2(new_n714), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n849), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n296), .A2(new_n848), .ZN(new_n862));
  OAI22_X1  g661(.A1(new_n860), .A2(new_n759), .B1(new_n721), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n861), .B1(new_n863), .B2(new_n693), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n845), .B1(new_n864), .B2(new_n758), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n569), .A2(new_n485), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n827), .A2(new_n727), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(G113gat), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n869), .A2(new_n870), .A3(new_n299), .ZN(new_n871));
  INV_X1    g670(.A(new_n869), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n788), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n871), .B1(new_n870), .B2(new_n873), .ZN(G1340gat));
  NAND2_X1  g673(.A1(new_n872), .A2(new_n722), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g675(.A1(new_n872), .A2(new_n758), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(G127gat), .ZN(G1342gat));
  OAI21_X1  g677(.A(G134gat), .B1(new_n869), .B2(new_n693), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n730), .A2(new_n693), .ZN(new_n880));
  INV_X1    g679(.A(G134gat), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n880), .A2(new_n881), .A3(new_n749), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n867), .A2(KEYINPUT56), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(KEYINPUT56), .B1(new_n867), .B2(new_n883), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n879), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  XOR2_X1   g685(.A(new_n886), .B(KEYINPUT117), .Z(G1343gat));
  NAND2_X1  g686(.A1(new_n865), .A2(new_n542), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n796), .A2(new_n749), .A3(new_n573), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n891), .A2(G141gat), .A3(new_n299), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT57), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n569), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n860), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n896), .B1(new_n297), .B2(new_n298), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n721), .A2(new_n862), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n747), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n746), .B1(new_n900), .B2(new_n861), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n895), .B1(new_n901), .B2(new_n845), .ZN(new_n902));
  XNOR2_X1  g701(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n903));
  AOI22_X1  g702(.A1(new_n902), .A2(KEYINPUT119), .B1(new_n888), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n788), .A2(KEYINPUT94), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n759), .A2(new_n293), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n860), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n693), .B1(new_n907), .B2(new_n898), .ZN(new_n908));
  INV_X1    g707(.A(new_n861), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n758), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(new_n845), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n894), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT119), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n889), .B1(new_n904), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(new_n788), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n892), .B1(new_n916), .B2(G141gat), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT58), .ZN(new_n918));
  INV_X1    g717(.A(new_n299), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n383), .B1(new_n915), .B2(new_n919), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n892), .A2(KEYINPUT58), .ZN(new_n921));
  OAI22_X1  g720(.A1(new_n917), .A2(new_n918), .B1(new_n920), .B2(new_n921), .ZN(G1344gat));
  INV_X1    g721(.A(new_n889), .ZN(new_n923));
  INV_X1    g722(.A(new_n888), .ZN(new_n924));
  INV_X1    g723(.A(new_n903), .ZN(new_n925));
  OAI22_X1  g724(.A1(new_n912), .A2(new_n913), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n902), .A2(KEYINPUT119), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n722), .B(new_n923), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n384), .A2(KEYINPUT59), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n865), .A2(new_n542), .A3(new_n925), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n725), .A2(new_n299), .A3(new_n723), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n542), .B1(new_n910), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n930), .B1(new_n932), .B2(new_n893), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n889), .A2(KEYINPUT120), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n889), .A2(KEYINPUT120), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n934), .A2(new_n722), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g735(.A(G148gat), .B1(new_n933), .B2(new_n936), .ZN(new_n937));
  AOI22_X1  g736(.A1(new_n928), .A2(new_n929), .B1(new_n937), .B2(KEYINPUT59), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n890), .A2(new_n384), .A3(new_n722), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(KEYINPUT121), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT121), .ZN(new_n942));
  INV_X1    g741(.A(new_n929), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n943), .B1(new_n915), .B2(new_n722), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT59), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n725), .A2(new_n299), .A3(new_n723), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n569), .B1(new_n901), .B2(new_n946), .ZN(new_n947));
  OAI22_X1  g746(.A1(new_n947), .A2(KEYINPUT57), .B1(new_n888), .B2(new_n903), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n948), .A2(new_n722), .A3(new_n934), .A4(new_n935), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n945), .B1(new_n949), .B2(G148gat), .ZN(new_n950));
  OAI211_X1 g749(.A(new_n942), .B(new_n939), .C1(new_n944), .C2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n941), .A2(new_n951), .ZN(G1345gat));
  NAND2_X1  g751(.A1(new_n393), .A2(new_n395), .ZN(new_n953));
  INV_X1    g752(.A(new_n915), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n953), .B1(new_n954), .B2(new_n746), .ZN(new_n955));
  OR2_X1    g754(.A1(new_n746), .A2(new_n953), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n955), .B1(new_n891), .B2(new_n956), .ZN(G1346gat));
  OAI21_X1  g756(.A(G162gat), .B1(new_n954), .B2(new_n693), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n880), .A2(new_n389), .A3(new_n749), .A4(new_n573), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n958), .B1(new_n888), .B2(new_n959), .ZN(G1347gat));
  NAND2_X1  g759(.A1(new_n730), .A2(new_n727), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT122), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n867), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g762(.A(G169gat), .B1(new_n963), .B2(new_n299), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n865), .A2(new_n727), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n827), .A2(new_n866), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n788), .A2(new_n325), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n964), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  XOR2_X1   g768(.A(new_n969), .B(KEYINPUT123), .Z(G1348gat));
  INV_X1    g769(.A(new_n967), .ZN(new_n971));
  AOI21_X1  g770(.A(G176gat), .B1(new_n971), .B2(new_n722), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n867), .A2(G176gat), .A3(new_n722), .A4(new_n962), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT124), .ZN(new_n974));
  AND2_X1   g773(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n973), .A2(new_n974), .ZN(new_n976));
  NOR3_X1   g775(.A1(new_n972), .A2(new_n975), .A3(new_n976), .ZN(G1349gat));
  OAI21_X1  g776(.A(G183gat), .B1(new_n963), .B2(new_n746), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n758), .A2(new_n346), .ZN(new_n979));
  OAI211_X1 g778(.A(new_n978), .B(KEYINPUT125), .C1(new_n967), .C2(new_n979), .ZN(new_n980));
  XNOR2_X1  g779(.A(new_n980), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g780(.A1(new_n971), .A2(new_n331), .A3(new_n747), .ZN(new_n982));
  OAI21_X1  g781(.A(G190gat), .B1(new_n963), .B2(new_n693), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n983), .A2(KEYINPUT61), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n983), .A2(KEYINPUT61), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n982), .B1(new_n984), .B2(new_n985), .ZN(G1351gat));
  AND4_X1   g785(.A1(new_n542), .A2(new_n965), .A3(new_n573), .A4(new_n827), .ZN(new_n987));
  AOI21_X1  g786(.A(G197gat), .B1(new_n987), .B2(new_n788), .ZN(new_n988));
  AND2_X1   g787(.A1(new_n962), .A2(new_n573), .ZN(new_n989));
  AND2_X1   g788(.A1(new_n948), .A2(new_n989), .ZN(new_n990));
  AND2_X1   g789(.A1(new_n919), .A2(G197gat), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n988), .B1(new_n990), .B2(new_n991), .ZN(G1352gat));
  AOI21_X1  g791(.A(G204gat), .B1(KEYINPUT126), .B2(KEYINPUT62), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n987), .A2(new_n722), .A3(new_n993), .ZN(new_n994));
  NOR2_X1   g793(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n995));
  XNOR2_X1  g794(.A(new_n994), .B(new_n995), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n990), .A2(new_n722), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n997), .A2(G204gat), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n996), .A2(new_n998), .ZN(G1353gat));
  NOR2_X1   g798(.A1(new_n746), .A2(new_n306), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n987), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g800(.A(KEYINPUT127), .ZN(new_n1002));
  NAND4_X1  g801(.A1(new_n948), .A2(new_n1002), .A3(new_n758), .A4(new_n989), .ZN(new_n1003));
  AND2_X1   g802(.A1(new_n1003), .A2(G211gat), .ZN(new_n1004));
  NAND3_X1  g803(.A1(new_n948), .A2(new_n758), .A3(new_n989), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1005), .A2(KEYINPUT127), .ZN(new_n1006));
  AOI21_X1  g805(.A(KEYINPUT63), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  AND4_X1   g806(.A1(KEYINPUT63), .A2(new_n1006), .A3(G211gat), .A4(new_n1003), .ZN(new_n1008));
  OAI21_X1  g807(.A(new_n1001), .B1(new_n1007), .B2(new_n1008), .ZN(G1354gat));
  INV_X1    g808(.A(G218gat), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n987), .A2(new_n1010), .A3(new_n747), .ZN(new_n1011));
  AND2_X1   g810(.A1(new_n990), .A2(new_n747), .ZN(new_n1012));
  OAI21_X1  g811(.A(new_n1011), .B1(new_n1012), .B2(new_n1010), .ZN(G1355gat));
endmodule


