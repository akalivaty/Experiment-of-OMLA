//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 0 1 0 1 0 1 0 0 0 1 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 1 0 0 1 1 0 1 0 1 0 0 0 1 0 1 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n842,
    new_n843, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1023, new_n1024, new_n1025, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1062,
    new_n1063;
  INV_X1    g000(.A(KEYINPUT91), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT36), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT69), .ZN(new_n204));
  INV_X1    g003(.A(G113gat), .ZN(new_n205));
  INV_X1    g004(.A(G120gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT1), .ZN(new_n208));
  NAND2_X1  g007(.A1(G113gat), .A2(G120gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G134gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G127gat), .ZN(new_n212));
  INV_X1    g011(.A(G127gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G134gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n210), .A2(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT1), .B1(new_n205), .B2(new_n206), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n217), .A2(new_n209), .B1(new_n212), .B2(new_n214), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n204), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n210), .A2(new_n215), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n217), .A2(new_n209), .A3(new_n212), .A4(new_n214), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(new_n221), .A3(KEYINPUT69), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224));
  AND2_X1   g023(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n224), .B1(new_n225), .B2(G190gat), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n227), .A2(KEYINPUT65), .ZN(new_n228));
  NAND2_X1  g027(.A1(G183gat), .A2(G190gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT24), .ZN(new_n230));
  AND3_X1   g029(.A1(new_n229), .A2(KEYINPUT65), .A3(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n226), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NOR2_X1   g033(.A1(G169gat), .A2(G176gat), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G169gat), .A2(G176gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT23), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n235), .A2(KEYINPUT23), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n239), .A2(KEYINPUT25), .A3(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n242), .B1(G183gat), .B2(G190gat), .ZN(new_n243));
  OR2_X1    g042(.A1(new_n227), .A2(KEYINPUT65), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n227), .A2(KEYINPUT65), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n241), .B1(new_n246), .B2(KEYINPUT66), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT23), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n248), .B1(G169gat), .B2(G176gat), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n240), .B1(new_n249), .B2(new_n235), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT64), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  OAI211_X1 g051(.A(KEYINPUT64), .B(new_n240), .C1(new_n249), .C2(new_n235), .ZN(new_n253));
  INV_X1    g052(.A(new_n227), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n226), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n252), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT25), .ZN(new_n257));
  AOI22_X1  g056(.A1(new_n234), .A2(new_n247), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT28), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT67), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT27), .B(G183gat), .ZN(new_n261));
  INV_X1    g060(.A(G190gat), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(G183gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT27), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT27), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(G183gat), .ZN(new_n267));
  AND4_X1   g066(.A1(new_n260), .A2(new_n265), .A3(new_n267), .A4(new_n262), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n259), .B1(new_n263), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n265), .A2(new_n267), .A3(new_n262), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT67), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n261), .A2(new_n260), .A3(new_n262), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n271), .A2(new_n272), .A3(KEYINPUT28), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT26), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n236), .A2(new_n274), .A3(new_n237), .ZN(new_n275));
  AOI22_X1  g074(.A1(new_n235), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT68), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT68), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n275), .A2(new_n276), .A3(new_n279), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n269), .A2(new_n273), .A3(new_n278), .A4(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n223), .B1(new_n258), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G227gat), .ZN(new_n284));
  INV_X1    g083(.A(G233gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI211_X1 g085(.A(KEYINPUT66), .B(new_n226), .C1(new_n228), .C2(new_n231), .ZN(new_n287));
  INV_X1    g086(.A(new_n241), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n234), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n253), .A2(new_n255), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT64), .B1(new_n239), .B2(new_n240), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n257), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  NOR3_X1   g092(.A1(new_n216), .A2(new_n218), .A3(new_n204), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT69), .B1(new_n220), .B2(new_n221), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n293), .A2(new_n296), .A3(new_n281), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n283), .A2(new_n286), .A3(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT33), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  XOR2_X1   g099(.A(G15gat), .B(G43gat), .Z(new_n301));
  XNOR2_X1  g100(.A(G71gat), .B(G99gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n301), .B(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  AOI211_X1 g103(.A(KEYINPUT34), .B(new_n286), .C1(new_n283), .C2(new_n297), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n283), .A2(new_n297), .ZN(new_n307));
  INV_X1    g106(.A(new_n286), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT34), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n304), .A2(new_n306), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n298), .A2(KEYINPUT32), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n303), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n314), .B1(new_n298), .B2(new_n299), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT34), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n316), .B1(new_n307), .B2(new_n308), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n315), .B1(new_n317), .B2(new_n305), .ZN(new_n318));
  AND3_X1   g117(.A1(new_n311), .A2(new_n313), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n313), .B1(new_n311), .B2(new_n318), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n203), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n311), .A2(new_n318), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(new_n312), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n311), .A2(new_n313), .A3(new_n318), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n323), .A2(KEYINPUT36), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT72), .ZN(new_n327));
  NAND2_X1  g126(.A1(G211gat), .A2(G218gat), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT22), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(G197gat), .ZN(new_n331));
  INV_X1    g130(.A(G204gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G197gat), .A2(G204gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(G211gat), .ZN(new_n336));
  INV_X1    g135(.A(G218gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT70), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n338), .A2(new_n339), .A3(new_n328), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n339), .B1(new_n338), .B2(new_n328), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n330), .B(new_n335), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n335), .A2(new_n330), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n338), .A2(new_n328), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT70), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n346), .A3(new_n340), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(G226gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n349), .A2(new_n285), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT71), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n352), .B1(new_n258), .B2(new_n282), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n293), .A2(KEYINPUT71), .A3(new_n281), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n351), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n350), .A2(KEYINPUT29), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n357), .B1(new_n293), .B2(new_n281), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n327), .B(new_n348), .C1(new_n355), .C2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n348), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n293), .A2(new_n281), .A3(new_n350), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n353), .A2(new_n354), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n360), .B(new_n361), .C1(new_n362), .C2(new_n357), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT30), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n358), .B1(new_n362), .B2(new_n350), .ZN(new_n367));
  OAI21_X1  g166(.A(KEYINPUT72), .B1(new_n367), .B2(new_n360), .ZN(new_n368));
  XNOR2_X1  g167(.A(G8gat), .B(G36gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(G64gat), .B(G92gat), .ZN(new_n370));
  XOR2_X1   g169(.A(new_n369), .B(new_n370), .Z(new_n371));
  NAND4_X1  g170(.A1(new_n365), .A2(new_n366), .A3(new_n368), .A4(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n371), .ZN(new_n373));
  AND3_X1   g172(.A1(new_n293), .A2(KEYINPUT71), .A3(new_n281), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT71), .B1(new_n293), .B2(new_n281), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n350), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n358), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n327), .B1(new_n378), .B2(new_n348), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n373), .B1(new_n364), .B2(new_n379), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n368), .A2(new_n359), .A3(new_n363), .A4(new_n371), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(KEYINPUT30), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n220), .A2(new_n221), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n383), .B(KEYINPUT77), .ZN(new_n384));
  INV_X1    g183(.A(G155gat), .ZN(new_n385));
  INV_X1    g184(.A(G162gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(G155gat), .A2(G162gat), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(KEYINPUT75), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(KEYINPUT2), .ZN(new_n390));
  AND2_X1   g189(.A1(G141gat), .A2(G148gat), .ZN(new_n391));
  NOR2_X1   g190(.A1(G141gat), .A2(G148gat), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AND3_X1   g192(.A1(new_n389), .A2(new_n390), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT75), .ZN(new_n395));
  INV_X1    g194(.A(new_n388), .ZN(new_n396));
  NOR2_X1   g195(.A1(G155gat), .A2(G162gat), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OR2_X1    g197(.A1(G141gat), .A2(G148gat), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT73), .ZN(new_n400));
  NAND2_X1  g199(.A1(G141gat), .A2(G148gat), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT73), .B1(new_n391), .B2(new_n392), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT2), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT74), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT74), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT2), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n402), .A2(new_n403), .A3(new_n408), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n396), .A2(new_n397), .ZN(new_n410));
  AOI22_X1  g209(.A1(new_n394), .A2(new_n398), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT76), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n409), .A2(new_n410), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n398), .A2(new_n389), .A3(new_n390), .A4(new_n393), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT76), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n384), .A2(new_n413), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT79), .ZN(new_n419));
  AND3_X1   g218(.A1(new_n414), .A2(new_n412), .A3(new_n415), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n412), .B1(new_n414), .B2(new_n415), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT79), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n422), .A2(new_n423), .A3(new_n384), .ZN(new_n424));
  INV_X1    g223(.A(new_n383), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n411), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT80), .B(KEYINPUT5), .ZN(new_n427));
  NAND2_X1  g226(.A1(G225gat), .A2(G233gat), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n419), .A2(new_n424), .A3(new_n426), .A4(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT4), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n411), .A2(new_n431), .A3(new_n425), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n431), .B1(new_n223), .B2(new_n411), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT78), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI211_X1 g234(.A(KEYINPUT78), .B(new_n431), .C1(new_n223), .C2(new_n411), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n427), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT3), .ZN(new_n439));
  NOR3_X1   g238(.A1(new_n420), .A2(new_n421), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n411), .A2(new_n439), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n384), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n438), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n428), .B1(new_n437), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n223), .A2(new_n431), .A3(new_n411), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT82), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT82), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n223), .A2(new_n411), .A3(new_n447), .A4(new_n431), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n426), .A2(KEYINPUT4), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n446), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n384), .A2(new_n441), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n413), .A2(new_n417), .A3(KEYINPUT3), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n438), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n430), .B1(new_n444), .B2(new_n454), .ZN(new_n455));
  XOR2_X1   g254(.A(G1gat), .B(G29gat), .Z(new_n456));
  XNOR2_X1  g255(.A(G57gat), .B(G85gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n456), .B(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n459));
  XOR2_X1   g258(.A(new_n458), .B(new_n459), .Z(new_n460));
  NAND2_X1  g259(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT6), .ZN(new_n462));
  INV_X1    g261(.A(new_n460), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n463), .B(new_n430), .C1(new_n444), .C2(new_n454), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n461), .A2(KEYINPUT83), .A3(new_n462), .A4(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT83), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n455), .B(new_n460), .C1(new_n466), .C2(KEYINPUT6), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n372), .A2(new_n382), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT88), .ZN(new_n469));
  XNOR2_X1  g268(.A(G78gat), .B(G106gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(KEYINPUT31), .B(G50gat), .ZN(new_n471));
  XOR2_X1   g270(.A(new_n470), .B(new_n471), .Z(new_n472));
  NOR2_X1   g271(.A1(new_n472), .A2(KEYINPUT87), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT29), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n441), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n360), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n344), .A2(new_n346), .A3(KEYINPUT84), .A4(new_n340), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n477), .A2(new_n474), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT84), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n343), .A2(new_n347), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT3), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n476), .B1(new_n411), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(G228gat), .A2(G233gat), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT29), .B1(new_n343), .B2(new_n347), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n439), .B1(new_n484), .B2(KEYINPUT85), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n348), .A2(KEYINPUT85), .A3(new_n474), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n422), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n483), .B1(new_n475), .B2(new_n360), .ZN(new_n488));
  AOI22_X1  g287(.A1(new_n482), .A2(new_n483), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(G22gat), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n473), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n481), .A2(new_n411), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n348), .B1(new_n441), .B2(new_n474), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n483), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n487), .A2(new_n488), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n473), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(G22gat), .A3(new_n497), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n491), .A2(new_n498), .B1(new_n490), .B2(new_n489), .ZN(new_n499));
  INV_X1    g298(.A(new_n472), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT86), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n489), .A2(new_n501), .A3(new_n490), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n494), .A2(new_n495), .A3(new_n490), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT86), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n500), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n469), .B1(new_n499), .B2(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n501), .B1(new_n489), .B2(new_n490), .ZN(new_n507));
  AND4_X1   g306(.A1(new_n501), .A2(new_n494), .A3(new_n495), .A4(new_n490), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n472), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n497), .B1(new_n496), .B2(G22gat), .ZN(new_n510));
  AOI211_X1 g309(.A(new_n490), .B(new_n473), .C1(new_n494), .C2(new_n495), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n503), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n509), .A2(new_n512), .A3(KEYINPUT88), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n506), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n326), .B1(new_n468), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n455), .A2(KEYINPUT6), .A3(new_n460), .ZN(new_n516));
  INV_X1    g315(.A(new_n428), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT4), .B1(new_n296), .B2(new_n416), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT78), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n433), .A2(new_n434), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(new_n520), .A3(new_n432), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n427), .B1(new_n451), .B2(new_n452), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n517), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n450), .A2(new_n453), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(new_n427), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n419), .A2(new_n424), .A3(new_n426), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  AOI22_X1  g326(.A1(new_n523), .A2(new_n525), .B1(new_n527), .B2(new_n429), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n462), .B1(new_n528), .B2(new_n463), .ZN(new_n529));
  INV_X1    g328(.A(new_n464), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n381), .B(new_n516), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT37), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n533), .B1(new_n365), .B2(new_n368), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n368), .A2(new_n533), .A3(new_n359), .A4(new_n363), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(new_n373), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT38), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(KEYINPUT90), .B1(new_n378), .B2(new_n348), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT90), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n367), .A2(new_n539), .A3(new_n360), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n361), .B1(new_n362), .B2(new_n357), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(new_n348), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n538), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT38), .B1(new_n543), .B2(KEYINPUT37), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n544), .A2(new_n373), .A3(new_n535), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n532), .A2(new_n537), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n509), .A2(new_n512), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n382), .A2(new_n372), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n527), .A2(KEYINPUT89), .A3(new_n428), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n428), .B1(new_n450), .B2(new_n453), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT39), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT89), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(new_n526), .B2(new_n517), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n551), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n460), .B1(new_n552), .B2(new_n553), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT40), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n557), .A2(new_n558), .A3(KEYINPUT40), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n561), .A2(new_n461), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n548), .B1(new_n550), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n515), .B1(new_n546), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n516), .B1(new_n529), .B2(new_n530), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT35), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n547), .A2(new_n324), .A3(new_n323), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n465), .A2(new_n467), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n319), .A2(new_n320), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n549), .A2(new_n571), .A3(new_n572), .A4(new_n547), .ZN(new_n573));
  AOI22_X1  g372(.A1(new_n549), .A2(new_n570), .B1(new_n573), .B2(KEYINPUT35), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n202), .B1(new_n565), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n514), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n549), .A2(new_n571), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AND3_X1   g377(.A1(new_n532), .A2(new_n537), .A3(new_n545), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n561), .A2(new_n461), .A3(new_n562), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n547), .B1(new_n580), .B2(new_n549), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n578), .B(new_n326), .C1(new_n579), .C2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n570), .A2(new_n549), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n573), .A2(KEYINPUT35), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n582), .A2(new_n585), .A3(KEYINPUT91), .ZN(new_n586));
  XNOR2_X1  g385(.A(G113gat), .B(G141gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(G197gat), .ZN(new_n588));
  XOR2_X1   g387(.A(KEYINPUT11), .B(G169gat), .Z(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(new_n590), .B(KEYINPUT12), .Z(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT92), .B(G36gat), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT14), .ZN(new_n593));
  INV_X1    g392(.A(G29gat), .ZN(new_n594));
  INV_X1    g393(.A(G36gat), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n597));
  AOI22_X1  g396(.A1(new_n592), .A2(G29gat), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(G43gat), .B(G50gat), .Z(new_n599));
  INV_X1    g398(.A(KEYINPUT15), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G43gat), .B(G50gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT15), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n598), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(KEYINPUT94), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT94), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n598), .A2(new_n601), .A3(new_n606), .A4(new_n603), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT93), .ZN(new_n608));
  OR3_X1    g407(.A1(new_n598), .A2(new_n608), .A3(new_n603), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n608), .B1(new_n598), .B2(new_n603), .ZN(new_n610));
  AOI22_X1  g409(.A1(new_n605), .A2(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G15gat), .B(G22gat), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n612), .A2(G1gat), .ZN(new_n613));
  INV_X1    g412(.A(G8gat), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT16), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n612), .B1(new_n615), .B2(G1gat), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n613), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n614), .B1(new_n613), .B2(new_n616), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(KEYINPUT96), .B1(new_n611), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n607), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n609), .A2(new_n610), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT96), .ZN(new_n624));
  INV_X1    g423(.A(new_n619), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n620), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n627), .B1(new_n623), .B2(new_n625), .ZN(new_n628));
  NAND2_X1  g427(.A1(G229gat), .A2(G233gat), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n629), .B(KEYINPUT13), .Z(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT17), .ZN(new_n632));
  OAI21_X1  g431(.A(KEYINPUT95), .B1(new_n623), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT95), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n611), .A2(new_n634), .A3(KEYINPUT17), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n625), .B1(new_n623), .B2(new_n632), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n638), .A2(new_n629), .A3(new_n627), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT18), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n631), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AOI22_X1  g440(.A1(new_n636), .A2(new_n637), .B1(new_n620), .B2(new_n626), .ZN(new_n642));
  AOI21_X1  g441(.A(KEYINPUT18), .B1(new_n642), .B2(new_n629), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n591), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n639), .A2(new_n640), .ZN(new_n645));
  INV_X1    g444(.A(new_n591), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n642), .A2(KEYINPUT18), .A3(new_n629), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n645), .A2(new_n646), .A3(new_n647), .A4(new_n631), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT97), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n644), .A2(KEYINPUT97), .A3(new_n648), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  AND3_X1   g453(.A1(new_n575), .A2(new_n586), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G183gat), .B(G211gat), .ZN(new_n656));
  AND2_X1   g455(.A1(G71gat), .A2(G78gat), .ZN(new_n657));
  NOR2_X1   g456(.A1(G71gat), .A2(G78gat), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n657), .B1(KEYINPUT9), .B2(new_n658), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT98), .B(G57gat), .Z(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(G64gat), .ZN(new_n661));
  INV_X1    g460(.A(G64gat), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(G57gat), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n659), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  XOR2_X1   g463(.A(G57gat), .B(G64gat), .Z(new_n665));
  AOI211_X1 g464(.A(new_n657), .B(new_n658), .C1(new_n665), .C2(KEYINPUT9), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT21), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(G231gat), .A2(G233gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n213), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n671), .A2(new_n213), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n656), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n674), .ZN(new_n676));
  INV_X1    g475(.A(new_n656), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n676), .A2(new_n672), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n667), .A2(new_n668), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n680), .A2(new_n625), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT99), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(new_n385), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  OR2_X1    g484(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n682), .A2(new_n685), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n679), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n675), .A2(new_n678), .A3(new_n686), .A4(new_n687), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(G232gat), .A2(G233gat), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n694), .A2(KEYINPUT41), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT100), .ZN(new_n696));
  XNOR2_X1  g495(.A(G134gat), .B(G162gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n623), .A2(new_n632), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT8), .ZN(new_n701));
  NAND2_X1  g500(.A1(G99gat), .A2(G106gat), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT102), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(KEYINPUT102), .A2(G99gat), .A3(G106gat), .ZN(new_n705));
  INV_X1    g504(.A(G85gat), .ZN(new_n706));
  INV_X1    g505(.A(G92gat), .ZN(new_n707));
  AOI22_X1  g506(.A1(new_n704), .A2(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT103), .ZN(new_n709));
  AOI211_X1 g508(.A(new_n706), .B(new_n707), .C1(KEYINPUT101), .C2(KEYINPUT7), .ZN(new_n710));
  NOR2_X1   g509(.A1(KEYINPUT101), .A2(KEYINPUT7), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  XOR2_X1   g512(.A(G99gat), .B(G106gat), .Z(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n714), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n709), .A2(new_n716), .A3(new_n712), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n636), .A2(new_n700), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(G190gat), .B(G218gat), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT104), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n718), .ZN(new_n723));
  AOI22_X1  g522(.A1(new_n723), .A2(new_n623), .B1(KEYINPUT41), .B2(new_n694), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n719), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n722), .B1(new_n719), .B2(new_n724), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n699), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n719), .A2(new_n724), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n721), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n719), .A2(new_n722), .A3(new_n724), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n729), .A2(new_n698), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(G230gat), .A2(G233gat), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT105), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n667), .B1(new_n717), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n718), .A2(new_n736), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n715), .B(new_n717), .C1(new_n735), .C2(new_n667), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT10), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT10), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n718), .A2(new_n740), .A3(new_n667), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n734), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n734), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n737), .A2(new_n743), .A3(new_n738), .ZN(new_n744));
  XNOR2_X1  g543(.A(G120gat), .B(G148gat), .ZN(new_n745));
  XNOR2_X1  g544(.A(G176gat), .B(G204gat), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n745), .B(new_n746), .Z(new_n747));
  NAND3_X1  g546(.A1(new_n742), .A2(new_n744), .A3(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n747), .B1(new_n742), .B2(new_n744), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n692), .A2(new_n733), .A3(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT106), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n655), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n756), .A2(new_n571), .ZN(new_n757));
  XOR2_X1   g556(.A(new_n757), .B(G1gat), .Z(G1324gat));
  XOR2_X1   g557(.A(KEYINPUT16), .B(G8gat), .Z(new_n759));
  NAND4_X1  g558(.A1(new_n655), .A2(new_n550), .A3(new_n755), .A4(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(G8gat), .B1(new_n756), .B2(new_n549), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(new_n760), .ZN(new_n762));
  MUX2_X1   g561(.A(new_n760), .B(new_n762), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g562(.A(G15gat), .B1(new_n756), .B2(new_n326), .ZN(new_n764));
  INV_X1    g563(.A(new_n572), .ZN(new_n765));
  OR2_X1    g564(.A1(new_n765), .A2(G15gat), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n764), .B1(new_n756), .B2(new_n766), .ZN(G1326gat));
  INV_X1    g566(.A(KEYINPUT107), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(new_n756), .B2(new_n514), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n655), .A2(KEYINPUT107), .A3(new_n576), .A4(new_n755), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g570(.A(KEYINPUT43), .B(G22gat), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n771), .B(new_n772), .ZN(G1327gat));
  INV_X1    g572(.A(new_n751), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n692), .A2(new_n774), .A3(new_n733), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n575), .A2(new_n586), .A3(new_n654), .A4(new_n775), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n776), .A2(G29gat), .A3(new_n571), .ZN(new_n777));
  XOR2_X1   g576(.A(new_n777), .B(KEYINPUT45), .Z(new_n778));
  NAND3_X1  g577(.A1(new_n649), .A2(new_n691), .A3(new_n751), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n575), .A2(new_n586), .A3(new_n732), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT44), .ZN(new_n781));
  AND3_X1   g580(.A1(new_n727), .A2(new_n731), .A3(KEYINPUT109), .ZN(new_n782));
  AOI21_X1  g581(.A(KEYINPUT109), .B1(new_n727), .B2(new_n731), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT44), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n564), .A2(new_n546), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT108), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n578), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n576), .A2(new_n577), .A3(KEYINPUT108), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n787), .A2(new_n789), .A3(new_n326), .A4(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n786), .B1(new_n791), .B2(new_n585), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n779), .B1(new_n781), .B2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(G29gat), .B1(new_n795), .B2(new_n571), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n778), .A2(new_n796), .ZN(G1328gat));
  OAI21_X1  g596(.A(new_n592), .B1(new_n795), .B2(new_n549), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n549), .A2(new_n592), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(KEYINPUT46), .B1(new_n776), .B2(new_n800), .ZN(new_n801));
  OR3_X1    g600(.A1(new_n776), .A2(KEYINPUT46), .A3(new_n800), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n798), .A2(new_n801), .A3(new_n802), .ZN(G1329gat));
  AOI21_X1  g602(.A(new_n792), .B1(new_n780), .B2(KEYINPUT44), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n804), .A2(new_n326), .A3(new_n779), .ZN(new_n805));
  INV_X1    g604(.A(G43gat), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT110), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n655), .A2(new_n806), .A3(new_n572), .A4(new_n775), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n808), .B1(new_n805), .B2(new_n806), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT47), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n807), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  OAI221_X1 g610(.A(new_n808), .B1(KEYINPUT110), .B2(KEYINPUT47), .C1(new_n805), .C2(new_n806), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(G1330gat));
  INV_X1    g612(.A(KEYINPUT48), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n514), .A2(G50gat), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n776), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n817), .B(KEYINPUT111), .ZN(new_n818));
  INV_X1    g617(.A(G50gat), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n819), .B1(new_n794), .B2(new_n576), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n814), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT112), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n822), .B1(new_n794), .B2(new_n548), .ZN(new_n823));
  NOR4_X1   g622(.A1(new_n804), .A2(KEYINPUT112), .A3(new_n547), .A4(new_n779), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n823), .A2(new_n824), .A3(new_n819), .ZN(new_n825));
  OAI21_X1  g624(.A(KEYINPUT48), .B1(new_n776), .B2(new_n816), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n821), .B1(new_n825), .B2(new_n826), .ZN(G1331gat));
  NAND2_X1  g626(.A1(new_n791), .A2(new_n585), .ZN(new_n828));
  NOR4_X1   g627(.A1(new_n649), .A2(new_n751), .A3(new_n691), .A4(new_n732), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(new_n571), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n831), .B(new_n660), .ZN(G1332gat));
  NOR2_X1   g631(.A1(new_n830), .A2(new_n549), .ZN(new_n833));
  NOR2_X1   g632(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n834));
  AND2_X1   g633(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n836), .B1(new_n833), .B2(new_n834), .ZN(G1333gat));
  OR3_X1    g636(.A1(new_n830), .A2(G71gat), .A3(new_n765), .ZN(new_n838));
  OAI21_X1  g637(.A(G71gat), .B1(new_n830), .B2(new_n326), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XOR2_X1   g639(.A(new_n840), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g640(.A1(new_n830), .A2(new_n514), .ZN(new_n842));
  XOR2_X1   g641(.A(KEYINPUT113), .B(G78gat), .Z(new_n843));
  XNOR2_X1  g642(.A(new_n842), .B(new_n843), .ZN(G1335gat));
  NOR3_X1   g643(.A1(new_n692), .A2(new_n649), .A3(new_n733), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT51), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n846), .B(new_n847), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n848), .A2(new_n774), .ZN(new_n849));
  INV_X1    g648(.A(new_n571), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n849), .A2(new_n706), .A3(new_n850), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n692), .A2(new_n649), .A3(new_n751), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT114), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n804), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(G85gat), .B1(new_n854), .B2(new_n571), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n851), .A2(new_n855), .ZN(G1336gat));
  OAI21_X1  g655(.A(G92gat), .B1(new_n854), .B2(new_n549), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT52), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n549), .A2(G92gat), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n848), .A2(new_n774), .A3(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n857), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  AND3_X1   g660(.A1(new_n848), .A2(new_n774), .A3(new_n859), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n804), .A2(new_n853), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n707), .B1(new_n863), .B2(new_n550), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT52), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n861), .A2(new_n865), .ZN(G1337gat));
  INV_X1    g665(.A(G99gat), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n849), .A2(new_n867), .A3(new_n572), .ZN(new_n868));
  OAI21_X1  g667(.A(G99gat), .B1(new_n854), .B2(new_n326), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(G1338gat));
  OAI21_X1  g669(.A(G106gat), .B1(new_n854), .B2(new_n547), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n751), .A2(new_n547), .A3(G106gat), .ZN(new_n872));
  AOI21_X1  g671(.A(KEYINPUT53), .B1(new_n848), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n863), .A2(new_n576), .ZN(new_n875));
  XOR2_X1   g674(.A(new_n872), .B(KEYINPUT115), .Z(new_n876));
  AOI22_X1  g675(.A1(new_n875), .A2(G106gat), .B1(new_n848), .B2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n874), .B1(new_n877), .B2(new_n878), .ZN(G1339gat));
  NOR2_X1   g678(.A1(new_n752), .A2(new_n649), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n737), .A2(new_n738), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n740), .ZN(new_n882));
  INV_X1    g681(.A(new_n741), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n882), .A2(new_n743), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n884), .A2(KEYINPUT54), .A3(new_n742), .ZN(new_n885));
  INV_X1    g684(.A(new_n747), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n887), .B(new_n734), .C1(new_n739), .C2(new_n741), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n885), .A2(KEYINPUT55), .A3(new_n886), .A4(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n748), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n886), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(KEYINPUT55), .B1(new_n892), .B2(new_n885), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n642), .A2(new_n629), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n628), .A2(new_n630), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n590), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n648), .A2(new_n896), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n890), .A2(new_n893), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n784), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n751), .A2(new_n897), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n890), .A2(new_n893), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n900), .B1(new_n901), .B2(new_n649), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n899), .B1(new_n902), .B2(new_n784), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n880), .B1(new_n903), .B2(new_n691), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n904), .A2(new_n571), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n905), .A2(new_n549), .A3(new_n514), .A4(new_n572), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n906), .A2(new_n205), .A3(new_n653), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n905), .A2(new_n547), .A3(new_n572), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT116), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(new_n549), .A3(new_n649), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n907), .B1(new_n910), .B2(new_n205), .ZN(G1340gat));
  NOR3_X1   g710(.A1(new_n906), .A2(new_n206), .A3(new_n751), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n909), .A2(new_n549), .A3(new_n774), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n912), .B1(new_n913), .B2(new_n206), .ZN(G1341gat));
  OAI21_X1  g713(.A(G127gat), .B1(new_n906), .B2(new_n691), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n909), .A2(new_n549), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n692), .A2(new_n213), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(G1342gat));
  NOR2_X1   g717(.A1(new_n733), .A2(G134gat), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n908), .A2(KEYINPUT116), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n908), .A2(KEYINPUT116), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n549), .B(new_n919), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(KEYINPUT56), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT56), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n909), .A2(new_n924), .A3(new_n549), .A4(new_n919), .ZN(new_n925));
  OAI21_X1  g724(.A(G134gat), .B1(new_n906), .B2(new_n733), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n923), .A2(new_n925), .A3(new_n926), .ZN(G1343gat));
  NAND2_X1  g726(.A1(new_n326), .A2(new_n548), .ZN(new_n928));
  NOR4_X1   g727(.A1(new_n904), .A2(new_n571), .A3(new_n550), .A4(new_n928), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n653), .A2(G141gat), .ZN(new_n930));
  AOI21_X1  g729(.A(KEYINPUT58), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT119), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n326), .A2(new_n850), .A3(new_n549), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT55), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n884), .A2(KEYINPUT54), .A3(new_n742), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n935), .B1(new_n936), .B2(new_n891), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n649), .A2(new_n937), .A3(new_n748), .A4(new_n889), .ZN(new_n938));
  INV_X1    g737(.A(new_n897), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n774), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n784), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n939), .A2(new_n937), .A3(new_n748), .A4(new_n889), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT109), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n732), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n727), .A2(new_n731), .A3(KEYINPUT109), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n942), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n691), .B1(new_n941), .B2(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(new_n880), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n547), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n950), .A2(KEYINPUT57), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n576), .A2(KEYINPUT57), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT117), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n953), .B1(new_n936), .B2(new_n891), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n892), .A2(KEYINPUT117), .A3(new_n885), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n954), .A2(new_n935), .A3(new_n955), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n889), .A2(new_n748), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n956), .A2(new_n651), .A3(new_n957), .A4(new_n652), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n732), .B1(new_n958), .B2(new_n940), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n691), .B1(new_n959), .B2(new_n947), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n952), .B1(new_n960), .B2(new_n949), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n934), .B1(new_n951), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n932), .B1(new_n962), .B2(new_n653), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(G141gat), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n962), .A2(new_n932), .A3(new_n653), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n931), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI211_X1 g765(.A(new_n649), .B(new_n934), .C1(new_n951), .C2(new_n961), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(G141gat), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n929), .A2(new_n930), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g769(.A(KEYINPUT118), .B1(new_n970), .B2(KEYINPUT58), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT118), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT58), .ZN(new_n973));
  AOI211_X1 g772(.A(new_n972), .B(new_n973), .C1(new_n968), .C2(new_n969), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n966), .B1(new_n971), .B2(new_n974), .ZN(G1344gat));
  INV_X1    g774(.A(G148gat), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n929), .A2(new_n976), .A3(new_n774), .ZN(new_n977));
  INV_X1    g776(.A(new_n962), .ZN(new_n978));
  AOI211_X1 g777(.A(KEYINPUT59), .B(new_n976), .C1(new_n978), .C2(new_n774), .ZN(new_n979));
  XNOR2_X1  g778(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n514), .A2(KEYINPUT57), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n958), .A2(new_n940), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(new_n733), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n898), .A2(new_n732), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n692), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n754), .A2(new_n654), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n981), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g786(.A(KEYINPUT57), .B1(new_n904), .B2(new_n547), .ZN(new_n988));
  NAND4_X1  g787(.A1(new_n987), .A2(new_n988), .A3(new_n774), .A4(new_n934), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n980), .B1(new_n989), .B2(G148gat), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n977), .B1(new_n979), .B2(new_n990), .ZN(G1345gat));
  OAI21_X1  g790(.A(G155gat), .B1(new_n962), .B2(new_n691), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n929), .A2(new_n385), .A3(new_n692), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n992), .A2(new_n993), .ZN(G1346gat));
  NAND3_X1  g793(.A1(new_n929), .A2(new_n386), .A3(new_n732), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n978), .A2(new_n784), .ZN(new_n996));
  INV_X1    g795(.A(new_n996), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n995), .B1(new_n997), .B2(new_n386), .ZN(G1347gat));
  INV_X1    g797(.A(new_n904), .ZN(new_n999));
  NOR2_X1   g798(.A1(new_n850), .A2(new_n549), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n1000), .A2(new_n572), .ZN(new_n1001));
  AND2_X1   g800(.A1(new_n1001), .A2(KEYINPUT121), .ZN(new_n1002));
  NOR2_X1   g801(.A1(new_n1002), .A2(new_n576), .ZN(new_n1003));
  OAI211_X1 g802(.A(new_n999), .B(new_n1003), .C1(KEYINPUT121), .C2(new_n1001), .ZN(new_n1004));
  INV_X1    g803(.A(G169gat), .ZN(new_n1005));
  NOR3_X1   g804(.A1(new_n1004), .A2(new_n1005), .A3(new_n653), .ZN(new_n1006));
  NOR4_X1   g805(.A1(new_n904), .A2(new_n850), .A3(new_n549), .A4(new_n569), .ZN(new_n1007));
  AOI21_X1  g806(.A(G169gat), .B1(new_n1007), .B2(new_n649), .ZN(new_n1008));
  NOR2_X1   g807(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g808(.A(new_n1009), .B(KEYINPUT122), .ZN(G1348gat));
  INV_X1    g809(.A(G176gat), .ZN(new_n1011));
  NOR2_X1   g810(.A1(new_n751), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g811(.A(new_n1012), .ZN(new_n1013));
  OR3_X1    g812(.A1(new_n1004), .A2(KEYINPUT123), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1007), .A2(new_n774), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n1015), .A2(new_n1011), .ZN(new_n1016));
  OAI21_X1  g815(.A(KEYINPUT123), .B1(new_n1004), .B2(new_n1013), .ZN(new_n1017));
  NAND3_X1  g816(.A1(new_n1014), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g817(.A1(new_n1018), .A2(KEYINPUT124), .ZN(new_n1019));
  INV_X1    g818(.A(KEYINPUT124), .ZN(new_n1020));
  NAND4_X1  g819(.A1(new_n1014), .A2(new_n1020), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1021));
  NAND2_X1  g820(.A1(new_n1019), .A2(new_n1021), .ZN(G1349gat));
  OAI21_X1  g821(.A(G183gat), .B1(new_n1004), .B2(new_n691), .ZN(new_n1023));
  NAND3_X1  g822(.A1(new_n1007), .A2(new_n261), .A3(new_n692), .ZN(new_n1024));
  NAND2_X1  g823(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g824(.A(new_n1025), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g825(.A1(new_n1007), .A2(new_n262), .A3(new_n784), .ZN(new_n1027));
  OAI21_X1  g826(.A(G190gat), .B1(new_n1004), .B2(new_n733), .ZN(new_n1028));
  AND2_X1   g827(.A1(new_n1028), .A2(KEYINPUT61), .ZN(new_n1029));
  NOR2_X1   g828(.A1(new_n1028), .A2(KEYINPUT61), .ZN(new_n1030));
  OAI21_X1  g829(.A(new_n1027), .B1(new_n1029), .B2(new_n1030), .ZN(G1351gat));
  NOR2_X1   g830(.A1(new_n904), .A2(new_n850), .ZN(new_n1032));
  NOR2_X1   g831(.A1(new_n928), .A2(new_n549), .ZN(new_n1033));
  AND2_X1   g832(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g833(.A(G197gat), .B1(new_n1034), .B2(new_n649), .ZN(new_n1035));
  NAND2_X1  g834(.A1(new_n987), .A2(new_n988), .ZN(new_n1036));
  NAND2_X1  g835(.A1(new_n1000), .A2(new_n326), .ZN(new_n1037));
  XNOR2_X1  g836(.A(new_n1037), .B(KEYINPUT125), .ZN(new_n1038));
  NOR2_X1   g837(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g838(.A1(new_n653), .A2(new_n331), .ZN(new_n1040));
  AOI21_X1  g839(.A(new_n1035), .B1(new_n1039), .B2(new_n1040), .ZN(G1352gat));
  INV_X1    g840(.A(KEYINPUT126), .ZN(new_n1042));
  AOI21_X1  g841(.A(new_n332), .B1(new_n1039), .B2(new_n774), .ZN(new_n1043));
  NAND4_X1  g842(.A1(new_n1032), .A2(new_n332), .A3(new_n774), .A4(new_n1033), .ZN(new_n1044));
  XNOR2_X1  g843(.A(new_n1044), .B(KEYINPUT62), .ZN(new_n1045));
  OAI21_X1  g844(.A(new_n1042), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g845(.A(KEYINPUT62), .ZN(new_n1047));
  XNOR2_X1  g846(.A(new_n1044), .B(new_n1047), .ZN(new_n1048));
  NOR3_X1   g847(.A1(new_n1036), .A2(new_n751), .A3(new_n1038), .ZN(new_n1049));
  OAI211_X1 g848(.A(new_n1048), .B(KEYINPUT126), .C1(new_n332), .C2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g849(.A1(new_n1046), .A2(new_n1050), .ZN(G1353gat));
  NAND3_X1  g850(.A1(new_n1034), .A2(new_n336), .A3(new_n692), .ZN(new_n1052));
  NOR2_X1   g851(.A1(new_n1037), .A2(new_n691), .ZN(new_n1053));
  NAND3_X1  g852(.A1(new_n987), .A2(new_n988), .A3(new_n1053), .ZN(new_n1054));
  AND3_X1   g853(.A1(new_n1054), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1055));
  AOI21_X1  g854(.A(KEYINPUT63), .B1(new_n1054), .B2(G211gat), .ZN(new_n1056));
  OAI21_X1  g855(.A(new_n1052), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g856(.A(KEYINPUT127), .ZN(new_n1058));
  NAND2_X1  g857(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  OAI211_X1 g858(.A(KEYINPUT127), .B(new_n1052), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1060));
  NAND2_X1  g859(.A1(new_n1059), .A2(new_n1060), .ZN(G1354gat));
  NAND3_X1  g860(.A1(new_n1034), .A2(new_n337), .A3(new_n784), .ZN(new_n1062));
  NOR3_X1   g861(.A1(new_n1036), .A2(new_n733), .A3(new_n1038), .ZN(new_n1063));
  OAI21_X1  g862(.A(new_n1062), .B1(new_n1063), .B2(new_n337), .ZN(G1355gat));
endmodule


