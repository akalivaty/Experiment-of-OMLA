//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 1 0 1 1 0 1 0 0 1 1 0 0 1 1 1 1 0 0 0 0 0 1 0 0 0 1 0 1 1 0 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n560, new_n561, new_n562, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT67), .Z(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n460), .A2(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G101), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G137), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(KEYINPUT68), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(new_n460), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n470), .A2(new_n475), .A3(G125), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n467), .B1(new_n478), .B2(G2105), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT69), .ZN(G160));
  NAND2_X1  g055(.A1(new_n463), .A2(G2105), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT70), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G112), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(G2105), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n468), .A2(new_n469), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n487), .B1(new_n489), .B2(G136), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n484), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR3_X1   g068(.A1(new_n493), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n470), .A2(new_n475), .A3(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT72), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g072(.A(G138), .B(new_n464), .C1(new_n468), .C2(new_n469), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT71), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n470), .A2(new_n475), .A3(KEYINPUT72), .A4(new_n494), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n498), .A2(new_n502), .A3(KEYINPUT4), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n497), .A2(new_n500), .A3(new_n501), .A4(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n505));
  INV_X1    g080(.A(G114), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(G2105), .ZN(new_n507));
  INV_X1    g082(.A(new_n481), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(G126), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(G164));
  AND2_X1   g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  OR2_X1    g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT74), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NOR3_X1   g092(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AND2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n518), .B1(G50), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n516), .B1(new_n515), .B2(new_n517), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n512), .A2(new_n513), .ZN(new_n526));
  OR3_X1    g101(.A1(new_n526), .A2(new_n521), .A3(KEYINPUT73), .ZN(new_n527));
  OAI21_X1  g102(.A(KEYINPUT73), .B1(new_n526), .B2(new_n521), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G88), .ZN(new_n530));
  AND3_X1   g105(.A1(new_n524), .A2(new_n525), .A3(new_n530), .ZN(G166));
  NAND2_X1  g106(.A1(new_n529), .A2(G89), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  NAND2_X1  g109(.A1(G63), .A2(G651), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n526), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n536), .B1(G51), .B2(new_n523), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n532), .A2(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G64), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n526), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n542), .A2(G651), .B1(new_n523), .B2(G52), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n527), .A2(new_n528), .ZN(new_n544));
  INV_X1    g119(.A(G90), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  NAND2_X1  g122(.A1(new_n529), .A2(G81), .ZN(new_n548));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G56), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n526), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT75), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n517), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n553), .B1(new_n552), .B2(new_n551), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n523), .A2(G43), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n548), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g134(.A(KEYINPUT76), .B(KEYINPUT8), .Z(new_n560));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n560), .B(new_n561), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  NAND3_X1  g138(.A1(new_n527), .A2(G91), .A3(new_n528), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT77), .ZN(new_n565));
  INV_X1    g140(.A(new_n523), .ZN(new_n566));
  INV_X1    g141(.A(G53), .ZN(new_n567));
  OR3_X1    g142(.A1(new_n566), .A2(KEYINPUT9), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g143(.A(KEYINPUT9), .B1(new_n566), .B2(new_n567), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n526), .B2(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n568), .A2(new_n569), .B1(G651), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n565), .A2(new_n573), .ZN(G299));
  NAND3_X1  g149(.A1(new_n524), .A2(new_n525), .A3(new_n530), .ZN(G303));
  NAND2_X1  g150(.A1(new_n529), .A2(G87), .ZN(new_n576));
  OR2_X1    g151(.A1(new_n514), .A2(G74), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n577), .A2(G651), .B1(G49), .B2(new_n523), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(G288));
  NAND3_X1  g154(.A1(new_n527), .A2(G86), .A3(new_n528), .ZN(new_n580));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G61), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n526), .B2(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n583), .A2(G651), .B1(new_n523), .B2(G48), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n585), .A2(KEYINPUT78), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(KEYINPUT78), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G305));
  NAND2_X1  g164(.A1(new_n529), .A2(G85), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT79), .ZN(new_n591));
  NAND2_X1  g166(.A1(G72), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G60), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n526), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n594), .A2(G651), .B1(new_n523), .B2(G47), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n590), .A2(new_n591), .A3(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n591), .B1(new_n590), .B2(new_n595), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  XOR2_X1   g176(.A(new_n601), .B(KEYINPUT80), .Z(new_n602));
  NAND2_X1  g177(.A1(new_n523), .A2(G54), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n514), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(new_n517), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n529), .A2(G92), .ZN(new_n606));
  XNOR2_X1  g181(.A(KEYINPUT81), .B(KEYINPUT10), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n607), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n529), .A2(G92), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n602), .B1(G868), .B2(new_n612), .ZN(G321));
  XNOR2_X1  g188(.A(G321), .B(KEYINPUT82), .ZN(G284));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  INV_X1    g190(.A(G299), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G297));
  OAI21_X1  g192(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n612), .B1(new_n619), .B2(G860), .ZN(G148));
  NAND2_X1  g195(.A1(new_n612), .A2(new_n619), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G868), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n557), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g199(.A1(new_n470), .A2(new_n475), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(new_n461), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  INV_X1    g203(.A(G2100), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n489), .A2(G135), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n464), .A2(G111), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  INV_X1    g209(.A(G123), .ZN(new_n635));
  OAI221_X1 g210(.A(new_n632), .B1(new_n633), .B2(new_n634), .C1(new_n482), .C2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NAND3_X1  g212(.A1(new_n630), .A2(new_n631), .A3(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2435), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT83), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2427), .B(G2430), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n641), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(KEYINPUT14), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2451), .B(G2454), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n648), .B(new_n649), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n646), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  AND2_X1   g228(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g229(.A(G14), .B1(new_n651), .B2(new_n653), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(G401));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT84), .ZN(new_n659));
  NOR2_X1   g234(.A1(G2072), .A2(G2078), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n442), .A2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n657), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n661), .B(KEYINPUT17), .Z(new_n664));
  OAI21_X1  g239(.A(new_n663), .B1(new_n664), .B2(new_n659), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n661), .A2(new_n657), .A3(new_n658), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT18), .Z(new_n667));
  NAND3_X1  g242(.A1(new_n664), .A2(new_n659), .A3(new_n657), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n665), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(new_n629), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT85), .B(G2096), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G227));
  XOR2_X1   g247(.A(G1991), .B(G1996), .Z(new_n673));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT19), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  XOR2_X1   g252(.A(G1961), .B(G1966), .Z(new_n678));
  AND2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT20), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n677), .A2(new_n678), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n676), .A2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT86), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  OR3_X1    g260(.A1(new_n676), .A2(new_n679), .A3(new_n682), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n681), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT87), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g264(.A1(new_n681), .A2(new_n685), .A3(KEYINPUT87), .A4(new_n686), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n691), .B1(new_n689), .B2(new_n690), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n673), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n694), .ZN(new_n696));
  INV_X1    g271(.A(new_n673), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n696), .A2(new_n697), .A3(new_n692), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1981), .B(G1986), .ZN(new_n699));
  AND3_X1   g274(.A1(new_n695), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n699), .B1(new_n695), .B2(new_n698), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(G229));
  INV_X1    g277(.A(G16), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G22), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G166), .B2(new_n703), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(G1971), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT33), .B(G1976), .Z(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n703), .A2(G23), .ZN(new_n709));
  INV_X1    g284(.A(G288), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(new_n703), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT88), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n706), .B1(new_n708), .B2(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(G6), .A2(G16), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(new_n588), .B2(G16), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT32), .B(G1981), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n712), .A2(new_n708), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n713), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(KEYINPUT34), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT34), .ZN(new_n721));
  NAND4_X1  g296(.A1(new_n713), .A2(new_n721), .A3(new_n717), .A4(new_n718), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n703), .A2(G24), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(new_n599), .B2(new_n703), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G1986), .ZN(new_n725));
  INV_X1    g300(.A(G29), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G25), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n483), .A2(G119), .ZN(new_n728));
  OAI21_X1  g303(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n729));
  INV_X1    g304(.A(G107), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(G2105), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n489), .B2(G131), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n728), .A2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n727), .B1(new_n734), .B2(new_n726), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT35), .B(G1991), .Z(new_n736));
  XOR2_X1   g311(.A(new_n735), .B(new_n736), .Z(new_n737));
  NOR2_X1   g312(.A1(new_n725), .A2(new_n737), .ZN(new_n738));
  AND3_X1   g313(.A1(new_n722), .A2(KEYINPUT89), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(KEYINPUT89), .B1(new_n722), .B2(new_n738), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n720), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(KEYINPUT36), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT36), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n743), .B(new_n720), .C1(new_n739), .C2(new_n740), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n489), .A2(G141), .ZN(new_n746));
  NAND3_X1  g321(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT26), .Z(new_n748));
  NAND3_X1  g323(.A1(new_n464), .A2(G105), .A3(G2104), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT92), .ZN(new_n750));
  AND3_X1   g325(.A1(new_n746), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G129), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n751), .B1(new_n752), .B2(new_n482), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n753), .A2(KEYINPUT93), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(KEYINPUT93), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n757), .A2(new_n726), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n726), .B2(G32), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT27), .B(G1996), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n703), .A2(G5), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G171), .B2(new_n703), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT94), .Z(new_n763));
  OAI22_X1  g338(.A1(new_n759), .A2(new_n760), .B1(G1961), .B2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(G2084), .ZN(new_n765));
  NAND2_X1  g340(.A1(G160), .A2(G29), .ZN(new_n766));
  INV_X1    g341(.A(G34), .ZN(new_n767));
  AOI21_X1  g342(.A(G29), .B1(new_n767), .B2(KEYINPUT24), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(KEYINPUT24), .B2(new_n767), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n764), .B1(new_n765), .B2(new_n770), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT95), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n703), .A2(G20), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT23), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n616), .B2(new_n703), .ZN(new_n775));
  INV_X1    g350(.A(G1956), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(G16), .A2(G19), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n557), .B2(G16), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT90), .B(G1341), .Z(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n726), .A2(G33), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n625), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n783), .A2(new_n464), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT25), .Z(new_n786));
  INV_X1    g361(.A(G139), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(new_n787), .B2(new_n465), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n784), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n782), .B1(new_n789), .B2(new_n726), .ZN(new_n790));
  AOI22_X1  g365(.A1(new_n779), .A2(new_n781), .B1(G2072), .B2(new_n790), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n790), .A2(G2072), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n791), .B(new_n792), .C1(new_n779), .C2(new_n781), .ZN(new_n793));
  INV_X1    g368(.A(new_n770), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n793), .B1(G2084), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n759), .A2(new_n760), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n763), .A2(G1961), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n612), .A2(G16), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G4), .B2(G16), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(G1348), .ZN(new_n801));
  NAND2_X1  g376(.A1(G164), .A2(G29), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G27), .B2(G29), .ZN(new_n803));
  INV_X1    g378(.A(G2078), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n796), .A2(new_n797), .A3(new_n801), .A4(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT30), .B(G28), .ZN(new_n807));
  OR2_X1    g382(.A1(KEYINPUT31), .A2(G11), .ZN(new_n808));
  NAND2_X1  g383(.A1(KEYINPUT31), .A2(G11), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n807), .A2(new_n726), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n726), .A2(KEYINPUT28), .A3(G26), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT28), .ZN(new_n812));
  INV_X1    g387(.A(G26), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n812), .B1(new_n813), .B2(G29), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n483), .A2(G128), .ZN(new_n815));
  OAI21_X1  g390(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n816));
  INV_X1    g391(.A(G116), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(G2105), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(new_n489), .B2(G140), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n811), .B(new_n814), .C1(new_n821), .C2(new_n726), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT91), .B(G2067), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  OAI221_X1 g399(.A(new_n810), .B1(new_n726), .B2(new_n636), .C1(new_n822), .C2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n703), .A2(G21), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(G168), .B2(new_n703), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(G1966), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(G29), .A2(G35), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(G162), .B2(G29), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT29), .B(G2090), .ZN(new_n832));
  AOI22_X1  g407(.A1(new_n822), .A2(new_n824), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n829), .B(new_n833), .C1(new_n831), .C2(new_n832), .ZN(new_n834));
  OAI22_X1  g409(.A1(new_n800), .A2(G1348), .B1(new_n804), .B2(new_n803), .ZN(new_n835));
  NOR3_X1   g410(.A1(new_n806), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  AND4_X1   g411(.A1(new_n772), .A2(new_n777), .A3(new_n795), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n745), .A2(new_n837), .ZN(G150));
  INV_X1    g413(.A(G150), .ZN(G311));
  AOI22_X1  g414(.A1(new_n529), .A2(G93), .B1(G55), .B2(new_n523), .ZN(new_n840));
  NAND2_X1  g415(.A1(G80), .A2(G543), .ZN(new_n841));
  INV_X1    g416(.A(G67), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n841), .B1(new_n526), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n517), .B1(new_n843), .B2(KEYINPUT97), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(KEYINPUT97), .B2(new_n843), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(G860), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT37), .Z(new_n848));
  NOR2_X1   g423(.A1(new_n611), .A2(new_n619), .ZN(new_n849));
  XOR2_X1   g424(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT98), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n849), .B(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n846), .A2(new_n556), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n846), .A2(new_n556), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n852), .B(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n857), .A2(KEYINPUT39), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT99), .Z(new_n859));
  AOI21_X1  g434(.A(G860), .B1(new_n857), .B2(KEYINPUT39), .ZN(new_n860));
  AND3_X1   g435(.A1(new_n859), .A2(KEYINPUT100), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(KEYINPUT100), .B1(new_n859), .B2(new_n860), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n848), .B1(new_n861), .B2(new_n862), .ZN(G145));
  NAND2_X1  g438(.A1(new_n756), .A2(new_n820), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n754), .A2(new_n821), .A3(new_n755), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n864), .A2(new_n510), .A3(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n510), .B1(new_n864), .B2(new_n865), .ZN(new_n868));
  OAI22_X1  g443(.A1(new_n867), .A2(new_n868), .B1(new_n784), .B2(new_n788), .ZN(new_n869));
  INV_X1    g444(.A(new_n868), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n870), .A2(new_n789), .A3(new_n866), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n489), .A2(G142), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n464), .A2(G118), .ZN(new_n874));
  OAI21_X1  g449(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n876), .B1(new_n483), .B2(G130), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n627), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n734), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n872), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT101), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n869), .A2(new_n871), .A3(new_n879), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(G160), .B(new_n636), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n491), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n869), .A2(new_n871), .A3(KEYINPUT101), .A4(new_n879), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n884), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n883), .A2(new_n886), .ZN(new_n890));
  AOI21_X1  g465(.A(G37), .B1(new_n890), .B2(new_n881), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n892), .B(new_n893), .ZN(G395));
  NAND2_X1  g469(.A1(new_n611), .A2(G299), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n608), .A2(new_n565), .A3(new_n573), .A4(new_n610), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(KEYINPUT103), .B1(new_n897), .B2(KEYINPUT41), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(KEYINPUT41), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT41), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n895), .A2(new_n900), .A3(new_n896), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n898), .B1(new_n902), .B2(KEYINPUT103), .ZN(new_n903));
  XOR2_X1   g478(.A(new_n856), .B(new_n621), .Z(new_n904));
  AND2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  XOR2_X1   g480(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n906));
  INV_X1    g481(.A(new_n897), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  OR3_X1    g483(.A1(new_n905), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(G166), .A2(new_n586), .A3(new_n587), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n588), .A2(G303), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(KEYINPUT104), .ZN(new_n913));
  OAI21_X1  g488(.A(G288), .B1(new_n597), .B2(new_n598), .ZN(new_n914));
  INV_X1    g489(.A(new_n598), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n915), .A2(new_n710), .A3(new_n596), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT104), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n910), .A2(new_n911), .A3(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n913), .A2(new_n918), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n917), .A2(new_n912), .A3(KEYINPUT104), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n906), .B1(new_n905), .B2(new_n908), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n909), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n923), .B1(new_n909), .B2(new_n924), .ZN(new_n926));
  OAI21_X1  g501(.A(G868), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n846), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n927), .B1(G868), .B2(new_n928), .ZN(G295));
  OAI21_X1  g504(.A(new_n927), .B1(G868), .B2(new_n928), .ZN(G331));
  NAND2_X1  g505(.A1(new_n921), .A2(new_n922), .ZN(new_n931));
  INV_X1    g506(.A(new_n901), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n900), .B1(new_n895), .B2(new_n896), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT103), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n898), .ZN(new_n935));
  XNOR2_X1  g510(.A(G286), .B(G301), .ZN(new_n936));
  INV_X1    g511(.A(new_n855), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n936), .B1(new_n937), .B2(new_n853), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT106), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n856), .A2(KEYINPUT106), .A3(new_n936), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n936), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n943), .A2(new_n855), .A3(new_n854), .ZN(new_n944));
  AOI22_X1  g519(.A1(new_n934), .A2(new_n935), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n944), .A2(new_n907), .A3(new_n938), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n931), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G37), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n856), .A2(new_n936), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n950), .B1(new_n940), .B2(new_n941), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n923), .B(new_n946), .C1(new_n903), .C2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n948), .A2(new_n949), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT43), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n944), .A2(new_n907), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n955), .B1(new_n940), .B2(new_n941), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n944), .A2(new_n938), .B1(new_n899), .B2(new_n901), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n931), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT43), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n952), .A2(new_n958), .A3(new_n959), .A4(new_n949), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n954), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n948), .A2(new_n959), .A3(new_n952), .A4(new_n949), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n964), .A2(KEYINPUT44), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n952), .A2(new_n958), .A3(new_n949), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(KEYINPUT107), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT107), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n952), .A2(new_n958), .A3(new_n968), .A4(new_n949), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n967), .A2(KEYINPUT43), .A3(new_n969), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n965), .A2(new_n970), .A3(KEYINPUT108), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT108), .B1(new_n965), .B2(new_n970), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n963), .B1(new_n971), .B2(new_n972), .ZN(G397));
  AOI21_X1  g548(.A(G1384), .B1(new_n504), .B2(new_n509), .ZN(new_n974));
  OR2_X1    g549(.A1(new_n974), .A2(KEYINPUT45), .ZN(new_n975));
  INV_X1    g550(.A(G1996), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n478), .A2(G2105), .ZN(new_n977));
  INV_X1    g552(.A(new_n467), .ZN(new_n978));
  XNOR2_X1  g553(.A(KEYINPUT109), .B(G40), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n977), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT110), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT110), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n479), .A2(new_n983), .A3(new_n980), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n974), .A2(KEYINPUT45), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n975), .A2(new_n976), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n985), .A2(new_n974), .ZN(new_n988));
  XOR2_X1   g563(.A(KEYINPUT58), .B(G1341), .Z(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n556), .B1(new_n987), .B2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n991), .B(KEYINPUT59), .ZN(new_n992));
  XOR2_X1   g567(.A(G299), .B(KEYINPUT57), .Z(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G1384), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n510), .A2(new_n995), .ZN(new_n996));
  AOI22_X1  g571(.A1(new_n996), .A2(KEYINPUT50), .B1(new_n982), .B2(new_n984), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT115), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n510), .A2(new_n999), .A3(new_n995), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT116), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n974), .A2(KEYINPUT116), .A3(new_n999), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n997), .A2(new_n998), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n983), .B1(new_n479), .B2(new_n980), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n464), .B1(new_n476), .B2(new_n477), .ZN(new_n1006));
  NOR4_X1   g581(.A1(new_n1006), .A2(new_n467), .A3(KEYINPUT110), .A4(new_n979), .ZN(new_n1007));
  OAI22_X1  g582(.A1(new_n999), .A2(new_n974), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT115), .ZN(new_n1009));
  AOI21_X1  g584(.A(G1956), .B1(new_n1004), .B2(new_n1009), .ZN(new_n1010));
  OAI22_X1  g585(.A1(KEYINPUT45), .A2(new_n974), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n974), .A2(KEYINPUT45), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g588(.A(KEYINPUT56), .B(G2072), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n994), .B1(new_n1010), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n997), .A2(new_n998), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1018), .A2(new_n1009), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(new_n776), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1021), .A2(new_n993), .A3(new_n1015), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1017), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT61), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n992), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1017), .A2(new_n1022), .A3(KEYINPUT61), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT118), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n996), .A2(new_n1029), .A3(KEYINPUT50), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT112), .B1(new_n974), .B2(new_n999), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1030), .A2(new_n1031), .A3(new_n985), .A4(new_n1000), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G1348), .ZN(new_n1035));
  AOI22_X1  g610(.A1(new_n984), .A2(new_n982), .B1(new_n974), .B2(new_n999), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1036), .A2(new_n1030), .A3(KEYINPUT117), .A4(new_n1031), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1034), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G2067), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n985), .A2(new_n1039), .A3(new_n974), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1038), .A2(KEYINPUT60), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(new_n611), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT60), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1038), .A2(KEYINPUT60), .A3(new_n612), .A4(new_n1040), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1042), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1017), .A2(new_n1022), .A3(KEYINPUT118), .A4(KEYINPUT61), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1025), .A2(new_n1028), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1017), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n611), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1022), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G1971), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1054), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT111), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g632(.A(KEYINPUT111), .B(new_n1054), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1058));
  INV_X1    g633(.A(G2090), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1036), .A2(new_n1030), .A3(new_n1059), .A4(new_n1031), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1057), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(G303), .A2(G8), .ZN(new_n1062));
  AND2_X1   g637(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1063));
  NOR2_X1   g638(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1062), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1065), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1061), .A2(G8), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT114), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n585), .A2(G1981), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n585), .A2(G1981), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1068), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT49), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT49), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1068), .B(new_n1073), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1072), .A2(G8), .A3(new_n988), .A4(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n710), .A2(G1976), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n988), .A2(new_n1076), .A3(G8), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT52), .ZN(new_n1078));
  INV_X1    g653(.A(G1976), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT52), .B1(G288), .B2(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n988), .A2(new_n1076), .A3(new_n1080), .A4(G8), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1075), .A2(new_n1078), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1067), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1004), .A2(new_n1059), .A3(new_n1009), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n1055), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1066), .B1(new_n1085), .B2(G8), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1013), .A2(new_n804), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT53), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(G301), .ZN(new_n1091));
  INV_X1    g666(.A(G1961), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1034), .A2(new_n1092), .A3(new_n1037), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1013), .A2(KEYINPUT53), .A3(new_n804), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1093), .A2(KEYINPUT120), .A3(new_n1094), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1091), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n479), .A2(G40), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1100), .B1(new_n974), .B2(KEYINPUT45), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT121), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n1101), .B(new_n1102), .ZN(new_n1103));
  NOR3_X1   g678(.A1(new_n1012), .A2(new_n1089), .A3(G2078), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1093), .A2(new_n1090), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(G171), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT54), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1087), .B1(new_n1099), .B2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1036), .A2(new_n1030), .A3(new_n765), .A4(new_n1031), .ZN(new_n1110));
  INV_X1    g685(.A(G1966), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1111), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1110), .A2(new_n1112), .A3(G168), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(G8), .ZN(new_n1114));
  AOI21_X1  g689(.A(G168), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT51), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT51), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1113), .A2(new_n1117), .A3(G8), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(KEYINPUT119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT119), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1116), .A2(new_n1121), .A3(new_n1118), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1109), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT54), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1126));
  AOI21_X1  g701(.A(G301), .B1(new_n1126), .B2(new_n1090), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1106), .A2(G171), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1125), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1053), .A2(new_n1124), .A3(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1120), .A2(KEYINPUT62), .A3(new_n1122), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT122), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1120), .A2(KEYINPUT122), .A3(KEYINPUT62), .A4(new_n1122), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT62), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1122), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1121), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1135), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  AOI22_X1  g713(.A1(new_n1097), .A2(new_n1098), .B1(new_n1089), .B2(new_n1088), .ZN(new_n1139));
  INV_X1    g714(.A(G8), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1140), .B1(new_n1084), .B2(new_n1055), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1067), .B(new_n1082), .C1(new_n1141), .C2(new_n1066), .ZN(new_n1142));
  NOR3_X1   g717(.A1(new_n1139), .A2(new_n1142), .A3(G301), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1133), .A2(new_n1134), .A3(new_n1138), .A4(new_n1143), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1061), .A2(G8), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1145), .A2(new_n1066), .A3(new_n1082), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1075), .A2(new_n1079), .A3(new_n710), .ZN(new_n1147));
  OAI211_X1 g722(.A(G8), .B(new_n988), .C1(new_n1147), .C2(new_n1070), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  AOI211_X1 g724(.A(new_n1140), .B(G286), .C1(new_n1110), .C2(new_n1112), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1087), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT63), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1145), .A2(new_n1066), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1150), .A2(KEYINPUT63), .ZN(new_n1155));
  OR3_X1    g730(.A1(new_n1154), .A2(new_n1083), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1149), .B1(new_n1153), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1130), .A2(new_n1144), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n975), .B1(new_n984), .B2(new_n982), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n820), .B(new_n1039), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1160), .B1(new_n757), .B2(new_n976), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1161), .B1(new_n976), .B2(new_n757), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n734), .A2(new_n736), .ZN(new_n1163));
  OR2_X1    g738(.A1(new_n734), .A2(new_n736), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  XOR2_X1   g740(.A(new_n599), .B(G1986), .Z(new_n1166));
  OAI21_X1  g741(.A(new_n1159), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1158), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1159), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1163), .B(KEYINPUT123), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1162), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n821), .A2(new_n1039), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1169), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  OR3_X1    g748(.A1(new_n1169), .A2(G1986), .A3(G290), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1174), .ZN(new_n1175));
  AOI22_X1  g750(.A1(new_n1165), .A2(new_n1159), .B1(new_n1175), .B2(KEYINPUT48), .ZN(new_n1176));
  OR2_X1    g751(.A1(new_n1175), .A2(KEYINPUT48), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1173), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(KEYINPUT46), .B1(new_n1159), .B2(new_n976), .ZN(new_n1179));
  AND2_X1   g754(.A1(new_n1179), .A2(KEYINPUT124), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1179), .A2(KEYINPUT124), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n756), .B1(KEYINPUT46), .B2(new_n976), .ZN(new_n1182));
  AND2_X1   g757(.A1(new_n1182), .A2(new_n1160), .ZN(new_n1183));
  OAI22_X1  g758(.A1(new_n1180), .A2(new_n1181), .B1(new_n1169), .B2(new_n1183), .ZN(new_n1184));
  XOR2_X1   g759(.A(new_n1184), .B(KEYINPUT125), .Z(new_n1185));
  INV_X1    g760(.A(KEYINPUT47), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1178), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1187), .B1(new_n1186), .B2(new_n1185), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1168), .A2(new_n1188), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g764(.A(G319), .B1(new_n654), .B2(new_n655), .ZN(new_n1191));
  NOR2_X1   g765(.A1(G227), .A2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g766(.A(new_n1192), .B1(new_n700), .B2(new_n701), .ZN(new_n1193));
  INV_X1    g767(.A(KEYINPUT126), .ZN(new_n1194));
  NAND2_X1  g768(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  OAI211_X1 g769(.A(KEYINPUT126), .B(new_n1192), .C1(new_n700), .C2(new_n701), .ZN(new_n1196));
  AOI22_X1  g770(.A1(new_n889), .A2(new_n891), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  AND3_X1   g771(.A1(new_n1197), .A2(new_n961), .A3(KEYINPUT127), .ZN(new_n1198));
  AOI21_X1  g772(.A(KEYINPUT127), .B1(new_n1197), .B2(new_n961), .ZN(new_n1199));
  NOR2_X1   g773(.A1(new_n1198), .A2(new_n1199), .ZN(G308));
  NAND2_X1  g774(.A1(new_n1197), .A2(new_n961), .ZN(G225));
endmodule


