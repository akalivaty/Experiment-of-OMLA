//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0 0 0 1 1 0 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 1 1 1 1 1 0 1 1 1 1 1 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028;
  XNOR2_X1  g000(.A(KEYINPUT26), .B(G101), .ZN(new_n187));
  NOR2_X1   g001(.A1(G237), .A2(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G210), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT72), .B(KEYINPUT73), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  XOR2_X1   g008(.A(G116), .B(G119), .Z(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT2), .B(G113), .ZN(new_n196));
  XNOR2_X1  g010(.A(new_n195), .B(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT65), .B1(new_n198), .B2(G146), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT65), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(G146), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n199), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT1), .B1(new_n198), .B2(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G128), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n201), .A2(G143), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT1), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n208), .A2(new_n203), .A3(new_n209), .A4(G128), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT69), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n207), .A2(KEYINPUT69), .A3(new_n210), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(G134), .B(G137), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT11), .ZN(new_n217));
  INV_X1    g031(.A(G134), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n217), .B1(new_n218), .B2(G137), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(G137), .ZN(new_n220));
  INV_X1    g034(.A(G137), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(KEYINPUT11), .A3(G134), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n219), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G131), .ZN(new_n224));
  MUX2_X1   g038(.A(new_n216), .B(new_n223), .S(new_n224), .Z(new_n225));
  AOI21_X1  g039(.A(new_n197), .B1(new_n215), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(KEYINPUT64), .A2(KEYINPUT0), .ZN(new_n227));
  INV_X1    g041(.A(G128), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT64), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT0), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n230), .A2(new_n231), .A3(new_n228), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n204), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n208), .A2(new_n203), .A3(KEYINPUT0), .A4(G128), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT67), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n223), .B(G131), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n235), .A2(new_n240), .A3(new_n236), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n238), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(KEYINPUT28), .B1(new_n226), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT66), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n235), .A2(new_n245), .A3(new_n236), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n245), .B1(new_n235), .B2(new_n236), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n223), .B(new_n224), .ZN(new_n248));
  NOR3_X1   g062(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n225), .A2(new_n211), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n197), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT75), .ZN(new_n253));
  INV_X1    g067(.A(new_n247), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n235), .A2(new_n245), .A3(new_n236), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n239), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(new_n250), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT75), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(new_n258), .A3(new_n197), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n253), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT68), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n242), .A2(new_n261), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n238), .A2(KEYINPUT68), .A3(new_n239), .A4(new_n241), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(new_n226), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT70), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n262), .A2(new_n226), .A3(KEYINPUT70), .A4(new_n263), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n260), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT28), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n194), .B(new_n244), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n266), .A2(new_n267), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n215), .A2(new_n225), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n262), .A2(KEYINPUT30), .A3(new_n272), .A4(new_n263), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT30), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n257), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n273), .A2(new_n197), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n271), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n194), .ZN(new_n278));
  AOI21_X1  g092(.A(KEYINPUT29), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(G902), .B1(new_n270), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n262), .A2(new_n272), .A3(new_n263), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n197), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT76), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n271), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n266), .A2(KEYINPUT76), .A3(new_n267), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n283), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OAI211_X1 g101(.A(KEYINPUT29), .B(new_n244), .C1(new_n287), .C2(new_n269), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n280), .B1(new_n288), .B2(new_n278), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G472), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n271), .A2(new_n276), .A3(new_n194), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT31), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT74), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n252), .A2(KEYINPUT75), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n258), .B1(new_n257), .B2(new_n197), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n269), .B1(new_n271), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n278), .B1(new_n298), .B2(new_n243), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n271), .A2(new_n276), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT31), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(new_n301), .A3(new_n194), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n291), .A2(KEYINPUT74), .A3(KEYINPUT31), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n294), .A2(new_n299), .A3(new_n302), .A4(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT32), .ZN(new_n305));
  NOR2_X1   g119(.A1(G472), .A2(G902), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n305), .B1(new_n304), .B2(new_n306), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n290), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G953), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(G221), .A3(G234), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n311), .B(KEYINPUT22), .ZN(new_n312));
  AND2_X1   g126(.A1(new_n312), .A2(new_n221), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n312), .A2(new_n221), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT79), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT79), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n317), .B1(new_n313), .B2(new_n314), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G110), .ZN(new_n320));
  INV_X1    g134(.A(G119), .ZN(new_n321));
  OAI21_X1  g135(.A(KEYINPUT23), .B1(new_n321), .B2(G128), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT23), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(new_n228), .A3(G119), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n228), .A2(G119), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n320), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n328), .B(KEYINPUT77), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT78), .ZN(new_n330));
  INV_X1    g144(.A(G140), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G125), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n330), .B1(new_n332), .B2(KEYINPUT16), .ZN(new_n333));
  INV_X1    g147(.A(G125), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G140), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n332), .A2(new_n335), .A3(KEYINPUT16), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT16), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n337), .A2(new_n331), .A3(KEYINPUT78), .A4(G125), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n333), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n201), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n333), .A2(new_n336), .A3(G146), .A4(new_n338), .ZN(new_n341));
  XNOR2_X1  g155(.A(G119), .B(G128), .ZN(new_n342));
  XOR2_X1   g156(.A(KEYINPUT24), .B(G110), .Z(new_n343));
  AOI22_X1  g157(.A1(new_n340), .A2(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n325), .A2(new_n320), .A3(new_n327), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n345), .B1(new_n342), .B2(new_n343), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n332), .A2(new_n335), .A3(new_n201), .ZN(new_n347));
  AND2_X1   g161(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  AOI22_X1  g162(.A1(new_n329), .A2(new_n344), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  OR3_X1    g163(.A1(new_n319), .A2(new_n349), .A3(KEYINPUT80), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n315), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT80), .B1(new_n319), .B2(new_n349), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT25), .ZN(new_n355));
  INV_X1    g169(.A(G902), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(KEYINPUT25), .B1(new_n353), .B2(G902), .ZN(new_n358));
  INV_X1    g172(.A(G217), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n359), .B1(G234), .B2(new_n356), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n357), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n360), .A2(G902), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n363), .B(KEYINPUT81), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n353), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n366), .B(KEYINPUT82), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n362), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(G110), .B(G140), .ZN(new_n369));
  AND2_X1   g183(.A1(new_n310), .A2(G227), .ZN(new_n370));
  XOR2_X1   g184(.A(new_n369), .B(new_n370), .Z(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n235), .A2(new_n240), .A3(new_n236), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n240), .B1(new_n235), .B2(new_n236), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G104), .ZN(new_n376));
  OAI21_X1  g190(.A(KEYINPUT3), .B1(new_n376), .B2(G107), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT3), .ZN(new_n378));
  INV_X1    g192(.A(G107), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n379), .A3(G104), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n376), .A2(G107), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n377), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G101), .ZN(new_n383));
  OR2_X1    g197(.A1(new_n383), .A2(KEYINPUT4), .ZN(new_n384));
  INV_X1    g198(.A(G101), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n377), .A2(new_n380), .A3(new_n385), .A4(new_n381), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n383), .A2(KEYINPUT4), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT85), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n383), .A2(KEYINPUT85), .A3(KEYINPUT4), .A4(new_n386), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n375), .A2(new_n384), .A3(new_n389), .A4(new_n390), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n379), .A2(G104), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n376), .A2(G107), .ZN(new_n393));
  OAI21_X1  g207(.A(G101), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n386), .A2(new_n394), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n207), .A2(KEYINPUT69), .A3(new_n210), .ZN(new_n396));
  AOI21_X1  g210(.A(KEYINPUT69), .B1(new_n207), .B2(new_n210), .ZN(new_n397));
  OAI211_X1 g211(.A(KEYINPUT10), .B(new_n395), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n210), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n205), .A2(G128), .B1(new_n208), .B2(new_n203), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n395), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(KEYINPUT86), .B(KEYINPUT10), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n391), .A2(KEYINPUT87), .A3(new_n398), .A4(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n389), .A2(new_n384), .A3(new_n390), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n238), .A2(new_n241), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n398), .B(new_n403), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT87), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n248), .B1(new_n404), .B2(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n407), .A2(new_n239), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n372), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n401), .B1(new_n211), .B2(new_n395), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n239), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(KEYINPUT12), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n371), .B1(new_n407), .B2(new_n239), .ZN(new_n416));
  OR2_X1    g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n412), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G469), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n419), .A3(new_n356), .ZN(new_n420));
  NAND2_X1  g234(.A1(G469), .A2(G902), .ZN(new_n421));
  XOR2_X1   g235(.A(new_n371), .B(KEYINPUT84), .Z(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(new_n415), .B2(new_n411), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n423), .B(G469), .C1(new_n410), .C2(new_n416), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n420), .A2(new_n421), .A3(new_n424), .ZN(new_n425));
  XOR2_X1   g239(.A(KEYINPUT9), .B(G234), .Z(new_n426));
  XNOR2_X1  g240(.A(new_n426), .B(KEYINPUT83), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n356), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(G221), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(G475), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n340), .A2(new_n341), .ZN(new_n433));
  INV_X1    g247(.A(G237), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(new_n310), .A3(G214), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n198), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n188), .A2(G143), .A3(G214), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(KEYINPUT91), .B1(new_n438), .B2(G131), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT91), .ZN(new_n440));
  AOI211_X1 g254(.A(new_n440), .B(new_n224), .C1(new_n436), .C2(new_n437), .ZN(new_n441));
  OAI21_X1  g255(.A(KEYINPUT17), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(KEYINPUT90), .B1(new_n438), .B2(G131), .ZN(new_n443));
  AND4_X1   g257(.A1(G143), .A2(new_n434), .A3(new_n310), .A4(G214), .ZN(new_n444));
  AOI21_X1  g258(.A(G143), .B1(new_n188), .B2(G214), .ZN(new_n445));
  OAI21_X1  g259(.A(G131), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n440), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n438), .A2(KEYINPUT91), .A3(G131), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT90), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n436), .A2(new_n449), .A3(new_n224), .A4(new_n437), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n443), .A2(new_n447), .A3(new_n448), .A4(new_n450), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n433), .B(new_n442), .C1(new_n451), .C2(KEYINPUT17), .ZN(new_n452));
  XNOR2_X1  g266(.A(G113), .B(G122), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(new_n376), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n332), .A2(new_n335), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n455), .A2(KEYINPUT89), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT89), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n457), .B1(new_n332), .B2(new_n335), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n347), .B1(new_n459), .B2(new_n201), .ZN(new_n460));
  NAND2_X1  g274(.A1(KEYINPUT18), .A2(G131), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n438), .B(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n452), .A2(new_n454), .A3(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(KEYINPUT19), .B1(new_n456), .B2(new_n458), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n465), .B(new_n201), .C1(KEYINPUT19), .C2(new_n455), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n451), .A2(new_n466), .A3(new_n341), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n454), .B1(new_n467), .B2(new_n463), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n432), .B(new_n356), .C1(new_n464), .C2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT20), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n454), .B1(new_n452), .B2(new_n463), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n356), .B1(new_n464), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(G475), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n452), .A2(new_n454), .A3(new_n463), .ZN(new_n475));
  AND2_X1   g289(.A1(new_n467), .A2(new_n463), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n475), .B1(new_n476), .B2(new_n454), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n477), .A2(KEYINPUT20), .A3(new_n432), .A4(new_n356), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n471), .A2(new_n474), .A3(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G122), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(G116), .ZN(new_n482));
  INV_X1    g296(.A(G116), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(G122), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n482), .A2(new_n484), .A3(new_n379), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n379), .B1(new_n482), .B2(new_n484), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT92), .ZN(new_n487));
  NOR3_X1   g301(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n483), .A2(G122), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n481), .A2(G116), .ZN(new_n490));
  OAI21_X1  g304(.A(G107), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n482), .A2(new_n484), .A3(new_n379), .ZN(new_n492));
  AOI21_X1  g306(.A(KEYINPUT92), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n198), .A2(G128), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n228), .A2(G143), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n495), .A2(new_n496), .A3(new_n218), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(KEYINPUT95), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT13), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n499), .B1(new_n228), .B2(G143), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n496), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT93), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n218), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT94), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n198), .A2(KEYINPUT13), .A3(G128), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n500), .A2(new_n505), .A3(KEYINPUT93), .A4(new_n496), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n503), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n504), .B1(new_n503), .B2(new_n506), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n494), .B(new_n498), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n490), .A2(KEYINPUT14), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n482), .A2(new_n484), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n510), .B(G107), .C1(new_n511), .C2(KEYINPUT14), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n495), .A2(new_n496), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n513), .A2(G134), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n218), .B1(new_n495), .B2(new_n496), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n512), .B(new_n492), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n427), .A2(G217), .A3(new_n310), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n509), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n518), .B1(new_n509), .B2(new_n516), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n356), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT96), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(G478), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n524), .A2(KEYINPUT15), .ZN(new_n525));
  OAI211_X1 g339(.A(KEYINPUT96), .B(new_n356), .C1(new_n519), .C2(new_n520), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  OR2_X1    g341(.A1(new_n521), .A2(new_n525), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n310), .A2(G952), .ZN(new_n531));
  NAND2_X1  g345(.A1(G234), .A2(G237), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  XOR2_X1   g347(.A(KEYINPUT21), .B(G898), .Z(new_n534));
  NAND3_X1  g348(.A1(new_n532), .A2(G902), .A3(G953), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n480), .A2(new_n530), .A3(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(G214), .B1(G237), .B2(G902), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n389), .A2(new_n197), .A3(new_n384), .A4(new_n390), .ZN(new_n540));
  OR2_X1    g354(.A1(new_n195), .A2(new_n196), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT5), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n542), .A2(new_n321), .A3(G116), .ZN(new_n543));
  OAI211_X1 g357(.A(G113), .B(new_n543), .C1(new_n195), .C2(new_n542), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n395), .A2(new_n541), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g360(.A(G110), .B(G122), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n540), .A2(new_n547), .A3(new_n545), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(KEYINPUT6), .A3(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT88), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n207), .A2(new_n334), .A3(new_n210), .ZN(new_n553));
  INV_X1    g367(.A(new_n237), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n552), .B(new_n553), .C1(new_n554), .C2(new_n334), .ZN(new_n555));
  INV_X1    g369(.A(G224), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n556), .A2(G953), .ZN(new_n557));
  INV_X1    g371(.A(new_n553), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n334), .B1(new_n235), .B2(new_n236), .ZN(new_n559));
  OAI21_X1  g373(.A(KEYINPUT88), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n555), .A2(new_n557), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n557), .B1(new_n555), .B2(new_n560), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT6), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n546), .A2(new_n564), .A3(new_n548), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n551), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n544), .A2(new_n541), .ZN(new_n567));
  INV_X1    g381(.A(new_n395), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n545), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n547), .B(KEYINPUT8), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT7), .ZN(new_n573));
  OAI22_X1  g387(.A1(new_n558), .A2(new_n559), .B1(new_n573), .B2(new_n557), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n557), .A2(new_n573), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n553), .B(new_n575), .C1(new_n554), .C2(new_n334), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n550), .A2(new_n572), .A3(new_n574), .A4(new_n576), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n577), .A2(new_n356), .ZN(new_n578));
  OAI21_X1  g392(.A(G210), .B1(G237), .B2(G902), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n566), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n579), .B1(new_n566), .B2(new_n578), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n537), .A2(new_n539), .A3(new_n583), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n309), .A2(new_n368), .A3(new_n431), .A4(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(G101), .ZN(G3));
  NAND2_X1  g400(.A1(new_n304), .A2(new_n306), .ZN(new_n587));
  INV_X1    g401(.A(new_n303), .ZN(new_n588));
  AOI21_X1  g402(.A(KEYINPUT74), .B1(new_n291), .B2(KEYINPUT31), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n291), .A2(KEYINPUT31), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n244), .B1(new_n268), .B2(new_n269), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n591), .B1(new_n592), .B2(new_n278), .ZN(new_n593));
  AOI21_X1  g407(.A(G902), .B1(new_n590), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(G472), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n587), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n368), .ZN(new_n597));
  NOR3_X1   g411(.A1(new_n596), .A2(new_n597), .A3(new_n430), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n509), .A2(new_n516), .A3(new_n518), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT98), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n509), .A2(new_n516), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n517), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n509), .A2(KEYINPUT98), .A3(new_n516), .A4(new_n518), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n601), .A2(new_n603), .A3(KEYINPUT33), .A4(new_n604), .ZN(new_n605));
  XOR2_X1   g419(.A(KEYINPUT97), .B(KEYINPUT33), .Z(new_n606));
  OAI21_X1  g420(.A(new_n606), .B1(new_n519), .B2(new_n520), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT99), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n608), .A2(new_n609), .A3(G478), .A4(new_n356), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n523), .A2(new_n524), .A3(new_n526), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n605), .A2(G478), .A3(new_n356), .A4(new_n607), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(KEYINPUT99), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n479), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n566), .A2(new_n578), .ZN(new_n616));
  INV_X1    g430(.A(new_n579), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n580), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n619), .A2(new_n538), .A3(new_n536), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n615), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n598), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(G104), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n622), .B(new_n624), .ZN(G6));
  INV_X1    g439(.A(new_n620), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n530), .A2(new_n479), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n598), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT35), .B(G107), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G9));
  NAND2_X1  g446(.A1(new_n619), .A2(new_n538), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n349), .B(KEYINPUT101), .ZN(new_n634));
  INV_X1    g448(.A(new_n319), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n635), .A2(KEYINPUT36), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n634), .B(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n364), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n361), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n430), .A2(new_n633), .A3(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n537), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n595), .B1(new_n304), .B2(new_n356), .ZN(new_n644));
  INV_X1    g458(.A(new_n306), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n645), .B1(new_n590), .B2(new_n593), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n642), .A2(new_n643), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT37), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(new_n320), .ZN(G12));
  OAI21_X1  g464(.A(new_n533), .B1(G900), .B2(new_n535), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n530), .A2(new_n479), .A3(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n309), .A2(new_n642), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G128), .ZN(G30));
  NAND2_X1  g469(.A1(new_n587), .A2(KEYINPUT32), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n277), .A2(new_n194), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n266), .A2(KEYINPUT76), .A3(new_n267), .ZN(new_n659));
  AOI21_X1  g473(.A(KEYINPUT76), .B1(new_n266), .B2(new_n267), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n282), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OAI211_X1 g475(.A(new_n356), .B(new_n658), .C1(new_n661), .C2(new_n194), .ZN(new_n662));
  AOI22_X1  g476(.A1(new_n656), .A2(new_n657), .B1(G472), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n479), .A2(new_n529), .A3(new_n538), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n583), .A2(KEYINPUT38), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT38), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n619), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n651), .B(KEYINPUT39), .Z(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n425), .A2(new_n429), .A3(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT102), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n673), .A2(new_n674), .ZN(new_n676));
  OAI21_X1  g490(.A(KEYINPUT40), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n665), .A2(new_n670), .A3(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n676), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT40), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n673), .A2(new_n674), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n641), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n678), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(new_n198), .ZN(G45));
  NOR2_X1   g499(.A1(new_n615), .A2(new_n652), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n309), .A2(new_n642), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G146), .ZN(G48));
  AND2_X1   g502(.A1(new_n407), .A2(new_n408), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n407), .A2(new_n408), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n239), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n411), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n371), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n417), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n356), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(G469), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n696), .A2(new_n429), .A3(new_n420), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n309), .A2(new_n368), .A3(new_n621), .A4(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(KEYINPUT41), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G113), .ZN(G15));
  NAND4_X1  g515(.A1(new_n309), .A2(new_n368), .A3(new_n629), .A4(new_n698), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G116), .ZN(G18));
  NOR2_X1   g517(.A1(new_n697), .A2(new_n633), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n309), .A2(new_n643), .A3(new_n640), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G119), .ZN(G21));
  AOI21_X1  g520(.A(new_n243), .B1(new_n661), .B2(KEYINPUT28), .ZN(new_n707));
  OAI211_X1 g521(.A(new_n302), .B(new_n292), .C1(new_n707), .C2(new_n194), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n644), .B1(new_n306), .B2(new_n708), .ZN(new_n709));
  OR3_X1    g523(.A1(new_n664), .A2(new_n583), .A3(KEYINPUT103), .ZN(new_n710));
  OAI21_X1  g524(.A(KEYINPUT103), .B1(new_n664), .B2(new_n583), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n697), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n709), .A2(new_n368), .A3(new_n712), .A4(new_n536), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G122), .ZN(G24));
  NAND4_X1  g528(.A1(new_n709), .A2(new_n640), .A3(new_n686), .A4(new_n704), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G125), .ZN(G27));
  NAND2_X1  g530(.A1(new_n656), .A2(new_n657), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n597), .B1(new_n717), .B2(new_n290), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n581), .A2(new_n582), .A3(new_n539), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n686), .A2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n718), .A2(KEYINPUT42), .A3(new_n431), .A4(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n309), .A2(new_n721), .A3(new_n368), .A4(new_n431), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT42), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G131), .ZN(G33));
  INV_X1    g541(.A(new_n719), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n430), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n718), .A2(new_n653), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G134), .ZN(G36));
  INV_X1    g545(.A(new_n429), .ZN(new_n732));
  AOI211_X1 g546(.A(G469), .B(G902), .C1(new_n412), .C2(new_n417), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n423), .B1(new_n410), .B2(new_n416), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT45), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n423), .B(KEYINPUT45), .C1(new_n410), .C2(new_n416), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n736), .A2(G469), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n421), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT46), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n733), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n738), .A2(KEYINPUT46), .A3(new_n421), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n732), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n672), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT43), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT104), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n479), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n471), .A2(new_n474), .A3(new_n478), .A4(KEYINPUT104), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n745), .B1(new_n749), .B2(new_n614), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n614), .A2(new_n745), .A3(new_n480), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(KEYINPUT105), .B1(new_n596), .B2(new_n640), .ZN(new_n753));
  OAI211_X1 g567(.A(KEYINPUT105), .B(new_n640), .C1(new_n644), .C2(new_n646), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n752), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT44), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n744), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n752), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT105), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n760), .B1(new_n647), .B2(new_n641), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n759), .B1(new_n761), .B2(new_n754), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n728), .B1(new_n762), .B2(KEYINPUT44), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n758), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G137), .ZN(G39));
  INV_X1    g579(.A(KEYINPUT47), .ZN(new_n766));
  INV_X1    g580(.A(new_n742), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT46), .B1(new_n738), .B2(new_n421), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n767), .A2(new_n768), .A3(new_n733), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n766), .B1(new_n769), .B2(new_n732), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n743), .A2(KEYINPUT47), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n290), .B(new_n597), .C1(new_n307), .C2(new_n308), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n772), .A2(new_n721), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G140), .ZN(G42));
  NAND2_X1  g590(.A1(new_n663), .A2(new_n368), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n669), .A2(new_n614), .A3(new_n749), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n779), .A2(new_n732), .A3(new_n539), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n419), .B1(new_n418), .B2(new_n356), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n781), .A2(new_n733), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(KEYINPUT49), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n778), .A2(new_n780), .A3(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n785));
  AOI211_X1 g599(.A(new_n766), .B(new_n732), .C1(new_n741), .C2(new_n742), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n739), .A2(new_n740), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n787), .A2(new_n420), .A3(new_n742), .ZN(new_n788));
  AOI21_X1  g602(.A(KEYINPUT47), .B1(new_n788), .B2(new_n429), .ZN(new_n789));
  OAI21_X1  g603(.A(KEYINPUT110), .B1(new_n786), .B2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT110), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n770), .A2(new_n771), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n696), .A2(new_n420), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n429), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n790), .A2(new_n792), .A3(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n533), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n709), .A2(new_n368), .A3(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT109), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n798), .A2(new_n799), .A3(new_n719), .A4(new_n752), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n304), .A2(new_n356), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(G472), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n708), .A2(new_n306), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n802), .A2(new_n368), .A3(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n804), .A2(new_n797), .A3(new_n752), .ZN(new_n805));
  OAI21_X1  g619(.A(KEYINPUT109), .B1(new_n805), .B2(new_n728), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n796), .A2(new_n800), .A3(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT50), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT111), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n782), .A2(new_n429), .A3(new_n539), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n809), .B1(new_n810), .B2(new_n670), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n698), .A2(KEYINPUT111), .A3(new_n539), .A4(new_n669), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n808), .B1(new_n805), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n811), .A2(new_n812), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n798), .A2(KEYINPUT50), .A3(new_n752), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n696), .A2(new_n429), .A3(new_n420), .A4(new_n719), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(KEYINPUT112), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT112), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n782), .A2(new_n820), .A3(new_n429), .A4(new_n719), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n752), .A2(new_n819), .A3(new_n797), .A4(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT113), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n533), .B1(new_n818), .B2(KEYINPUT112), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n825), .A2(new_n752), .A3(KEYINPUT113), .A4(new_n821), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n827), .A2(new_n640), .A3(new_n709), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n819), .A2(new_n821), .A3(new_n797), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n778), .A2(new_n480), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n817), .A2(new_n828), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n785), .B1(new_n807), .B2(new_n832), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n817), .A2(new_n831), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n806), .B(new_n800), .C1(new_n772), .C2(new_n794), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n834), .A2(KEYINPUT51), .A3(new_n828), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n827), .A2(new_n718), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT48), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT48), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n827), .A2(new_n839), .A3(new_n718), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n615), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n830), .A2(new_n368), .A3(new_n842), .A4(new_n663), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n804), .A2(new_n797), .A3(new_n704), .A4(new_n752), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n843), .A2(new_n844), .A3(new_n531), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT114), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT114), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n843), .A2(new_n844), .A3(new_n847), .A4(new_n531), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n841), .A2(new_n849), .A3(KEYINPUT115), .ZN(new_n850));
  AOI21_X1  g664(.A(KEYINPUT115), .B1(new_n841), .B2(new_n849), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n833), .B(new_n836), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n853));
  AND4_X1   g667(.A1(new_n309), .A2(new_n530), .A3(new_n640), .A4(new_n729), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n479), .A2(new_n652), .ZN(new_n855));
  AOI21_X1  g669(.A(KEYINPUT107), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n309), .A2(new_n530), .A3(new_n640), .A4(new_n729), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT107), .ZN(new_n858));
  INV_X1    g672(.A(new_n855), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n726), .B1(new_n856), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n842), .A2(KEYINPUT106), .A3(new_n626), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT106), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n863), .B1(new_n615), .B2(new_n620), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n862), .A2(new_n628), .A3(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n597), .A2(new_n430), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n865), .A2(new_n647), .A3(new_n866), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n585), .A2(new_n867), .A3(new_n648), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n309), .A2(new_n368), .A3(new_n653), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n709), .A2(new_n640), .A3(new_n686), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(new_n729), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n699), .A2(new_n705), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n702), .A2(new_n713), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n868), .A2(new_n872), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n861), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n662), .A2(G472), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n877), .B1(new_n307), .B2(new_n308), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n710), .A2(new_n711), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT108), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n880), .B1(new_n640), .B2(new_n652), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n361), .A2(new_n639), .A3(KEYINPUT108), .A4(new_n651), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n430), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n878), .A2(new_n879), .A3(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n654), .A2(new_n715), .A3(new_n687), .A4(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT52), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n885), .B(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT53), .B1(new_n876), .B2(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n699), .A2(new_n702), .A3(new_n705), .A4(new_n713), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n585), .A2(new_n867), .A3(new_n648), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n309), .A2(new_n530), .A3(new_n640), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n892), .A2(KEYINPUT107), .A3(new_n729), .A4(new_n855), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n858), .B1(new_n857), .B2(new_n859), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n891), .A2(new_n895), .A3(new_n726), .A4(new_n872), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT53), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n715), .A2(new_n687), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n898), .A2(new_n886), .A3(new_n654), .A4(new_n884), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n885), .A2(KEYINPUT52), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n896), .A2(new_n897), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n853), .B1(new_n888), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n897), .B1(new_n896), .B2(new_n901), .ZN(new_n904));
  AND4_X1   g718(.A1(new_n872), .A2(new_n868), .A3(new_n874), .A4(new_n873), .ZN(new_n905));
  AOI22_X1  g719(.A1(new_n893), .A2(new_n894), .B1(new_n725), .B2(new_n722), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n887), .A2(new_n905), .A3(KEYINPUT53), .A4(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n904), .A2(KEYINPUT54), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n852), .B1(new_n903), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(G952), .A2(G953), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n784), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(KEYINPUT116), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT116), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n913), .B(new_n784), .C1(new_n909), .C2(new_n910), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n912), .A2(new_n914), .ZN(G75));
  AOI21_X1  g729(.A(new_n356), .B1(new_n904), .B2(new_n907), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(G210), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT56), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT117), .B1(new_n916), .B2(G210), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n551), .A2(new_n565), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(new_n563), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT55), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n919), .B1(new_n920), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n310), .A2(G952), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n917), .A2(KEYINPUT117), .A3(new_n918), .A4(new_n923), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n925), .A2(new_n927), .A3(new_n928), .ZN(G51));
  OR2_X1    g743(.A1(new_n738), .A2(KEYINPUT118), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n738), .A2(KEYINPUT118), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n916), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT119), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n421), .B(KEYINPUT57), .Z(new_n934));
  NAND3_X1  g748(.A1(new_n903), .A2(new_n908), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n418), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n926), .B1(new_n933), .B2(new_n936), .ZN(G54));
  NAND2_X1  g751(.A1(new_n904), .A2(new_n907), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n938), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n939));
  INV_X1    g753(.A(new_n477), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n927), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n939), .A2(new_n940), .ZN(new_n942));
  OR2_X1    g756(.A1(new_n942), .A2(KEYINPUT120), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(KEYINPUT120), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n941), .B1(new_n943), .B2(new_n944), .ZN(G60));
  NAND2_X1  g759(.A1(G478), .A2(G902), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT59), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n903), .A2(new_n908), .A3(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n608), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n948), .A2(new_n949), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n950), .A2(new_n951), .A3(new_n926), .ZN(G63));
  NAND2_X1  g766(.A1(G217), .A2(G902), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT60), .Z(new_n954));
  NAND3_X1  g768(.A1(new_n938), .A2(new_n638), .A3(new_n954), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n938), .A2(new_n954), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n927), .B(new_n955), .C1(new_n956), .C2(new_n354), .ZN(new_n957));
  AOI21_X1  g771(.A(KEYINPUT61), .B1(new_n955), .B2(KEYINPUT121), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n957), .B(new_n958), .ZN(G66));
  INV_X1    g773(.A(new_n534), .ZN(new_n960));
  OAI21_X1  g774(.A(G953), .B1(new_n960), .B2(new_n556), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n961), .B1(new_n891), .B2(G953), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n921), .B1(G898), .B2(new_n310), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(G69));
  AOI21_X1  g778(.A(new_n310), .B1(G227), .B2(G900), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT124), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n715), .A2(new_n654), .A3(new_n687), .ZN(new_n967));
  OAI21_X1  g781(.A(KEYINPUT62), .B1(new_n684), .B2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(new_n967), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT62), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n969), .B(new_n970), .C1(new_n683), .C2(new_n678), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  AOI211_X1 g786(.A(new_n720), .B(new_n773), .C1(new_n770), .C2(new_n771), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n973), .B1(new_n758), .B2(new_n763), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n675), .A2(new_n676), .A3(new_n728), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n975), .B(new_n718), .C1(new_n842), .C2(new_n627), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n972), .A2(KEYINPUT123), .A3(new_n974), .A4(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT123), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n974), .A2(new_n976), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n968), .A2(new_n971), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n978), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(G953), .B1(new_n977), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n273), .A2(new_n275), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n465), .B1(KEYINPUT19), .B2(new_n455), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT122), .Z(new_n985));
  XNOR2_X1  g799(.A(new_n983), .B(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n966), .B1(new_n982), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n719), .B1(new_n756), .B2(new_n757), .ZN(new_n989));
  INV_X1    g803(.A(new_n744), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n990), .B1(new_n762), .B2(KEYINPUT44), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n726), .B(new_n775), .C1(new_n989), .C2(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT125), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n990), .A2(new_n718), .A3(new_n994), .A4(new_n879), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n743), .A2(new_n309), .A3(new_n368), .A4(new_n672), .ZN(new_n996));
  INV_X1    g810(.A(new_n879), .ZN(new_n997));
  OAI21_X1  g811(.A(KEYINPUT125), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n967), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n993), .A2(KEYINPUT126), .A3(new_n730), .A4(new_n999), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n974), .A2(new_n726), .A3(new_n730), .A4(new_n999), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT126), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n1000), .A2(new_n1003), .A3(new_n310), .ZN(new_n1004));
  NAND2_X1  g818(.A1(G900), .A2(G953), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1004), .A2(new_n987), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n965), .B1(new_n988), .B2(new_n1007), .ZN(new_n1008));
  AND2_X1   g822(.A1(new_n977), .A2(new_n981), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n986), .B1(new_n1009), .B2(G953), .ZN(new_n1010));
  INV_X1    g824(.A(new_n965), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n1010), .A2(new_n966), .A3(new_n1011), .A4(new_n1006), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1008), .A2(new_n1012), .ZN(G72));
  NAND3_X1  g827(.A1(new_n1000), .A2(new_n1003), .A3(new_n891), .ZN(new_n1014));
  NAND2_X1  g828(.A1(G472), .A2(G902), .ZN(new_n1015));
  XOR2_X1   g829(.A(new_n1015), .B(KEYINPUT63), .Z(new_n1016));
  NAND2_X1  g830(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n1017), .A2(new_n300), .A3(new_n278), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n277), .A2(new_n278), .ZN(new_n1019));
  AOI22_X1  g833(.A1(new_n904), .A2(new_n907), .B1(new_n291), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n926), .B1(new_n1020), .B2(new_n1016), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n977), .A2(new_n981), .A3(new_n891), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1023), .A2(new_n1016), .ZN(new_n1024));
  INV_X1    g838(.A(new_n658), .ZN(new_n1025));
  AOI21_X1  g839(.A(KEYINPUT127), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g840(.A(KEYINPUT127), .ZN(new_n1027));
  AOI211_X1 g841(.A(new_n1027), .B(new_n658), .C1(new_n1023), .C2(new_n1016), .ZN(new_n1028));
  NOR3_X1   g842(.A1(new_n1022), .A2(new_n1026), .A3(new_n1028), .ZN(G57));
endmodule


