//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 1 0 1 0 0 0 0 1 0 0 1 0 0 1 0 0 1 1 0 0 0 0 1 1 0 1 0 1 1 1 0 0 0 0 1 1 0 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:54 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1279,
    new_n1280, new_n1281, new_n1282, new_n1283, new_n1284, new_n1285,
    new_n1286, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT0), .Z(new_n206));
  INV_X1    g0006(.A(G87), .ZN(new_n207));
  INV_X1    g0007(.A(G250), .ZN(new_n208));
  INV_X1    g0008(.A(G97), .ZN(new_n209));
  INV_X1    g0009(.A(G257), .ZN(new_n210));
  OAI22_X1  g0010(.A1(new_n207), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g0011(.A(new_n211), .B1(G68), .B2(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G107), .ZN(new_n213));
  INV_X1    g0013(.A(G264), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(G116), .B2(G270), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G50), .A2(G226), .ZN(new_n217));
  INV_X1    g0017(.A(G77), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n216), .B(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G58), .ZN(new_n221));
  INV_X1    g0021(.A(G232), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n203), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT64), .B(G20), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(G50), .B1(G58), .B2(G68), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT65), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n206), .B(new_n225), .C1(new_n228), .C2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G264), .ZN(new_n237));
  INV_X1    g0037(.A(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n235), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  OAI21_X1  g0048(.A(KEYINPUT66), .B1(new_n203), .B2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT66), .ZN(new_n250));
  NAND4_X1  g0050(.A1(new_n250), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n249), .A2(new_n227), .A3(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G1), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n252), .B1(new_n253), .B2(G20), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n253), .A2(G13), .A3(G20), .ZN(new_n255));
  OAI21_X1  g0055(.A(KEYINPUT12), .B1(new_n255), .B2(G68), .ZN(new_n256));
  OR3_X1    g0056(.A1(new_n255), .A2(KEYINPUT12), .A3(G68), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n254), .A2(G68), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G50), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n260), .B(KEYINPUT72), .ZN(new_n261));
  INV_X1    g0061(.A(G68), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G20), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n226), .A2(G33), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n261), .B(new_n263), .C1(new_n218), .C2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT11), .ZN(new_n266));
  AND3_X1   g0066(.A1(new_n265), .A2(new_n266), .A3(new_n252), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n266), .B1(new_n265), .B2(new_n252), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n258), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT73), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT73), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n271), .B(new_n258), .C1(new_n267), .C2(new_n268), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G169), .ZN(new_n274));
  INV_X1    g0074(.A(G41), .ZN(new_n275));
  INV_X1    g0075(.A(G45), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(new_n253), .A3(G274), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G226), .A2(G1698), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n280), .B1(new_n222), .B2(G1698), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT3), .B(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G33), .A2(G97), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AND2_X1   g0085(.A1(G1), .A2(G13), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n279), .B1(new_n285), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT13), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n253), .A2(new_n277), .B1(new_n286), .B2(new_n287), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G238), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n290), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n281), .A2(new_n282), .B1(G33), .B2(G97), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n293), .B(new_n278), .C1(new_n295), .C2(new_n288), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT13), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n274), .B1(new_n294), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT14), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n298), .B(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G179), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n294), .A2(new_n297), .A3(KEYINPUT71), .ZN(new_n302));
  OR3_X1    g0102(.A1(new_n296), .A2(KEYINPUT71), .A3(KEYINPUT13), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n273), .B1(new_n300), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n302), .A2(new_n303), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n269), .B1(new_n306), .B2(G190), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n294), .A2(new_n297), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(G200), .ZN(new_n309));
  OR2_X1    g0109(.A1(new_n309), .A2(KEYINPUT70), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(KEYINPUT70), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n307), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT8), .B(G58), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  AND2_X1   g0114(.A1(KEYINPUT64), .A2(G20), .ZN(new_n315));
  NOR2_X1   g0115(.A1(KEYINPUT64), .A2(G20), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n314), .A2(new_n259), .B1(new_n317), .B2(G77), .ZN(new_n318));
  XOR2_X1   g0118(.A(KEYINPUT15), .B(G87), .Z(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n318), .B1(new_n264), .B2(new_n320), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n321), .A2(new_n252), .B1(new_n254), .B2(G77), .ZN(new_n322));
  INV_X1    g0122(.A(new_n255), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n218), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(G238), .A2(G1698), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n282), .B(new_n326), .C1(new_n222), .C2(G1698), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n327), .B(new_n289), .C1(G107), .C2(new_n282), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n292), .A2(G244), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n328), .A2(new_n278), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G200), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(KEYINPUT69), .B1(new_n325), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT69), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n331), .A2(new_n322), .A3(new_n334), .A4(new_n324), .ZN(new_n335));
  INV_X1    g0135(.A(G190), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n333), .B(new_n335), .C1(new_n336), .C2(new_n330), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n305), .A2(new_n312), .A3(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n255), .A2(G50), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n254), .A2(G50), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G20), .ZN(new_n342));
  NOR2_X1   g0142(.A1(G58), .A2(G68), .ZN(new_n343));
  INV_X1    g0143(.A(G50), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n345), .B1(G150), .B2(new_n259), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT67), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n347), .A2(new_n221), .A3(KEYINPUT8), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(new_n314), .B2(new_n347), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n346), .B1(new_n349), .B2(new_n264), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n252), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT68), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n350), .A2(KEYINPUT68), .A3(new_n252), .ZN(new_n354));
  AOI211_X1 g0154(.A(new_n339), .B(new_n341), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G1698), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(G222), .ZN(new_n357));
  INV_X1    g0157(.A(G223), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n282), .B(new_n357), .C1(new_n358), .C2(new_n356), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n359), .B(new_n289), .C1(G77), .C2(new_n282), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n292), .A2(G226), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n360), .A2(new_n278), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n274), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(G179), .B2(new_n362), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n355), .A2(new_n364), .ZN(new_n365));
  OR2_X1    g0165(.A1(new_n330), .A2(G179), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n330), .A2(new_n274), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n325), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n362), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n355), .A2(KEYINPUT9), .B1(G190), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT10), .ZN(new_n372));
  INV_X1    g0172(.A(new_n339), .ZN(new_n373));
  INV_X1    g0173(.A(new_n354), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT68), .B1(new_n350), .B2(new_n252), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n373), .B(new_n340), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT9), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n362), .A2(G200), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n371), .A2(new_n372), .A3(new_n378), .A4(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n378), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n370), .A2(G190), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n379), .B(new_n382), .C1(new_n376), .C2(new_n377), .ZN(new_n383));
  OAI21_X1  g0183(.A(KEYINPUT10), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  AOI211_X1 g0184(.A(new_n365), .B(new_n369), .C1(new_n380), .C2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT74), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT3), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n386), .B1(new_n387), .B2(G33), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n248), .A2(KEYINPUT74), .A3(KEYINPUT3), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n387), .A2(G33), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT7), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n392), .A2(new_n393), .A3(new_n226), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n248), .A2(KEYINPUT3), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n395), .B1(new_n388), .B2(new_n389), .ZN(new_n396));
  OAI21_X1  g0196(.A(KEYINPUT7), .B1(new_n396), .B2(G20), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n394), .A2(G68), .A3(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n221), .A2(new_n262), .ZN(new_n399));
  OAI21_X1  g0199(.A(G20), .B1(new_n399), .B2(new_n343), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n259), .A2(G159), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n398), .A2(KEYINPUT16), .A3(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT16), .ZN(new_n405));
  OAI21_X1  g0205(.A(KEYINPUT75), .B1(new_n387), .B2(G33), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT75), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n407), .A2(new_n248), .A3(KEYINPUT3), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n406), .A2(new_n408), .A3(new_n391), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n409), .A2(KEYINPUT7), .A3(new_n226), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n393), .B1(new_n282), .B2(G20), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n262), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n405), .B1(new_n412), .B2(new_n402), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n404), .A2(new_n413), .A3(new_n252), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n349), .A2(new_n255), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n254), .B2(new_n349), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G226), .A2(G1698), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n358), .B2(G1698), .ZN(new_n419));
  AND3_X1   g0219(.A1(new_n248), .A2(KEYINPUT74), .A3(KEYINPUT3), .ZN(new_n420));
  AOI21_X1  g0220(.A(KEYINPUT74), .B1(new_n248), .B2(KEYINPUT3), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n391), .B(new_n419), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(G33), .A2(G87), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n288), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n253), .B1(G41), .B2(G45), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n288), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n278), .B1(new_n426), .B2(new_n222), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT76), .ZN(new_n428));
  NOR4_X1   g0228(.A1(new_n424), .A2(new_n427), .A3(new_n428), .A4(G179), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n274), .B1(new_n424), .B2(new_n427), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT76), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n422), .A2(new_n423), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n427), .B1(new_n432), .B2(new_n289), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n301), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n429), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n417), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT18), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT18), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n417), .A2(new_n438), .A3(new_n435), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT17), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT77), .ZN(new_n441));
  NOR4_X1   g0241(.A1(new_n424), .A2(new_n427), .A3(new_n441), .A4(G190), .ZN(new_n442));
  OAI21_X1  g0242(.A(KEYINPUT77), .B1(new_n433), .B2(G200), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n433), .A2(new_n336), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n440), .B1(new_n417), .B2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n442), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n279), .B1(new_n292), .B2(G232), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n396), .A2(new_n419), .B1(G33), .B2(G87), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n448), .B1(new_n449), .B2(new_n288), .ZN(new_n450));
  INV_X1    g0250(.A(G200), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n441), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n450), .A2(G190), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n447), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n454), .A2(KEYINPUT17), .A3(new_n414), .A4(new_n416), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n437), .A2(new_n439), .A3(new_n446), .A4(new_n455), .ZN(new_n456));
  OR2_X1    g0256(.A1(new_n456), .A2(KEYINPUT78), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(KEYINPUT78), .ZN(new_n458));
  AND4_X1   g0258(.A1(new_n338), .A2(new_n385), .A3(new_n457), .A4(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n255), .A2(G97), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n255), .B1(G1), .B2(new_n248), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n252), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G97), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n410), .A2(new_n411), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G107), .ZN(new_n467));
  INV_X1    g0267(.A(new_n259), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(new_n218), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT6), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n209), .A2(new_n213), .ZN(new_n472));
  NOR2_X1   g0272(.A1(G97), .A2(G107), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n213), .A2(KEYINPUT6), .A3(G97), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n226), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n467), .A2(new_n470), .A3(new_n477), .ZN(new_n478));
  AOI211_X1 g0278(.A(new_n461), .B(new_n465), .C1(new_n478), .C2(new_n252), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n219), .A2(G1698), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n390), .A2(new_n391), .A3(new_n480), .ZN(new_n481));
  XOR2_X1   g0281(.A(KEYINPUT79), .B(KEYINPUT4), .Z(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT80), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n480), .A2(KEYINPUT4), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n486), .B1(new_n208), .B2(new_n356), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n487), .A2(new_n282), .B1(G33), .B2(G283), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n481), .A2(KEYINPUT80), .A3(new_n482), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n485), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n289), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n276), .A2(G1), .ZN(new_n492));
  AND2_X1   g0292(.A1(KEYINPUT5), .A2(G41), .ZN(new_n493));
  NOR2_X1   g0293(.A1(KEYINPUT5), .A2(G41), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(G274), .ZN(new_n496));
  OR2_X1    g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n495), .A2(new_n288), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n497), .B1(new_n498), .B2(new_n210), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(G200), .B1(new_n491), .B2(new_n500), .ZN(new_n501));
  AOI211_X1 g0301(.A(G190), .B(new_n499), .C1(new_n490), .C2(new_n289), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n479), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n491), .A2(new_n301), .A3(new_n500), .ZN(new_n504));
  INV_X1    g0304(.A(new_n461), .ZN(new_n505));
  AOI211_X1 g0305(.A(new_n469), .B(new_n476), .C1(new_n466), .C2(G107), .ZN(new_n506));
  INV_X1    g0306(.A(new_n252), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n505), .B(new_n464), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n499), .B1(new_n490), .B2(new_n289), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n504), .B(new_n508), .C1(G169), .C2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT82), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT81), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n512), .B1(new_n253), .B2(G45), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n496), .B1(new_n208), .B2(KEYINPUT81), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n513), .A2(G250), .B1(new_n514), .B2(new_n492), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n511), .B1(new_n515), .B2(new_n289), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n492), .ZN(new_n517));
  OAI211_X1 g0317(.A(KEYINPUT81), .B(G250), .C1(new_n276), .C2(G1), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n519), .A2(KEYINPUT82), .A3(new_n288), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(G238), .A2(G1698), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n522), .B1(new_n219), .B2(G1698), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n396), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(G116), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT83), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT83), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G116), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(new_n528), .A3(G33), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n288), .B1(new_n524), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(G200), .B1(new_n521), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n319), .A2(new_n255), .ZN(new_n532));
  NAND3_X1  g0332(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n315), .B2(new_n316), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT85), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n207), .A2(new_n209), .A3(new_n213), .ZN(new_n537));
  OAI211_X1 g0337(.A(KEYINPUT85), .B(new_n533), .C1(new_n315), .C2(new_n316), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n226), .A2(G33), .A3(G97), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT19), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n396), .A2(G68), .A3(new_n226), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n539), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n532), .B1(new_n544), .B2(new_n252), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n463), .A2(G87), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n531), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT86), .ZN(new_n548));
  XNOR2_X1  g0348(.A(KEYINPUT83), .B(G116), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n396), .A2(new_n523), .B1(G33), .B2(new_n549), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n516), .B(new_n520), .C1(new_n288), .C2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n548), .B1(new_n551), .B2(new_n336), .ZN(new_n552));
  NOR3_X1   g0352(.A1(new_n515), .A2(new_n511), .A3(new_n289), .ZN(new_n553));
  AOI21_X1  g0353(.A(KEYINPUT82), .B1(new_n519), .B2(new_n288), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n530), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n555), .A2(new_n556), .A3(KEYINPUT86), .A4(G190), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n547), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n463), .A2(new_n319), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n545), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(KEYINPUT84), .B1(new_n551), .B2(G179), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n551), .A2(new_n274), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT84), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n555), .A2(new_n556), .A3(new_n564), .A4(new_n301), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n561), .A2(new_n562), .A3(new_n563), .A4(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n503), .A2(new_n510), .A3(new_n559), .A4(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT24), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT23), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n529), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n342), .ZN(new_n571));
  NAND2_X1  g0371(.A1(KEYINPUT23), .A2(G107), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT22), .ZN(new_n573));
  OAI21_X1  g0373(.A(G87), .B1(new_n315), .B2(new_n316), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n248), .A2(KEYINPUT3), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n391), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n573), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n317), .A2(new_n569), .A3(new_n213), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n571), .A2(new_n572), .A3(new_n577), .A4(new_n578), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n396), .A2(KEYINPUT22), .A3(G87), .A4(new_n226), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n568), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  AND3_X1   g0382(.A1(new_n577), .A2(new_n572), .A3(new_n578), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n583), .A2(KEYINPUT24), .A3(new_n571), .A4(new_n580), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n582), .A2(new_n584), .A3(new_n252), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n323), .A2(KEYINPUT25), .A3(new_n213), .ZN(new_n586));
  XOR2_X1   g0386(.A(new_n586), .B(KEYINPUT88), .Z(new_n587));
  AOI21_X1  g0387(.A(KEYINPUT25), .B1(new_n323), .B2(new_n213), .ZN(new_n588));
  XNOR2_X1  g0388(.A(new_n588), .B(KEYINPUT89), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n587), .A2(new_n589), .B1(G107), .B2(new_n463), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n585), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n495), .A2(G264), .A3(new_n288), .ZN(new_n592));
  NAND2_X1  g0392(.A1(G257), .A2(G1698), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(new_n208), .B2(G1698), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n396), .A2(new_n594), .B1(G33), .B2(G294), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n497), .B(new_n592), .C1(new_n595), .C2(new_n288), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT90), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n390), .A2(new_n391), .A3(new_n594), .ZN(new_n598));
  NAND2_X1  g0398(.A1(G33), .A2(G294), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n289), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT90), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n601), .A2(new_n602), .A3(new_n497), .A4(new_n592), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n274), .B1(new_n597), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n596), .A2(new_n301), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n591), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n597), .A2(new_n603), .A3(new_n336), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n596), .A2(new_n451), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n609), .A2(new_n590), .A3(new_n585), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n210), .A2(G1698), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n390), .A2(new_n391), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT87), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n214), .A2(new_n356), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n396), .A2(new_n615), .B1(G303), .B2(new_n576), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT87), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n396), .A2(new_n617), .A3(new_n612), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n614), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n289), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n498), .A2(new_n238), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n620), .A2(G190), .A3(new_n497), .A4(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n527), .A2(G116), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n525), .A2(KEYINPUT83), .ZN(new_n625));
  OAI21_X1  g0425(.A(G20), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n248), .A2(G97), .ZN(new_n627));
  NAND2_X1  g0427(.A1(G33), .A2(G283), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n627), .B(new_n628), .C1(new_n315), .C2(new_n316), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n252), .A2(new_n626), .A3(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT20), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n252), .A2(new_n626), .A3(KEYINPUT20), .A4(new_n629), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n549), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n463), .A2(G116), .B1(new_n323), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n497), .ZN(new_n639));
  AOI211_X1 g0439(.A(new_n639), .B(new_n621), .C1(new_n619), .C2(new_n289), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n623), .B(new_n638), .C1(new_n640), .C2(new_n451), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT21), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n637), .A2(G169), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n642), .B1(new_n640), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n640), .A2(G179), .A3(new_n637), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n620), .A2(new_n497), .A3(new_n622), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n646), .A2(KEYINPUT21), .A3(G169), .A4(new_n637), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n641), .A2(new_n644), .A3(new_n645), .A4(new_n647), .ZN(new_n648));
  NOR4_X1   g0448(.A1(new_n460), .A2(new_n567), .A3(new_n611), .A4(new_n648), .ZN(G372));
  INV_X1    g0449(.A(new_n365), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n380), .A2(new_n384), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n446), .A2(new_n455), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n312), .A2(new_n369), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n652), .B1(new_n653), .B2(new_n305), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n437), .A2(new_n439), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n651), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(G169), .B1(new_n555), .B2(new_n556), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT91), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n657), .A2(new_n658), .B1(new_n545), .B2(new_n560), .ZN(new_n659));
  INV_X1    g0459(.A(new_n551), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n563), .A2(KEYINPUT91), .B1(new_n660), .B2(new_n301), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n659), .A2(new_n661), .B1(new_n547), .B2(new_n558), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n663), .A2(new_n503), .A3(new_n510), .A4(new_n610), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n644), .A2(new_n645), .A3(new_n647), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n597), .A2(new_n603), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(G169), .ZN(new_n667));
  INV_X1    g0467(.A(new_n605), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n667), .A2(new_n668), .B1(new_n590), .B2(new_n585), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n662), .B1(new_n664), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n510), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT26), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(new_n663), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n559), .A2(new_n566), .ZN(new_n675));
  OAI21_X1  g0475(.A(KEYINPUT26), .B1(new_n675), .B2(new_n510), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n671), .A2(new_n677), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n650), .B(new_n656), .C1(new_n460), .C2(new_n678), .ZN(G369));
  INV_X1    g0479(.A(G13), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n317), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  OR3_X1    g0482(.A1(new_n682), .A2(KEYINPUT27), .A3(G1), .ZN(new_n683));
  OAI21_X1  g0483(.A(KEYINPUT27), .B1(new_n682), .B2(G1), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G213), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(G343), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(new_n638), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n665), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n648), .A2(new_n689), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(G330), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT92), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n606), .B2(new_n688), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n669), .A2(KEYINPUT92), .A3(new_n687), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n591), .A2(new_n687), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n699), .B1(new_n611), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n695), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT93), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n665), .A2(new_n688), .ZN(new_n704));
  AOI22_X1  g0504(.A1(new_n701), .A2(new_n704), .B1(new_n669), .B2(new_n688), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n703), .A2(new_n705), .ZN(G399));
  INV_X1    g0506(.A(new_n204), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(G41), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(G1), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n537), .A2(G116), .ZN(new_n711));
  INV_X1    g0511(.A(new_n230), .ZN(new_n712));
  OAI22_X1  g0512(.A1(new_n710), .A2(new_n711), .B1(new_n712), .B2(new_n709), .ZN(new_n713));
  XOR2_X1   g0513(.A(KEYINPUT94), .B(KEYINPUT28), .Z(new_n714));
  XNOR2_X1  g0514(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n611), .A2(new_n648), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n503), .A2(new_n510), .ZN(new_n717));
  INV_X1    g0517(.A(new_n675), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n716), .A2(new_n717), .A3(new_n718), .A4(new_n688), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n640), .A2(G179), .A3(new_n660), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n601), .A2(new_n592), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n509), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(KEYINPUT95), .B2(KEYINPUT30), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT96), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n509), .A2(G179), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n551), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n646), .A2(new_n596), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n725), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(KEYINPUT95), .A2(KEYINPUT30), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(new_n720), .B2(new_n722), .ZN(new_n731));
  INV_X1    g0531(.A(new_n728), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n732), .A2(KEYINPUT96), .A3(new_n726), .A4(new_n551), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n724), .A2(new_n729), .A3(new_n731), .A4(new_n733), .ZN(new_n734));
  AOI22_X1  g0534(.A1(new_n719), .A2(KEYINPUT31), .B1(new_n687), .B2(new_n734), .ZN(new_n735));
  OAI211_X1 g0535(.A(new_n724), .B(new_n731), .C1(new_n727), .C2(new_n728), .ZN(new_n736));
  AND3_X1   g0536(.A1(new_n736), .A2(KEYINPUT31), .A3(new_n687), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n738), .A2(G330), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n718), .A2(new_n673), .A3(new_n672), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n662), .A2(new_n559), .ZN(new_n741));
  OAI21_X1  g0541(.A(KEYINPUT26), .B1(new_n741), .B2(new_n510), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n688), .B1(new_n671), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(KEYINPUT29), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT29), .ZN(new_n746));
  OAI211_X1 g0546(.A(new_n746), .B(new_n688), .C1(new_n671), .C2(new_n677), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n739), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n715), .B1(new_n749), .B2(G1), .ZN(G364));
  AOI21_X1  g0550(.A(new_n227), .B1(G20), .B2(new_n274), .ZN(new_n751));
  OAI21_X1  g0551(.A(KEYINPUT98), .B1(new_n226), .B2(new_n301), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT98), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n317), .A2(new_n753), .A3(G179), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n755), .A2(G190), .A3(new_n451), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n755), .A2(new_n336), .A3(new_n451), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n221), .A2(new_n756), .B1(new_n757), .B2(new_n218), .ZN(new_n758));
  XOR2_X1   g0558(.A(new_n758), .B(KEYINPUT99), .Z(new_n759));
  NAND3_X1  g0559(.A1(new_n755), .A2(G190), .A3(G200), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n759), .B1(new_n344), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT100), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G179), .A2(G200), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G190), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n317), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n209), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n451), .A2(G179), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n317), .A2(new_n336), .A3(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n213), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n755), .A2(new_n336), .A3(G200), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n770), .B1(new_n772), .B2(G68), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n768), .A2(G20), .A3(G190), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G87), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n317), .A2(new_n336), .A3(new_n763), .ZN(new_n777));
  XOR2_X1   g0577(.A(KEYINPUT101), .B(G159), .Z(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT32), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n773), .A2(new_n776), .A3(new_n781), .ZN(new_n782));
  NOR4_X1   g0582(.A1(new_n762), .A2(new_n576), .A3(new_n767), .A4(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(KEYINPUT33), .B(G317), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n772), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n760), .ZN(new_n786));
  XOR2_X1   g0586(.A(KEYINPUT102), .B(G326), .Z(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n282), .B1(new_n775), .B2(G303), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n765), .A2(G294), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n785), .A2(new_n788), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G311), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n757), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G322), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n756), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G283), .ZN(new_n796));
  INV_X1    g0596(.A(G329), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n796), .A2(new_n769), .B1(new_n777), .B2(new_n797), .ZN(new_n798));
  NOR4_X1   g0598(.A1(new_n791), .A2(new_n793), .A3(new_n795), .A4(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n751), .B1(new_n783), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(G13), .A2(G33), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(G20), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n693), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n681), .A2(G45), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n710), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n282), .A2(G355), .A3(new_n204), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n243), .A2(new_n276), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n396), .A2(new_n707), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(new_n712), .B2(G45), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n809), .B1(G116), .B2(new_n204), .C1(new_n810), .C2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n803), .A2(new_n751), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n808), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n815), .B(KEYINPUT97), .Z(new_n816));
  NAND3_X1  g0616(.A1(new_n800), .A2(new_n804), .A3(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n695), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n693), .A2(new_n694), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n818), .A2(new_n819), .A3(new_n808), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n817), .A2(new_n820), .ZN(G396));
  NAND2_X1  g0621(.A1(new_n738), .A2(G330), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n368), .A2(new_n687), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n687), .A2(new_n325), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n337), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n823), .B1(new_n825), .B2(new_n368), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n688), .B(new_n826), .C1(new_n671), .C2(new_n677), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n678), .A2(new_n687), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n826), .B(KEYINPUT103), .Z(new_n829));
  OAI211_X1 g0629(.A(new_n822), .B(new_n827), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n827), .B1(new_n829), .B2(new_n828), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n739), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n830), .A2(new_n832), .A3(new_n808), .ZN(new_n833));
  INV_X1    g0633(.A(G303), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n796), .A2(new_n771), .B1(new_n760), .B2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n757), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n549), .ZN(new_n837));
  INV_X1    g0637(.A(new_n777), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n767), .B1(G311), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n769), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(G87), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n837), .A2(new_n576), .A3(new_n839), .A4(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n756), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n835), .B(new_n842), .C1(G294), .C2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n213), .B2(new_n774), .ZN(new_n845));
  AOI22_X1  g0645(.A1(G143), .A2(new_n843), .B1(new_n836), .B2(new_n778), .ZN(new_n846));
  INV_X1    g0646(.A(G137), .ZN(new_n847));
  INV_X1    g0647(.A(G150), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n846), .B1(new_n847), .B2(new_n760), .C1(new_n848), .C2(new_n771), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT34), .Z(new_n850));
  AOI22_X1  g0650(.A1(new_n840), .A2(G68), .B1(G58), .B2(new_n765), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n392), .B1(G50), .B2(new_n775), .ZN(new_n852));
  INV_X1    g0652(.A(G132), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n851), .B(new_n852), .C1(new_n853), .C2(new_n777), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n845), .B1(new_n850), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n751), .A2(new_n801), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n855), .A2(new_n751), .B1(new_n218), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n857), .B1(new_n802), .B2(new_n826), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n807), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n833), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT104), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n860), .B(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(G384));
  INV_X1    g0663(.A(KEYINPUT38), .ZN(new_n864));
  INV_X1    g0664(.A(new_n685), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n404), .A2(new_n252), .ZN(new_n866));
  AOI21_X1  g0666(.A(KEYINPUT16), .B1(new_n398), .B2(new_n403), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n416), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT106), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OAI211_X1 g0670(.A(KEYINPUT106), .B(new_n416), .C1(new_n866), .C2(new_n867), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AND3_X1   g0672(.A1(new_n456), .A2(new_n865), .A3(new_n872), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n430), .A2(KEYINPUT76), .B1(new_n433), .B2(new_n301), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n685), .B1(new_n874), .B2(new_n429), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n417), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n454), .A2(new_n414), .A3(new_n416), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT37), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n870), .A2(new_n871), .A3(new_n875), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n877), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n879), .B1(new_n881), .B2(KEYINPUT37), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n864), .B1(new_n873), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n456), .A2(new_n865), .A3(new_n872), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n878), .B1(new_n880), .B2(new_n877), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n884), .B(KEYINPUT38), .C1(new_n885), .C2(new_n879), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n273), .A2(new_n687), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n305), .A2(new_n312), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n888), .B1(new_n305), .B2(new_n312), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT105), .ZN(new_n893));
  INV_X1    g0693(.A(new_n823), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n827), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n893), .B1(new_n827), .B2(new_n894), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n887), .B(new_n892), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  OR2_X1    g0698(.A1(new_n305), .A2(new_n687), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n456), .A2(new_n417), .A3(new_n865), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n878), .B1(new_n876), .B2(new_n877), .ZN(new_n901));
  OAI21_X1  g0701(.A(KEYINPUT107), .B1(new_n879), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n876), .A2(new_n877), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(KEYINPUT37), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT107), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n900), .A2(new_n902), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT108), .B1(new_n908), .B2(new_n864), .ZN(new_n909));
  OAI21_X1  g0709(.A(KEYINPUT39), .B1(new_n887), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n908), .A2(new_n864), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT39), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n911), .A2(KEYINPUT108), .A3(new_n912), .A4(new_n886), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n899), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n865), .B1(new_n437), .B2(new_n439), .ZN(new_n915));
  NOR3_X1   g0715(.A1(new_n898), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n656), .A2(new_n650), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n917), .B1(new_n748), .B2(new_n459), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n916), .B(new_n918), .Z(new_n919));
  OAI21_X1  g0719(.A(new_n826), .B1(new_n889), .B2(new_n890), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n734), .A2(new_n687), .ZN(new_n921));
  NOR4_X1   g0721(.A1(new_n567), .A2(new_n611), .A3(new_n648), .A4(new_n687), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT31), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n734), .A2(KEYINPUT31), .A3(new_n687), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n920), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT40), .B1(new_n926), .B2(new_n887), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT40), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(new_n911), .B2(new_n886), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n926), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT109), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n929), .A2(new_n926), .A3(KEYINPUT109), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n927), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n924), .A2(new_n925), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n934), .A2(new_n459), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n926), .A2(new_n887), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n928), .ZN(new_n938));
  AND3_X1   g0738(.A1(new_n929), .A2(KEYINPUT109), .A3(new_n926), .ZN(new_n939));
  AOI21_X1  g0739(.A(KEYINPUT109), .B1(new_n929), .B2(new_n926), .ZN(new_n940));
  OAI211_X1 g0740(.A(G330), .B(new_n938), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n694), .B1(new_n924), .B2(new_n925), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n459), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n936), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n919), .B(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n253), .B2(new_n681), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n474), .A2(new_n475), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n525), .B1(new_n948), .B2(KEYINPUT35), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n949), .B(new_n228), .C1(KEYINPUT35), .C2(new_n948), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT36), .ZN(new_n951));
  NOR3_X1   g0751(.A1(new_n712), .A2(new_n218), .A3(new_n399), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n262), .A2(G50), .ZN(new_n953));
  OAI211_X1 g0753(.A(G1), .B(new_n680), .C1(new_n952), .C2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n947), .A2(new_n951), .A3(new_n954), .ZN(G367));
  XNOR2_X1  g0755(.A(new_n708), .B(KEYINPUT41), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT113), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n702), .B(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n701), .B(new_n704), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n818), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n749), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n717), .B1(new_n479), .B2(new_n688), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n672), .A2(new_n687), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n965), .A2(KEYINPUT111), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT111), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(new_n963), .B2(new_n964), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n705), .ZN(new_n970));
  OAI21_X1  g0770(.A(KEYINPUT45), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n965), .B(KEYINPUT111), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT45), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n972), .A2(new_n973), .A3(new_n705), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n703), .ZN(new_n976));
  OAI211_X1 g0776(.A(KEYINPUT112), .B(KEYINPUT44), .C1(new_n972), .C2(new_n705), .ZN(new_n977));
  XOR2_X1   g0777(.A(KEYINPUT112), .B(KEYINPUT44), .Z(new_n978));
  NAND3_X1  g0778(.A1(new_n969), .A2(new_n970), .A3(new_n978), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n975), .A2(new_n976), .A3(new_n977), .A4(new_n979), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n977), .A2(new_n971), .A3(new_n974), .A4(new_n979), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n703), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n962), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n749), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n956), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n806), .A2(new_n253), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n701), .A2(new_n704), .ZN(new_n988));
  OAI21_X1  g0788(.A(KEYINPUT42), .B1(new_n969), .B2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT42), .ZN(new_n990));
  INV_X1    g0790(.A(new_n988), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n972), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  AND2_X1   g0792(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT43), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n688), .B1(new_n546), .B2(new_n545), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n662), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n663), .B2(new_n995), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT110), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n669), .B1(new_n966), .B2(new_n968), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n687), .B1(new_n999), .B2(new_n510), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n993), .A2(new_n994), .A3(new_n998), .A4(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n998), .A2(new_n994), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n998), .A2(new_n994), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n989), .A2(new_n992), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n1003), .B(new_n1004), .C1(new_n1005), .C2(new_n1000), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n703), .A2(new_n969), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1002), .A2(new_n1008), .A3(new_n1006), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n987), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n811), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n814), .B1(new_n204), .B2(new_n320), .C1(new_n239), .C2(new_n1015), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n786), .A2(G143), .B1(G137), .B2(new_n838), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n576), .B1(new_n775), .B2(G58), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1017), .B(new_n1018), .C1(new_n848), .C2(new_n756), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n771), .A2(new_n779), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n757), .A2(new_n344), .B1(new_n262), .B2(new_n766), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n769), .A2(new_n218), .ZN(new_n1022));
  NOR4_X1   g0822(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .A4(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n392), .B1(new_n757), .B2(new_n796), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT46), .ZN(new_n1025));
  NOR3_X1   g0825(.A1(new_n774), .A2(new_n1025), .A3(new_n525), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n840), .A2(G97), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n213), .B2(new_n766), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1026), .B(new_n1028), .C1(G317), .C2(new_n838), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1025), .B1(new_n635), .B2(new_n774), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1029), .B(new_n1030), .C1(new_n834), .C2(new_n756), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n1024), .B(new_n1031), .C1(G311), .C2(new_n786), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n772), .A2(G294), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1023), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT47), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n751), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n807), .B(new_n1016), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n803), .B2(new_n998), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT114), .Z(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1014), .A2(new_n1040), .ZN(G387));
  INV_X1    g0841(.A(G317), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n834), .A2(new_n757), .B1(new_n756), .B2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT116), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n792), .B2(new_n771), .C1(new_n794), .C2(new_n760), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1045), .A2(KEYINPUT48), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(KEYINPUT48), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n1046), .A2(new_n1047), .B1(G294), .B2(new_n775), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n765), .A2(G283), .ZN(new_n1049));
  AND3_X1   g0849(.A1(new_n1048), .A2(KEYINPUT49), .A3(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(KEYINPUT49), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n392), .B1(new_n769), .B2(new_n635), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(new_n838), .B2(new_n787), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n766), .A2(new_n320), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n836), .B2(G68), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1057), .B(new_n1027), .C1(new_n344), .C2(new_n756), .ZN(new_n1058));
  INV_X1    g0858(.A(G159), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n396), .B1(new_n771), .B2(new_n349), .C1(new_n1059), .C2(new_n760), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n774), .A2(new_n218), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n777), .A2(new_n848), .ZN(new_n1062));
  NOR4_X1   g0862(.A1(new_n1058), .A2(new_n1060), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1055), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n751), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT117), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n314), .A2(new_n344), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT50), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n262), .A2(new_n218), .ZN(new_n1070));
  NOR4_X1   g0870(.A1(new_n1069), .A2(G45), .A3(new_n1070), .A4(new_n711), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n811), .B1(new_n235), .B2(new_n276), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n711), .A2(new_n204), .A3(new_n282), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1071), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n204), .A2(G107), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n814), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1066), .A2(new_n1067), .A3(new_n807), .A4(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1063), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n807), .B(new_n1076), .C1(new_n1078), .C2(new_n1036), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(KEYINPUT117), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n803), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1077), .B(new_n1080), .C1(new_n701), .C2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n958), .A2(new_n960), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1083), .A2(new_n986), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT115), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n984), .A2(new_n1083), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n962), .A2(new_n708), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1082), .A2(new_n1085), .A3(new_n1087), .ZN(G393));
  NAND2_X1  g0888(.A1(new_n969), .A2(new_n803), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n792), .A2(new_n756), .B1(new_n760), .B2(new_n1042), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT52), .Z(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(G322), .B2(new_n838), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n775), .A2(G283), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n772), .A2(G303), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n836), .A2(G294), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n766), .A2(new_n635), .ZN(new_n1097));
  NOR4_X1   g0897(.A1(new_n1096), .A2(new_n282), .A3(new_n770), .A4(new_n1097), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n848), .A2(new_n760), .B1(new_n756), .B2(new_n1059), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT51), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n396), .B1(new_n262), .B2(new_n774), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(G77), .B2(new_n765), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n836), .A2(new_n314), .B1(G143), .B2(new_n838), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1100), .A2(new_n841), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(G50), .B2(new_n772), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n751), .B1(new_n1098), .B2(new_n1105), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n814), .B1(new_n209), .B2(new_n204), .C1(new_n246), .C2(new_n1015), .ZN(new_n1107));
  AND4_X1   g0907(.A1(new_n807), .A2(new_n1089), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n980), .A2(new_n982), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n986), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1108), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n980), .A2(new_n962), .A3(new_n982), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n708), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1111), .B1(new_n1113), .B2(new_n983), .ZN(G390));
  NAND2_X1  g0914(.A1(new_n911), .A2(new_n886), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n899), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n825), .A2(new_n368), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n688), .B(new_n1117), .C1(new_n671), .C2(new_n743), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n891), .B1(new_n1118), .B2(new_n894), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g0920(.A(G330), .B(new_n826), .C1(new_n735), .C2(new_n737), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1121), .A2(new_n891), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n895), .A2(new_n896), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n899), .B1(new_n1123), .B2(new_n891), .ZN(new_n1124));
  AND2_X1   g0924(.A1(new_n910), .A2(new_n913), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n1120), .B(new_n1122), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n942), .A2(new_n826), .A3(new_n892), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n827), .A2(new_n894), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(KEYINPUT105), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n827), .A2(new_n893), .A3(new_n894), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n891), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n899), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n910), .B(new_n913), .C1(new_n1131), .C2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1120), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1127), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1126), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n1110), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1125), .A2(new_n801), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n843), .A2(G132), .B1(G125), .B2(new_n838), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n576), .B1(new_n840), .B2(G50), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(KEYINPUT120), .ZN(new_n1141));
  INV_X1    g0941(.A(G128), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1139), .B(new_n1141), .C1(new_n1142), .C2(new_n760), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n775), .A2(G150), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT53), .ZN(new_n1145));
  XOR2_X1   g0945(.A(KEYINPUT54), .B(G143), .Z(new_n1146));
  AND2_X1   g0946(.A1(new_n836), .A2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1140), .A2(KEYINPUT120), .ZN(new_n1148));
  NOR4_X1   g0948(.A1(new_n1143), .A2(new_n1145), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n1149), .B1(new_n847), .B2(new_n771), .C1(new_n1059), .C2(new_n766), .ZN(new_n1150));
  XOR2_X1   g0950(.A(new_n1150), .B(KEYINPUT121), .Z(new_n1151));
  AOI22_X1  g0951(.A1(G97), .A2(new_n836), .B1(new_n843), .B2(G116), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n772), .A2(G107), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1152), .A2(new_n776), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(G294), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n262), .A2(new_n769), .B1(new_n777), .B2(new_n1155), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n1156), .A2(KEYINPUT122), .B1(G77), .B2(new_n765), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1157), .B1(KEYINPUT122), .B2(new_n1156), .C1(new_n796), .C2(new_n760), .ZN(new_n1158));
  NOR3_X1   g0958(.A1(new_n1154), .A2(new_n282), .A3(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n751), .B1(new_n1151), .B2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n808), .B1(new_n349), .B2(new_n856), .ZN(new_n1161));
  XOR2_X1   g0961(.A(new_n1161), .B(KEYINPUT119), .Z(new_n1162));
  NAND3_X1  g0962(.A1(new_n1138), .A2(new_n1160), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n918), .A2(new_n943), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT118), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1164), .B(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1122), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n1118), .A2(new_n894), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n942), .A2(new_n829), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n891), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1167), .A2(new_n1168), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1121), .A2(new_n891), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n1172), .A2(new_n1127), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1171), .B1(new_n1173), .B2(new_n1123), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1166), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1133), .A2(new_n1134), .A3(new_n1167), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1120), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1176), .B1(new_n1177), .B2(new_n1127), .ZN(new_n1178));
  AND2_X1   g0978(.A1(new_n1175), .A2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n708), .B1(new_n1175), .B2(new_n1178), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1137), .B(new_n1163), .C1(new_n1179), .C2(new_n1180), .ZN(G378));
  NAND2_X1  g0981(.A1(new_n651), .A2(new_n650), .ZN(new_n1182));
  XOR2_X1   g0982(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1182), .B(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n355), .A2(new_n685), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1185), .B(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n941), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n932), .A2(new_n933), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1190), .A2(G330), .A3(new_n938), .A4(new_n1187), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n1189), .A2(new_n1191), .A3(new_n916), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n916), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1192), .A2(new_n1193), .A3(new_n986), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1188), .A2(new_n802), .ZN(new_n1195));
  NOR3_X1   g0995(.A1(new_n751), .A2(G50), .A3(new_n801), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n396), .A2(G41), .ZN(new_n1197));
  AOI211_X1 g0997(.A(G50), .B(new_n1197), .C1(new_n248), .C2(new_n275), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n843), .A2(G128), .B1(new_n775), .B2(new_n1146), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1199), .B1(new_n853), .B2(new_n771), .C1(new_n847), .C2(new_n757), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(G150), .B2(new_n765), .ZN(new_n1201));
  INV_X1    g1001(.A(G125), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1201), .B1(new_n1202), .B2(new_n760), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT59), .Z(new_n1204));
  INV_X1    g1004(.A(G124), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n248), .B(new_n275), .C1(new_n777), .C2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(new_n840), .B2(new_n778), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1198), .B1(new_n1204), .B2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1061), .B1(new_n843), .B2(G107), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1209), .B1(new_n221), .B2(new_n769), .C1(new_n796), .C2(new_n777), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n766), .A2(new_n262), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1197), .B1(new_n757), .B2(new_n320), .C1(new_n209), .C2(new_n771), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n760), .A2(new_n525), .ZN(new_n1213));
  NOR4_X1   g1013(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  XOR2_X1   g1014(.A(new_n1214), .B(KEYINPUT58), .Z(new_n1215));
  AOI21_X1  g1015(.A(new_n1036), .B1(new_n1208), .B2(new_n1215), .ZN(new_n1216));
  NOR4_X1   g1016(.A1(new_n1195), .A2(new_n808), .A3(new_n1196), .A4(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(KEYINPUT123), .B1(new_n1194), .B2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT123), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1217), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n916), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1187), .B1(new_n934), .B2(G330), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n941), .A2(new_n1188), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1221), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1189), .A2(new_n1191), .A3(new_n916), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1219), .B(new_n1220), .C1(new_n1226), .C2(new_n986), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1218), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT57), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1164), .B(KEYINPUT118), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n1136), .B2(new_n1174), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1229), .B1(new_n1231), .B2(new_n1226), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1123), .B1(new_n1127), .B2(new_n1172), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1122), .B1(new_n891), .B2(new_n1169), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1234), .B1(new_n1235), .B2(new_n1168), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1166), .B1(new_n1178), .B2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1233), .A2(new_n1237), .A3(KEYINPUT57), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1232), .A2(new_n708), .A3(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1228), .A2(new_n1239), .ZN(G375));
  NAND2_X1  g1040(.A1(new_n1230), .A2(new_n1236), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1241), .A2(new_n1175), .A3(new_n956), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n757), .A2(new_n848), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n760), .A2(new_n853), .B1(new_n1142), .B2(new_n777), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n1243), .B(new_n1244), .C1(G137), .C2(new_n843), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n772), .A2(new_n1146), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n765), .A2(G50), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n396), .B1(new_n1059), .B2(new_n774), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(G58), .B2(new_n840), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .A4(new_n1249), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n756), .A2(new_n796), .B1(new_n834), .B2(new_n777), .ZN(new_n1251));
  OR3_X1    g1051(.A1(new_n1022), .A2(KEYINPUT124), .A3(new_n282), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n1251), .B(new_n1253), .C1(new_n549), .C2(new_n772), .ZN(new_n1254));
  OAI21_X1  g1054(.A(KEYINPUT124), .B1(new_n1022), .B2(new_n282), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n836), .A2(G107), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1056), .B1(new_n786), .B2(G294), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .A4(new_n1257), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n774), .A2(new_n209), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1250), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n751), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n807), .B(new_n1261), .C1(new_n892), .C2(new_n802), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1262), .B1(new_n262), .B2(new_n856), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(new_n1174), .B2(new_n1110), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1242), .A2(new_n1264), .ZN(G381));
  INV_X1    g1065(.A(G378), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT125), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n1228), .A2(new_n1239), .A3(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1267), .B1(new_n1228), .B2(new_n1239), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n862), .B(new_n1266), .C1(new_n1268), .C2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(G390), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1014), .A2(new_n1271), .A3(new_n1040), .ZN(new_n1272));
  INV_X1    g1072(.A(G396), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1082), .A2(new_n1273), .A3(new_n1085), .A4(new_n1087), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1272), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NOR3_X1   g1076(.A1(new_n1270), .A2(G381), .A3(new_n1276), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(new_n1277), .B(KEYINPUT126), .ZN(G407));
  INV_X1    g1078(.A(G213), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1280), .A2(G378), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1279), .B1(new_n1281), .B2(new_n686), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1270), .A2(G381), .ZN(new_n1283));
  AOI21_X1  g1083(.A(KEYINPUT126), .B1(new_n1283), .B2(new_n1275), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT126), .ZN(new_n1285));
  NOR4_X1   g1085(.A1(new_n1270), .A2(new_n1285), .A3(G381), .A4(new_n1276), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1282), .B1(new_n1284), .B2(new_n1286), .ZN(G409));
  NAND2_X1  g1087(.A1(G393), .A2(G396), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n1274), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1012), .B1(new_n985), .B2(new_n986), .ZN(new_n1290));
  OAI21_X1  g1090(.A(G390), .B1(new_n1290), .B2(new_n1039), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1272), .A2(new_n1289), .A3(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1289), .B1(new_n1272), .B2(new_n1291), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT61), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1279), .A2(G343), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1228), .A2(new_n1239), .A3(G378), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1233), .A2(new_n1237), .A3(new_n956), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1298), .B(new_n1220), .C1(new_n986), .C2(new_n1226), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n1266), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1296), .B1(new_n1297), .B2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT60), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1302), .B1(new_n1166), .B2(new_n1174), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1230), .A2(KEYINPUT60), .A3(new_n1236), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1303), .A2(new_n1304), .A3(new_n708), .A4(new_n1175), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1264), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(G384), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1305), .A2(new_n862), .A3(new_n1264), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1296), .A2(G2897), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1307), .A2(G2897), .A3(new_n1296), .A4(new_n1308), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  OAI211_X1 g1113(.A(new_n1294), .B(new_n1295), .C1(new_n1301), .C2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1308), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n862), .B1(new_n1305), .B2(new_n1264), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  AOI211_X1 g1118(.A(new_n1296), .B(new_n1318), .C1(new_n1297), .C2(new_n1300), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT127), .ZN(new_n1320));
  OAI21_X1  g1120(.A(KEYINPUT63), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1301), .A2(new_n1309), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT63), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1322), .A2(KEYINPUT127), .A3(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1315), .A2(new_n1321), .A3(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT62), .ZN(new_n1326));
  AND3_X1   g1126(.A1(new_n1301), .A2(new_n1326), .A3(new_n1309), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1295), .B1(new_n1301), .B2(new_n1313), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1326), .B1(new_n1301), .B2(new_n1309), .ZN(new_n1329));
  NOR3_X1   g1129(.A1(new_n1327), .A2(new_n1328), .A3(new_n1329), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1325), .B1(new_n1330), .B2(new_n1294), .ZN(G405));
  NAND2_X1  g1131(.A1(G375), .A2(new_n1266), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(new_n1297), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1333), .A2(new_n1318), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1332), .A2(new_n1297), .A3(new_n1309), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  XNOR2_X1  g1136(.A(new_n1336), .B(new_n1294), .ZN(G402));
endmodule


