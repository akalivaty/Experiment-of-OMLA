

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U553 ( .A(n525), .B(n524), .ZN(n553) );
  INV_X1 U554 ( .A(KEYINPUT26), .ZN(n684) );
  INV_X1 U555 ( .A(KEYINPUT64), .ZN(n689) );
  OR2_X1 U556 ( .A1(n697), .A2(n696), .ZN(n694) );
  NOR2_X1 U557 ( .A1(n745), .A2(n744), .ZN(n767) );
  NOR2_X1 U558 ( .A1(n682), .A2(G1384), .ZN(n785) );
  NAND2_X1 U559 ( .A1(G160), .A2(G40), .ZN(n786) );
  NOR2_X2 U560 ( .A1(G2104), .A2(n520), .ZN(n859) );
  NOR2_X2 U561 ( .A1(n530), .A2(n529), .ZN(G160) );
  INV_X1 U562 ( .A(G2105), .ZN(n520) );
  AND2_X1 U563 ( .A1(n520), .A2(G2104), .ZN(n863) );
  NAND2_X1 U564 ( .A1(G101), .A2(n863), .ZN(n519) );
  XOR2_X1 U565 ( .A(KEYINPUT23), .B(n519), .Z(n523) );
  NAND2_X1 U566 ( .A1(G125), .A2(n859), .ZN(n521) );
  XOR2_X1 U567 ( .A(KEYINPUT65), .B(n521), .Z(n522) );
  NAND2_X1 U568 ( .A1(n523), .A2(n522), .ZN(n530) );
  XNOR2_X1 U569 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n525) );
  NOR2_X1 U570 ( .A1(G2105), .A2(G2104), .ZN(n524) );
  NAND2_X1 U571 ( .A1(G137), .A2(n553), .ZN(n528) );
  AND2_X1 U572 ( .A1(G2104), .A2(G2105), .ZN(n526) );
  XNOR2_X2 U573 ( .A(KEYINPUT66), .B(n526), .ZN(n860) );
  NAND2_X1 U574 ( .A1(G113), .A2(n860), .ZN(n527) );
  NAND2_X1 U575 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U576 ( .A1(G543), .A2(G651), .ZN(n643) );
  NAND2_X1 U577 ( .A1(G85), .A2(n643), .ZN(n532) );
  XOR2_X1 U578 ( .A(KEYINPUT0), .B(G543), .Z(n638) );
  INV_X1 U579 ( .A(G651), .ZN(n533) );
  NOR2_X1 U580 ( .A1(n638), .A2(n533), .ZN(n646) );
  NAND2_X1 U581 ( .A1(G72), .A2(n646), .ZN(n531) );
  NAND2_X1 U582 ( .A1(n532), .A2(n531), .ZN(n538) );
  NOR2_X1 U583 ( .A1(G543), .A2(n533), .ZN(n534) );
  XOR2_X1 U584 ( .A(KEYINPUT1), .B(n534), .Z(n642) );
  NAND2_X1 U585 ( .A1(G60), .A2(n642), .ZN(n536) );
  NOR2_X2 U586 ( .A1(n638), .A2(G651), .ZN(n650) );
  NAND2_X1 U587 ( .A1(G47), .A2(n650), .ZN(n535) );
  NAND2_X1 U588 ( .A1(n536), .A2(n535), .ZN(n537) );
  OR2_X1 U589 ( .A1(n538), .A2(n537), .ZN(G290) );
  AND2_X1 U590 ( .A1(G452), .A2(G94), .ZN(G173) );
  XOR2_X1 U591 ( .A(KEYINPUT18), .B(KEYINPUT75), .Z(n540) );
  NAND2_X1 U592 ( .A1(G123), .A2(n859), .ZN(n539) );
  XNOR2_X1 U593 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U594 ( .A(KEYINPUT74), .B(n541), .ZN(n543) );
  NAND2_X1 U595 ( .A1(n553), .A2(G135), .ZN(n542) );
  NAND2_X1 U596 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U597 ( .A(KEYINPUT76), .B(n544), .ZN(n548) );
  NAND2_X1 U598 ( .A1(G99), .A2(n863), .ZN(n546) );
  NAND2_X1 U599 ( .A1(G111), .A2(n860), .ZN(n545) );
  NAND2_X1 U600 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U601 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U602 ( .A(KEYINPUT77), .B(n549), .ZN(n1000) );
  XNOR2_X1 U603 ( .A(G2096), .B(n1000), .ZN(n550) );
  OR2_X1 U604 ( .A1(G2100), .A2(n550), .ZN(G156) );
  NAND2_X1 U605 ( .A1(G126), .A2(n859), .ZN(n552) );
  NAND2_X1 U606 ( .A1(G102), .A2(n863), .ZN(n551) );
  NAND2_X1 U607 ( .A1(n552), .A2(n551), .ZN(n560) );
  NAND2_X1 U608 ( .A1(n553), .A2(G138), .ZN(n555) );
  INV_X1 U609 ( .A(KEYINPUT87), .ZN(n554) );
  XNOR2_X1 U610 ( .A(n555), .B(n554), .ZN(n558) );
  NAND2_X1 U611 ( .A1(n860), .A2(G114), .ZN(n556) );
  XNOR2_X1 U612 ( .A(n556), .B(KEYINPUT86), .ZN(n557) );
  NAND2_X1 U613 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X1 U614 ( .A1(n560), .A2(n559), .ZN(n682) );
  BUF_X1 U615 ( .A(n682), .Z(G164) );
  INV_X1 U616 ( .A(G57), .ZN(G237) );
  INV_X1 U617 ( .A(G132), .ZN(G219) );
  INV_X1 U618 ( .A(G82), .ZN(G220) );
  NAND2_X1 U619 ( .A1(G88), .A2(n643), .ZN(n562) );
  NAND2_X1 U620 ( .A1(G75), .A2(n646), .ZN(n561) );
  NAND2_X1 U621 ( .A1(n562), .A2(n561), .ZN(n566) );
  NAND2_X1 U622 ( .A1(G62), .A2(n642), .ZN(n564) );
  NAND2_X1 U623 ( .A1(G50), .A2(n650), .ZN(n563) );
  NAND2_X1 U624 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U625 ( .A1(n566), .A2(n565), .ZN(G166) );
  NAND2_X1 U626 ( .A1(G64), .A2(n642), .ZN(n568) );
  NAND2_X1 U627 ( .A1(G52), .A2(n650), .ZN(n567) );
  NAND2_X1 U628 ( .A1(n568), .A2(n567), .ZN(n573) );
  NAND2_X1 U629 ( .A1(G90), .A2(n643), .ZN(n570) );
  NAND2_X1 U630 ( .A1(G77), .A2(n646), .ZN(n569) );
  NAND2_X1 U631 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U632 ( .A(KEYINPUT9), .B(n571), .Z(n572) );
  NOR2_X1 U633 ( .A1(n573), .A2(n572), .ZN(G171) );
  NAND2_X1 U634 ( .A1(G7), .A2(G661), .ZN(n574) );
  XNOR2_X1 U635 ( .A(n574), .B(KEYINPUT68), .ZN(n575) );
  XNOR2_X1 U636 ( .A(KEYINPUT10), .B(n575), .ZN(G223) );
  INV_X1 U637 ( .A(G223), .ZN(n825) );
  NAND2_X1 U638 ( .A1(n825), .A2(G567), .ZN(n576) );
  XOR2_X1 U639 ( .A(KEYINPUT11), .B(n576), .Z(G234) );
  NAND2_X1 U640 ( .A1(G56), .A2(n642), .ZN(n577) );
  XOR2_X1 U641 ( .A(KEYINPUT14), .B(n577), .Z(n583) );
  NAND2_X1 U642 ( .A1(n643), .A2(G81), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(KEYINPUT12), .ZN(n580) );
  NAND2_X1 U644 ( .A1(G68), .A2(n646), .ZN(n579) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U646 ( .A(KEYINPUT13), .B(n581), .Z(n582) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n585) );
  NAND2_X1 U648 ( .A1(n650), .A2(G43), .ZN(n584) );
  NAND2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n923) );
  INV_X1 U650 ( .A(G860), .ZN(n616) );
  OR2_X1 U651 ( .A1(n923), .A2(n616), .ZN(G153) );
  INV_X1 U652 ( .A(G171), .ZN(G301) );
  NAND2_X1 U653 ( .A1(G868), .A2(G301), .ZN(n595) );
  NAND2_X1 U654 ( .A1(G79), .A2(n646), .ZN(n592) );
  NAND2_X1 U655 ( .A1(G66), .A2(n642), .ZN(n587) );
  NAND2_X1 U656 ( .A1(G92), .A2(n643), .ZN(n586) );
  NAND2_X1 U657 ( .A1(n587), .A2(n586), .ZN(n590) );
  NAND2_X1 U658 ( .A1(G54), .A2(n650), .ZN(n588) );
  XNOR2_X1 U659 ( .A(KEYINPUT69), .B(n588), .ZN(n589) );
  NOR2_X1 U660 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U661 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U662 ( .A(n593), .B(KEYINPUT15), .ZN(n918) );
  INV_X1 U663 ( .A(n918), .ZN(n697) );
  INV_X1 U664 ( .A(G868), .ZN(n653) );
  NAND2_X1 U665 ( .A1(n697), .A2(n653), .ZN(n594) );
  NAND2_X1 U666 ( .A1(n595), .A2(n594), .ZN(G284) );
  NAND2_X1 U667 ( .A1(n643), .A2(G89), .ZN(n596) );
  XNOR2_X1 U668 ( .A(n596), .B(KEYINPUT4), .ZN(n598) );
  NAND2_X1 U669 ( .A1(G76), .A2(n646), .ZN(n597) );
  NAND2_X1 U670 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U671 ( .A(n599), .B(KEYINPUT5), .ZN(n604) );
  NAND2_X1 U672 ( .A1(G63), .A2(n642), .ZN(n601) );
  NAND2_X1 U673 ( .A1(G51), .A2(n650), .ZN(n600) );
  NAND2_X1 U674 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U675 ( .A(KEYINPUT6), .B(n602), .Z(n603) );
  NAND2_X1 U676 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U677 ( .A(n605), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U678 ( .A(G168), .B(KEYINPUT8), .Z(n606) );
  XNOR2_X1 U679 ( .A(KEYINPUT70), .B(n606), .ZN(G286) );
  NAND2_X1 U680 ( .A1(G65), .A2(n642), .ZN(n608) );
  NAND2_X1 U681 ( .A1(G53), .A2(n650), .ZN(n607) );
  NAND2_X1 U682 ( .A1(n608), .A2(n607), .ZN(n612) );
  NAND2_X1 U683 ( .A1(G91), .A2(n643), .ZN(n610) );
  NAND2_X1 U684 ( .A1(G78), .A2(n646), .ZN(n609) );
  NAND2_X1 U685 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U686 ( .A1(n612), .A2(n611), .ZN(n928) );
  INV_X1 U687 ( .A(n928), .ZN(G299) );
  XNOR2_X1 U688 ( .A(KEYINPUT71), .B(G868), .ZN(n613) );
  NOR2_X1 U689 ( .A1(G286), .A2(n613), .ZN(n615) );
  NOR2_X1 U690 ( .A1(G868), .A2(G299), .ZN(n614) );
  NOR2_X1 U691 ( .A1(n615), .A2(n614), .ZN(G297) );
  NAND2_X1 U692 ( .A1(n616), .A2(G559), .ZN(n617) );
  NAND2_X1 U693 ( .A1(n617), .A2(n918), .ZN(n618) );
  XNOR2_X1 U694 ( .A(n618), .B(KEYINPUT72), .ZN(n619) );
  XNOR2_X1 U695 ( .A(KEYINPUT16), .B(n619), .ZN(G148) );
  NOR2_X1 U696 ( .A1(G868), .A2(n923), .ZN(n620) );
  XOR2_X1 U697 ( .A(KEYINPUT73), .B(n620), .Z(n623) );
  NAND2_X1 U698 ( .A1(G868), .A2(n918), .ZN(n621) );
  NOR2_X1 U699 ( .A1(G559), .A2(n621), .ZN(n622) );
  NOR2_X1 U700 ( .A1(n623), .A2(n622), .ZN(G282) );
  NAND2_X1 U701 ( .A1(G80), .A2(n646), .ZN(n624) );
  XNOR2_X1 U702 ( .A(n624), .B(KEYINPUT78), .ZN(n631) );
  NAND2_X1 U703 ( .A1(G93), .A2(n643), .ZN(n626) );
  NAND2_X1 U704 ( .A1(G55), .A2(n650), .ZN(n625) );
  NAND2_X1 U705 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U706 ( .A1(G67), .A2(n642), .ZN(n627) );
  XNOR2_X1 U707 ( .A(KEYINPUT79), .B(n627), .ZN(n628) );
  NOR2_X1 U708 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U709 ( .A1(n631), .A2(n630), .ZN(n661) );
  NAND2_X1 U710 ( .A1(n918), .A2(G559), .ZN(n664) );
  XNOR2_X1 U711 ( .A(n923), .B(n664), .ZN(n632) );
  NOR2_X1 U712 ( .A1(G860), .A2(n632), .ZN(n633) );
  XOR2_X1 U713 ( .A(n661), .B(n633), .Z(G145) );
  NAND2_X1 U714 ( .A1(G49), .A2(n650), .ZN(n635) );
  NAND2_X1 U715 ( .A1(G74), .A2(G651), .ZN(n634) );
  NAND2_X1 U716 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U717 ( .A1(n642), .A2(n636), .ZN(n637) );
  XNOR2_X1 U718 ( .A(KEYINPUT80), .B(n637), .ZN(n641) );
  NAND2_X1 U719 ( .A1(n638), .A2(G87), .ZN(n639) );
  XOR2_X1 U720 ( .A(KEYINPUT81), .B(n639), .Z(n640) );
  NAND2_X1 U721 ( .A1(n641), .A2(n640), .ZN(G288) );
  NAND2_X1 U722 ( .A1(G61), .A2(n642), .ZN(n645) );
  NAND2_X1 U723 ( .A1(G86), .A2(n643), .ZN(n644) );
  NAND2_X1 U724 ( .A1(n645), .A2(n644), .ZN(n649) );
  NAND2_X1 U725 ( .A1(n646), .A2(G73), .ZN(n647) );
  XOR2_X1 U726 ( .A(KEYINPUT2), .B(n647), .Z(n648) );
  NOR2_X1 U727 ( .A1(n649), .A2(n648), .ZN(n652) );
  NAND2_X1 U728 ( .A1(n650), .A2(G48), .ZN(n651) );
  NAND2_X1 U729 ( .A1(n652), .A2(n651), .ZN(G305) );
  NAND2_X1 U730 ( .A1(n653), .A2(n661), .ZN(n654) );
  XNOR2_X1 U731 ( .A(n654), .B(KEYINPUT84), .ZN(n667) );
  XNOR2_X1 U732 ( .A(KEYINPUT82), .B(KEYINPUT19), .ZN(n656) );
  XNOR2_X1 U733 ( .A(G290), .B(KEYINPUT83), .ZN(n655) );
  XNOR2_X1 U734 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U735 ( .A(G288), .B(n657), .ZN(n659) );
  XNOR2_X1 U736 ( .A(n928), .B(G166), .ZN(n658) );
  XNOR2_X1 U737 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U738 ( .A(n660), .B(G305), .ZN(n662) );
  XNOR2_X1 U739 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U740 ( .A(n663), .B(n923), .ZN(n905) );
  XNOR2_X1 U741 ( .A(n905), .B(n664), .ZN(n665) );
  NAND2_X1 U742 ( .A1(G868), .A2(n665), .ZN(n666) );
  NAND2_X1 U743 ( .A1(n667), .A2(n666), .ZN(n668) );
  XOR2_X1 U744 ( .A(KEYINPUT85), .B(n668), .Z(G295) );
  NAND2_X1 U745 ( .A1(G2078), .A2(G2084), .ZN(n669) );
  XOR2_X1 U746 ( .A(KEYINPUT20), .B(n669), .Z(n670) );
  NAND2_X1 U747 ( .A1(G2090), .A2(n670), .ZN(n671) );
  XNOR2_X1 U748 ( .A(KEYINPUT21), .B(n671), .ZN(n672) );
  NAND2_X1 U749 ( .A1(n672), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U750 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U751 ( .A1(G220), .A2(G219), .ZN(n673) );
  XOR2_X1 U752 ( .A(KEYINPUT22), .B(n673), .Z(n674) );
  NOR2_X1 U753 ( .A1(G218), .A2(n674), .ZN(n675) );
  NAND2_X1 U754 ( .A1(G96), .A2(n675), .ZN(n829) );
  NAND2_X1 U755 ( .A1(n829), .A2(G2106), .ZN(n679) );
  NAND2_X1 U756 ( .A1(G69), .A2(G120), .ZN(n676) );
  NOR2_X1 U757 ( .A1(G237), .A2(n676), .ZN(n677) );
  NAND2_X1 U758 ( .A1(G108), .A2(n677), .ZN(n830) );
  NAND2_X1 U759 ( .A1(n830), .A2(G567), .ZN(n678) );
  NAND2_X1 U760 ( .A1(n679), .A2(n678), .ZN(n917) );
  NAND2_X1 U761 ( .A1(G661), .A2(G483), .ZN(n680) );
  NOR2_X1 U762 ( .A1(n917), .A2(n680), .ZN(n828) );
  NAND2_X1 U763 ( .A1(n828), .A2(G36), .ZN(G176) );
  INV_X1 U764 ( .A(G166), .ZN(G303) );
  NOR2_X1 U765 ( .A1(G1976), .A2(G288), .ZN(n681) );
  XOR2_X1 U766 ( .A(KEYINPUT103), .B(n681), .Z(n920) );
  INV_X1 U767 ( .A(n786), .ZN(n683) );
  NAND2_X2 U768 ( .A1(n785), .A2(n683), .ZN(n728) );
  INV_X1 U769 ( .A(G1996), .ZN(n972) );
  NOR2_X1 U770 ( .A1(n728), .A2(n972), .ZN(n685) );
  XNOR2_X1 U771 ( .A(n685), .B(n684), .ZN(n687) );
  NAND2_X1 U772 ( .A1(n728), .A2(G1341), .ZN(n686) );
  NAND2_X1 U773 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U774 ( .A1(n923), .A2(n688), .ZN(n690) );
  XNOR2_X1 U775 ( .A(n690), .B(n689), .ZN(n695) );
  NAND2_X1 U776 ( .A1(G1348), .A2(n728), .ZN(n692) );
  INV_X1 U777 ( .A(n728), .ZN(n711) );
  NAND2_X1 U778 ( .A1(n711), .A2(G2067), .ZN(n691) );
  NAND2_X1 U779 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U780 ( .A(n693), .B(KEYINPUT97), .Z(n696) );
  NAND2_X1 U781 ( .A1(n695), .A2(n694), .ZN(n699) );
  NAND2_X1 U782 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U783 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U784 ( .A(n700), .B(KEYINPUT98), .ZN(n705) );
  NAND2_X1 U785 ( .A1(n711), .A2(G2072), .ZN(n701) );
  XNOR2_X1 U786 ( .A(n701), .B(KEYINPUT27), .ZN(n703) );
  AND2_X1 U787 ( .A1(G1956), .A2(n728), .ZN(n702) );
  NOR2_X1 U788 ( .A1(n703), .A2(n702), .ZN(n706) );
  NAND2_X1 U789 ( .A1(n706), .A2(n928), .ZN(n704) );
  NAND2_X1 U790 ( .A1(n705), .A2(n704), .ZN(n709) );
  NOR2_X1 U791 ( .A1(n706), .A2(n928), .ZN(n707) );
  XOR2_X1 U792 ( .A(n707), .B(KEYINPUT28), .Z(n708) );
  NAND2_X1 U793 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U794 ( .A(n710), .B(KEYINPUT29), .ZN(n716) );
  XNOR2_X1 U795 ( .A(G1961), .B(KEYINPUT95), .ZN(n952) );
  NAND2_X1 U796 ( .A1(n952), .A2(n728), .ZN(n713) );
  XNOR2_X1 U797 ( .A(G2078), .B(KEYINPUT25), .ZN(n971) );
  NAND2_X1 U798 ( .A1(n711), .A2(n971), .ZN(n712) );
  NAND2_X1 U799 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U800 ( .A(n714), .B(KEYINPUT96), .Z(n722) );
  NOR2_X1 U801 ( .A1(G301), .A2(n722), .ZN(n715) );
  NOR2_X1 U802 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U803 ( .A(n717), .B(KEYINPUT99), .ZN(n727) );
  NAND2_X1 U804 ( .A1(G8), .A2(n728), .ZN(n768) );
  NOR2_X1 U805 ( .A1(G1966), .A2(n768), .ZN(n743) );
  NOR2_X1 U806 ( .A1(G2084), .A2(n728), .ZN(n738) );
  NOR2_X1 U807 ( .A1(n743), .A2(n738), .ZN(n718) );
  NAND2_X1 U808 ( .A1(G8), .A2(n718), .ZN(n719) );
  XNOR2_X1 U809 ( .A(KEYINPUT30), .B(n719), .ZN(n720) );
  NOR2_X1 U810 ( .A1(G168), .A2(n720), .ZN(n721) );
  XNOR2_X1 U811 ( .A(n721), .B(KEYINPUT100), .ZN(n724) );
  AND2_X1 U812 ( .A1(G301), .A2(n722), .ZN(n723) );
  NOR2_X1 U813 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U814 ( .A(KEYINPUT31), .B(n725), .Z(n726) );
  NAND2_X1 U815 ( .A1(n727), .A2(n726), .ZN(n740) );
  NAND2_X1 U816 ( .A1(n740), .A2(G286), .ZN(n734) );
  NOR2_X1 U817 ( .A1(G1971), .A2(n768), .ZN(n730) );
  NOR2_X1 U818 ( .A1(G2090), .A2(n728), .ZN(n729) );
  NOR2_X1 U819 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U820 ( .A1(n731), .A2(G303), .ZN(n732) );
  XOR2_X1 U821 ( .A(KEYINPUT101), .B(n732), .Z(n733) );
  NAND2_X1 U822 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U823 ( .A(n735), .B(KEYINPUT102), .ZN(n736) );
  AND2_X1 U824 ( .A1(n736), .A2(G8), .ZN(n737) );
  XNOR2_X1 U825 ( .A(KEYINPUT32), .B(n737), .ZN(n745) );
  NAND2_X1 U826 ( .A1(G8), .A2(n738), .ZN(n739) );
  XNOR2_X1 U827 ( .A(n739), .B(KEYINPUT94), .ZN(n741) );
  NAND2_X1 U828 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U829 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U830 ( .A1(n920), .A2(n767), .ZN(n750) );
  NOR2_X1 U831 ( .A1(G1971), .A2(G303), .ZN(n746) );
  XOR2_X1 U832 ( .A(n746), .B(KEYINPUT104), .Z(n748) );
  INV_X1 U833 ( .A(KEYINPUT33), .ZN(n747) );
  AND2_X1 U834 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U835 ( .A1(n750), .A2(n749), .ZN(n760) );
  INV_X1 U836 ( .A(n768), .ZN(n751) );
  NAND2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n921) );
  AND2_X1 U838 ( .A1(n751), .A2(n921), .ZN(n752) );
  NOR2_X1 U839 ( .A1(KEYINPUT33), .A2(n752), .ZN(n754) );
  XNOR2_X1 U840 ( .A(G1981), .B(KEYINPUT106), .ZN(n753) );
  XNOR2_X1 U841 ( .A(n753), .B(G305), .ZN(n934) );
  NOR2_X1 U842 ( .A1(n754), .A2(n934), .ZN(n758) );
  NAND2_X1 U843 ( .A1(KEYINPUT33), .A2(n920), .ZN(n755) );
  NOR2_X1 U844 ( .A1(n768), .A2(n755), .ZN(n756) );
  XNOR2_X1 U845 ( .A(KEYINPUT105), .B(n756), .ZN(n757) );
  AND2_X1 U846 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U847 ( .A1(n760), .A2(n759), .ZN(n773) );
  NOR2_X1 U848 ( .A1(G2090), .A2(G303), .ZN(n761) );
  AND2_X1 U849 ( .A1(G8), .A2(n761), .ZN(n765) );
  NOR2_X1 U850 ( .A1(G1981), .A2(G305), .ZN(n762) );
  XNOR2_X1 U851 ( .A(n762), .B(KEYINPUT93), .ZN(n763) );
  XNOR2_X1 U852 ( .A(n763), .B(KEYINPUT24), .ZN(n764) );
  NOR2_X1 U853 ( .A1(n764), .A2(n768), .ZN(n769) );
  OR2_X1 U854 ( .A1(n765), .A2(n769), .ZN(n766) );
  OR2_X1 U855 ( .A1(n767), .A2(n766), .ZN(n771) );
  OR2_X1 U856 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U857 ( .A1(n771), .A2(n770), .ZN(n772) );
  AND2_X1 U858 ( .A1(n773), .A2(n772), .ZN(n808) );
  XNOR2_X1 U859 ( .A(G2067), .B(KEYINPUT37), .ZN(n818) );
  NAND2_X1 U860 ( .A1(G104), .A2(n863), .ZN(n775) );
  NAND2_X1 U861 ( .A1(G140), .A2(n553), .ZN(n774) );
  NAND2_X1 U862 ( .A1(n775), .A2(n774), .ZN(n777) );
  XOR2_X1 U863 ( .A(KEYINPUT34), .B(KEYINPUT89), .Z(n776) );
  XNOR2_X1 U864 ( .A(n777), .B(n776), .ZN(n783) );
  NAND2_X1 U865 ( .A1(n859), .A2(G128), .ZN(n778) );
  XNOR2_X1 U866 ( .A(n778), .B(KEYINPUT90), .ZN(n780) );
  NAND2_X1 U867 ( .A1(G116), .A2(n860), .ZN(n779) );
  NAND2_X1 U868 ( .A1(n780), .A2(n779), .ZN(n781) );
  XOR2_X1 U869 ( .A(KEYINPUT35), .B(n781), .Z(n782) );
  NOR2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U871 ( .A(KEYINPUT36), .B(n784), .ZN(n882) );
  NOR2_X1 U872 ( .A1(n818), .A2(n882), .ZN(n1003) );
  NOR2_X1 U873 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U874 ( .A(n787), .B(KEYINPUT88), .ZN(n820) );
  NAND2_X1 U875 ( .A1(n1003), .A2(n820), .ZN(n816) );
  INV_X1 U876 ( .A(n820), .ZN(n804) );
  NAND2_X1 U877 ( .A1(G129), .A2(n859), .ZN(n789) );
  NAND2_X1 U878 ( .A1(G141), .A2(n553), .ZN(n788) );
  NAND2_X1 U879 ( .A1(n789), .A2(n788), .ZN(n792) );
  NAND2_X1 U880 ( .A1(n863), .A2(G105), .ZN(n790) );
  XOR2_X1 U881 ( .A(KEYINPUT38), .B(n790), .Z(n791) );
  NOR2_X1 U882 ( .A1(n792), .A2(n791), .ZN(n794) );
  NAND2_X1 U883 ( .A1(G117), .A2(n860), .ZN(n793) );
  NAND2_X1 U884 ( .A1(n794), .A2(n793), .ZN(n876) );
  NAND2_X1 U885 ( .A1(G1996), .A2(n876), .ZN(n802) );
  NAND2_X1 U886 ( .A1(G119), .A2(n859), .ZN(n796) );
  NAND2_X1 U887 ( .A1(G131), .A2(n553), .ZN(n795) );
  NAND2_X1 U888 ( .A1(n796), .A2(n795), .ZN(n800) );
  NAND2_X1 U889 ( .A1(G95), .A2(n863), .ZN(n798) );
  NAND2_X1 U890 ( .A1(G107), .A2(n860), .ZN(n797) );
  NAND2_X1 U891 ( .A1(n798), .A2(n797), .ZN(n799) );
  OR2_X1 U892 ( .A1(n800), .A2(n799), .ZN(n869) );
  NAND2_X1 U893 ( .A1(G1991), .A2(n869), .ZN(n801) );
  NAND2_X1 U894 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U895 ( .A(KEYINPUT91), .B(n803), .ZN(n994) );
  NOR2_X1 U896 ( .A1(n804), .A2(n994), .ZN(n813) );
  INV_X1 U897 ( .A(n813), .ZN(n805) );
  NAND2_X1 U898 ( .A1(n816), .A2(n805), .ZN(n806) );
  XNOR2_X1 U899 ( .A(n806), .B(KEYINPUT92), .ZN(n807) );
  NOR2_X1 U900 ( .A1(n808), .A2(n807), .ZN(n810) );
  XNOR2_X1 U901 ( .A(G1986), .B(G290), .ZN(n932) );
  NAND2_X1 U902 ( .A1(n932), .A2(n820), .ZN(n809) );
  NAND2_X1 U903 ( .A1(n810), .A2(n809), .ZN(n823) );
  NOR2_X1 U904 ( .A1(G1996), .A2(n876), .ZN(n996) );
  NOR2_X1 U905 ( .A1(G1991), .A2(n869), .ZN(n992) );
  NOR2_X1 U906 ( .A1(G1986), .A2(G290), .ZN(n811) );
  NOR2_X1 U907 ( .A1(n992), .A2(n811), .ZN(n812) );
  NOR2_X1 U908 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U909 ( .A1(n996), .A2(n814), .ZN(n815) );
  XNOR2_X1 U910 ( .A(n815), .B(KEYINPUT39), .ZN(n817) );
  NAND2_X1 U911 ( .A1(n817), .A2(n816), .ZN(n819) );
  NAND2_X1 U912 ( .A1(n818), .A2(n882), .ZN(n1012) );
  NAND2_X1 U913 ( .A1(n819), .A2(n1012), .ZN(n821) );
  NAND2_X1 U914 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U915 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U916 ( .A(KEYINPUT40), .B(n824), .ZN(G329) );
  NAND2_X1 U917 ( .A1(G2106), .A2(n825), .ZN(G217) );
  AND2_X1 U918 ( .A1(G15), .A2(G2), .ZN(n826) );
  NAND2_X1 U919 ( .A1(G661), .A2(n826), .ZN(G259) );
  NAND2_X1 U920 ( .A1(G3), .A2(G1), .ZN(n827) );
  NAND2_X1 U921 ( .A1(n828), .A2(n827), .ZN(G188) );
  INV_X1 U923 ( .A(G120), .ZN(G236) );
  INV_X1 U924 ( .A(G96), .ZN(G221) );
  INV_X1 U925 ( .A(G69), .ZN(G235) );
  NOR2_X1 U926 ( .A1(n830), .A2(n829), .ZN(G325) );
  INV_X1 U927 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U928 ( .A(G2446), .B(G2454), .ZN(n840) );
  XOR2_X1 U929 ( .A(G2430), .B(KEYINPUT108), .Z(n832) );
  XNOR2_X1 U930 ( .A(G2451), .B(G2443), .ZN(n831) );
  XNOR2_X1 U931 ( .A(n832), .B(n831), .ZN(n836) );
  XOR2_X1 U932 ( .A(G2427), .B(KEYINPUT107), .Z(n834) );
  XNOR2_X1 U933 ( .A(G1341), .B(G1348), .ZN(n833) );
  XNOR2_X1 U934 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U935 ( .A(n836), .B(n835), .Z(n838) );
  XNOR2_X1 U936 ( .A(G2438), .B(G2435), .ZN(n837) );
  XNOR2_X1 U937 ( .A(n838), .B(n837), .ZN(n839) );
  XNOR2_X1 U938 ( .A(n840), .B(n839), .ZN(n841) );
  NAND2_X1 U939 ( .A1(n841), .A2(G14), .ZN(n842) );
  XNOR2_X1 U940 ( .A(KEYINPUT109), .B(n842), .ZN(G401) );
  NAND2_X1 U941 ( .A1(G100), .A2(n863), .ZN(n844) );
  NAND2_X1 U942 ( .A1(G112), .A2(n860), .ZN(n843) );
  NAND2_X1 U943 ( .A1(n844), .A2(n843), .ZN(n850) );
  NAND2_X1 U944 ( .A1(n859), .A2(G124), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n845), .B(KEYINPUT44), .ZN(n847) );
  NAND2_X1 U946 ( .A1(G136), .A2(n553), .ZN(n846) );
  NAND2_X1 U947 ( .A1(n847), .A2(n846), .ZN(n848) );
  XOR2_X1 U948 ( .A(KEYINPUT113), .B(n848), .Z(n849) );
  NOR2_X1 U949 ( .A1(n850), .A2(n849), .ZN(G162) );
  NAND2_X1 U950 ( .A1(G103), .A2(n863), .ZN(n852) );
  NAND2_X1 U951 ( .A1(G139), .A2(n553), .ZN(n851) );
  NAND2_X1 U952 ( .A1(n852), .A2(n851), .ZN(n858) );
  NAND2_X1 U953 ( .A1(G115), .A2(n860), .ZN(n853) );
  XNOR2_X1 U954 ( .A(n853), .B(KEYINPUT114), .ZN(n855) );
  NAND2_X1 U955 ( .A1(G127), .A2(n859), .ZN(n854) );
  NAND2_X1 U956 ( .A1(n855), .A2(n854), .ZN(n856) );
  XOR2_X1 U957 ( .A(KEYINPUT47), .B(n856), .Z(n857) );
  NOR2_X1 U958 ( .A1(n858), .A2(n857), .ZN(n1005) );
  NAND2_X1 U959 ( .A1(G130), .A2(n859), .ZN(n862) );
  NAND2_X1 U960 ( .A1(G118), .A2(n860), .ZN(n861) );
  NAND2_X1 U961 ( .A1(n862), .A2(n861), .ZN(n868) );
  NAND2_X1 U962 ( .A1(G106), .A2(n863), .ZN(n865) );
  NAND2_X1 U963 ( .A1(G142), .A2(n553), .ZN(n864) );
  NAND2_X1 U964 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U965 ( .A(n866), .B(KEYINPUT45), .Z(n867) );
  NOR2_X1 U966 ( .A1(n868), .A2(n867), .ZN(n870) );
  XNOR2_X1 U967 ( .A(n870), .B(n869), .ZN(n874) );
  XOR2_X1 U968 ( .A(KEYINPUT46), .B(KEYINPUT115), .Z(n872) );
  XNOR2_X1 U969 ( .A(KEYINPUT116), .B(KEYINPUT48), .ZN(n871) );
  XNOR2_X1 U970 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U971 ( .A(n874), .B(n873), .Z(n879) );
  XOR2_X1 U972 ( .A(G160), .B(G162), .Z(n875) );
  XNOR2_X1 U973 ( .A(n876), .B(n875), .ZN(n877) );
  XNOR2_X1 U974 ( .A(G164), .B(n877), .ZN(n878) );
  XNOR2_X1 U975 ( .A(n879), .B(n878), .ZN(n880) );
  XOR2_X1 U976 ( .A(n1005), .B(n880), .Z(n881) );
  XNOR2_X1 U977 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U978 ( .A(n883), .B(n1000), .ZN(n884) );
  NOR2_X1 U979 ( .A1(G37), .A2(n884), .ZN(G395) );
  XOR2_X1 U980 ( .A(KEYINPUT112), .B(KEYINPUT42), .Z(n886) );
  XNOR2_X1 U981 ( .A(G2678), .B(G2096), .ZN(n885) );
  XNOR2_X1 U982 ( .A(n886), .B(n885), .ZN(n887) );
  XOR2_X1 U983 ( .A(n887), .B(KEYINPUT43), .Z(n889) );
  XNOR2_X1 U984 ( .A(G2067), .B(G2090), .ZN(n888) );
  XNOR2_X1 U985 ( .A(n889), .B(n888), .ZN(n893) );
  XOR2_X1 U986 ( .A(G2100), .B(G2084), .Z(n891) );
  XNOR2_X1 U987 ( .A(G2078), .B(G2072), .ZN(n890) );
  XNOR2_X1 U988 ( .A(n891), .B(n890), .ZN(n892) );
  XOR2_X1 U989 ( .A(n893), .B(n892), .Z(n895) );
  XNOR2_X1 U990 ( .A(KEYINPUT111), .B(KEYINPUT110), .ZN(n894) );
  XNOR2_X1 U991 ( .A(n895), .B(n894), .ZN(G227) );
  XOR2_X1 U992 ( .A(G1976), .B(G1981), .Z(n897) );
  XNOR2_X1 U993 ( .A(G1966), .B(G1956), .ZN(n896) );
  XNOR2_X1 U994 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U995 ( .A(n898), .B(KEYINPUT41), .Z(n900) );
  XNOR2_X1 U996 ( .A(G1996), .B(G1991), .ZN(n899) );
  XNOR2_X1 U997 ( .A(n900), .B(n899), .ZN(n904) );
  XOR2_X1 U998 ( .A(G2474), .B(G1971), .Z(n902) );
  XNOR2_X1 U999 ( .A(G1986), .B(G1961), .ZN(n901) );
  XNOR2_X1 U1000 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(G229) );
  XOR2_X1 U1002 ( .A(KEYINPUT117), .B(n905), .Z(n907) );
  XNOR2_X1 U1003 ( .A(G171), .B(n918), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1005 ( .A(n908), .B(G286), .Z(n909) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n909), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(KEYINPUT118), .B(n910), .ZN(G397) );
  NOR2_X1 U1008 ( .A1(G401), .A2(n917), .ZN(n914) );
  NOR2_X1 U1009 ( .A1(G227), .A2(G229), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(KEYINPUT49), .B(n911), .ZN(n912) );
  NOR2_X1 U1011 ( .A1(G395), .A2(n912), .ZN(n913) );
  NAND2_X1 U1012 ( .A1(n914), .A2(n913), .ZN(n915) );
  NOR2_X1 U1013 ( .A1(n915), .A2(G397), .ZN(n916) );
  XNOR2_X1 U1014 ( .A(n916), .B(KEYINPUT119), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(n917), .ZN(G319) );
  INV_X1 U1017 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1018 ( .A(G16), .B(KEYINPUT56), .Z(n941) );
  XOR2_X1 U1019 ( .A(G1348), .B(n918), .Z(n919) );
  NOR2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n927) );
  XNOR2_X1 U1021 ( .A(G166), .B(G1971), .ZN(n922) );
  NAND2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(n925) );
  XNOR2_X1 U1023 ( .A(G1341), .B(n923), .ZN(n924) );
  NOR2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n939) );
  XNOR2_X1 U1026 ( .A(n928), .B(G1956), .ZN(n930) );
  XNOR2_X1 U1027 ( .A(G171), .B(G1961), .ZN(n929) );
  NAND2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n937) );
  XOR2_X1 U1030 ( .A(G168), .B(G1966), .Z(n933) );
  NOR2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1032 ( .A(KEYINPUT57), .B(n935), .Z(n936) );
  NAND2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n1021) );
  XNOR2_X1 U1036 ( .A(KEYINPUT125), .B(G1981), .ZN(n942) );
  XNOR2_X1 U1037 ( .A(n942), .B(G6), .ZN(n947) );
  XOR2_X1 U1038 ( .A(G1348), .B(KEYINPUT59), .Z(n943) );
  XNOR2_X1 U1039 ( .A(G4), .B(n943), .ZN(n945) );
  XNOR2_X1 U1040 ( .A(G20), .B(G1956), .ZN(n944) );
  NOR2_X1 U1041 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n950) );
  XNOR2_X1 U1043 ( .A(KEYINPUT124), .B(G1341), .ZN(n948) );
  XNOR2_X1 U1044 ( .A(G19), .B(n948), .ZN(n949) );
  NOR2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1046 ( .A(KEYINPUT60), .B(n951), .ZN(n962) );
  XNOR2_X1 U1047 ( .A(KEYINPUT123), .B(G5), .ZN(n953) );
  XNOR2_X1 U1048 ( .A(n953), .B(n952), .ZN(n960) );
  XNOR2_X1 U1049 ( .A(G1971), .B(G22), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(G23), .B(G1976), .ZN(n954) );
  NOR2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n957) );
  XOR2_X1 U1052 ( .A(G1986), .B(G24), .Z(n956) );
  NAND2_X1 U1053 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1054 ( .A(KEYINPUT58), .B(n958), .ZN(n959) );
  NOR2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(G21), .B(G1966), .ZN(n963) );
  NOR2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1059 ( .A(KEYINPUT61), .B(n965), .Z(n966) );
  NOR2_X1 U1060 ( .A1(G16), .A2(n966), .ZN(n990) );
  INV_X1 U1061 ( .A(KEYINPUT55), .ZN(n1015) );
  XNOR2_X1 U1062 ( .A(G2090), .B(G35), .ZN(n981) );
  XOR2_X1 U1063 ( .A(G1991), .B(G25), .Z(n967) );
  NAND2_X1 U1064 ( .A1(n967), .A2(G28), .ZN(n978) );
  XNOR2_X1 U1065 ( .A(G2067), .B(G26), .ZN(n969) );
  XNOR2_X1 U1066 ( .A(G2072), .B(G33), .ZN(n968) );
  NOR2_X1 U1067 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1068 ( .A(KEYINPUT122), .B(n970), .ZN(n976) );
  XOR2_X1 U1069 ( .A(n971), .B(G27), .Z(n974) );
  XOR2_X1 U1070 ( .A(n972), .B(G32), .Z(n973) );
  NOR2_X1 U1071 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n977) );
  NOR2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1074 ( .A(KEYINPUT53), .B(n979), .ZN(n980) );
  NOR2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n984) );
  XOR2_X1 U1076 ( .A(G2084), .B(G34), .Z(n982) );
  XNOR2_X1 U1077 ( .A(KEYINPUT54), .B(n982), .ZN(n983) );
  NAND2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1079 ( .A(n1015), .B(n985), .ZN(n987) );
  INV_X1 U1080 ( .A(G29), .ZN(n986) );
  NAND2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1082 ( .A1(G11), .A2(n988), .ZN(n989) );
  NOR2_X1 U1083 ( .A1(n990), .A2(n989), .ZN(n1019) );
  XOR2_X1 U1084 ( .A(G160), .B(G2084), .Z(n991) );
  NOR2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n999) );
  XOR2_X1 U1087 ( .A(G2090), .B(G162), .Z(n995) );
  NOR2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1089 ( .A(n997), .B(KEYINPUT51), .ZN(n998) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1001) );
  NAND2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NOR2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1093 ( .A(KEYINPUT120), .B(n1004), .Z(n1010) );
  XOR2_X1 U1094 ( .A(G2072), .B(n1005), .Z(n1007) );
  XOR2_X1 U1095 ( .A(G164), .B(G2078), .Z(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1097 ( .A(KEYINPUT50), .B(n1008), .Z(n1009) );
  NOR2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(n1013), .B(KEYINPUT121), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(KEYINPUT52), .B(n1014), .ZN(n1016) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1103 ( .A1(n1017), .A2(G29), .ZN(n1018) );
  NAND2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1105 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1106 ( .A(KEYINPUT126), .B(n1022), .Z(n1023) );
  XNOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1023), .ZN(G150) );
  INV_X1 U1108 ( .A(G150), .ZN(G311) );
endmodule

