//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 0 1 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 1 0 1 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1 1 1 1 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1254, new_n1255,
    new_n1256, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1300, new_n1301, new_n1302;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AND2_X1   g0005(.A1(KEYINPUT64), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(KEYINPUT64), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT65), .Z(new_n211));
  NAND2_X1  g0011(.A1(new_n203), .A2(G50), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G1), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT0), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n221));
  INV_X1    g0021(.A(G77), .ZN(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  INV_X1    g0023(.A(G107), .ZN(new_n224));
  INV_X1    g0024(.A(G264), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n217), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n220), .B1(KEYINPUT1), .B2(new_n230), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n213), .B(new_n231), .C1(KEYINPUT1), .C2(new_n230), .ZN(G361));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT66), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT67), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  INV_X1    g0050(.A(G41), .ZN(new_n251));
  OAI211_X1 g0051(.A(G1), .B(G13), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G45), .ZN(new_n253));
  AOI21_X1  g0053(.A(G1), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n252), .A2(G274), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT68), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT68), .ZN(new_n257));
  NAND4_X1  g0057(.A1(new_n252), .A2(new_n257), .A3(new_n254), .A4(G274), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n209), .B1(G33), .B2(G41), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(new_n254), .ZN(new_n261));
  OR2_X1    g0061(.A1(KEYINPUT69), .A2(G226), .ZN(new_n262));
  NAND2_X1  g0062(.A1(KEYINPUT69), .A2(G226), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT3), .B(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G1698), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT70), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n267), .B(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT71), .B(G223), .ZN(new_n270));
  AND2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n266), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G222), .ZN(new_n274));
  OAI22_X1  g0074(.A1(new_n273), .A2(new_n274), .B1(new_n222), .B2(new_n266), .ZN(new_n275));
  OR2_X1    g0075(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n265), .B1(new_n276), .B2(new_n260), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(G169), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n209), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n208), .A2(G33), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT8), .B(G58), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n284));
  INV_X1    g0084(.A(G150), .ZN(new_n285));
  NOR2_X1   g0085(.A1(G20), .A2(G33), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n284), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n280), .B1(new_n283), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(KEYINPUT72), .ZN(new_n290));
  INV_X1    g0090(.A(G13), .ZN(new_n291));
  NOR3_X1   g0091(.A1(new_n291), .A2(new_n215), .A3(G1), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(new_n280), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n214), .A2(G20), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n293), .A2(G50), .A3(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n291), .A2(G1), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G20), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n290), .B(new_n295), .C1(G50), .C2(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n289), .A2(KEYINPUT72), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n278), .A2(new_n300), .ZN(new_n301));
  OR2_X1    g0101(.A1(new_n301), .A2(KEYINPUT73), .ZN(new_n302));
  INV_X1    g0102(.A(G179), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n277), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n301), .A2(KEYINPUT73), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n302), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G200), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n277), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n308), .B1(G190), .B2(new_n277), .ZN(new_n309));
  XOR2_X1   g0109(.A(new_n300), .B(KEYINPUT9), .Z(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT76), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT10), .ZN(new_n313));
  OR2_X1    g0113(.A1(new_n312), .A2(KEYINPUT10), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n311), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n309), .A2(new_n312), .A3(KEYINPUT10), .A4(new_n310), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n306), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G226), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G1698), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n319), .B1(G223), .B2(G1698), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT3), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G33), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G87), .ZN(new_n325));
  OAI22_X1  g0125(.A1(new_n320), .A2(new_n324), .B1(new_n250), .B2(new_n325), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n256), .A2(new_n258), .B1(new_n326), .B2(new_n260), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT79), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n261), .A2(new_n328), .A3(G232), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n214), .B1(G41), .B2(G45), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n252), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G232), .ZN(new_n332));
  OAI21_X1  g0132(.A(KEYINPUT79), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n327), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G169), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT80), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n327), .A2(new_n303), .A3(new_n334), .ZN(new_n339));
  AND3_X1   g0139(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n338), .B1(new_n337), .B2(new_n339), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n282), .B1(new_n214), .B2(G20), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n343), .A2(new_n293), .B1(new_n292), .B2(new_n282), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT78), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT64), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n215), .ZN(new_n348));
  NAND2_X1  g0148(.A1(KEYINPUT64), .A2(G20), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(KEYINPUT7), .A3(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n321), .A2(G33), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT77), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n351), .B1(new_n352), .B2(new_n322), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n321), .A2(KEYINPUT77), .A3(G33), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n350), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(G20), .B1(new_n322), .B2(new_n323), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n356), .A2(KEYINPUT7), .ZN(new_n357));
  OAI21_X1  g0157(.A(G68), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  XNOR2_X1  g0158(.A(G58), .B(G68), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n359), .A2(G20), .B1(G159), .B2(new_n286), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT16), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT7), .ZN(new_n362));
  OAI21_X1  g0162(.A(G68), .B1(new_n356), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n348), .A2(new_n349), .ZN(new_n364));
  NOR3_X1   g0164(.A1(new_n364), .A2(new_n266), .A3(KEYINPUT7), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n360), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT16), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n280), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n346), .B1(new_n361), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n280), .ZN(new_n370));
  INV_X1    g0170(.A(new_n360), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n324), .A2(new_n215), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n202), .B1(new_n372), .B2(KEYINPUT7), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n324), .A2(new_n208), .A3(new_n362), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n371), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n370), .B1(new_n375), .B2(KEYINPUT16), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n322), .A2(new_n352), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n377), .A2(new_n323), .A3(new_n354), .ZN(new_n378));
  INV_X1    g0178(.A(new_n350), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n372), .A2(new_n362), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n202), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n367), .B1(new_n382), .B2(new_n371), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n376), .A2(new_n383), .A3(KEYINPUT78), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n345), .B1(new_n369), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT18), .B1(new_n342), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n369), .A2(new_n384), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n344), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n337), .A2(new_n339), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT80), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT18), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n388), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(KEYINPUT81), .B1(new_n335), .B2(G190), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n335), .A2(new_n307), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT81), .ZN(new_n397));
  INV_X1    g0197(.A(G190), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n327), .A2(new_n397), .A3(new_n398), .A4(new_n334), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n395), .A2(new_n396), .A3(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n387), .A2(new_n344), .A3(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT17), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n385), .A2(KEYINPUT17), .A3(new_n400), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n386), .A2(new_n394), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n332), .A2(G1698), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(G226), .B2(G1698), .ZN(new_n407));
  INV_X1    g0207(.A(G97), .ZN(new_n408));
  OAI22_X1  g0208(.A1(new_n407), .A2(new_n324), .B1(new_n250), .B2(new_n408), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n409), .A2(new_n260), .B1(G238), .B2(new_n261), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n259), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n411), .A2(KEYINPUT13), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n411), .A2(KEYINPUT13), .ZN(new_n413));
  OR2_X1    g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n414), .A2(G200), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n414), .A2(new_n398), .ZN(new_n416));
  INV_X1    g0216(.A(new_n296), .ZN(new_n417));
  NOR4_X1   g0217(.A1(new_n417), .A2(KEYINPUT12), .A3(new_n215), .A4(G68), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT75), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n297), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n292), .A2(KEYINPUT75), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n202), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n418), .B1(new_n424), .B2(KEYINPUT12), .ZN(new_n425));
  INV_X1    g0225(.A(new_n281), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(G77), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n286), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n370), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n425), .B1(KEYINPUT11), .B2(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n423), .A2(new_n280), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n431), .A2(G68), .A3(new_n294), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n430), .B(new_n432), .C1(KEYINPUT11), .C2(new_n429), .ZN(new_n433));
  OR3_X1    g0233(.A1(new_n415), .A2(new_n416), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT14), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n435), .B(G169), .C1(new_n412), .C2(new_n413), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(new_n414), .B2(new_n303), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n435), .B1(new_n414), .B2(G169), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n433), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n431), .A2(G77), .A3(new_n294), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(G77), .B2(new_n422), .ZN(new_n441));
  OAI22_X1  g0241(.A1(new_n208), .A2(new_n222), .B1(new_n282), .B2(new_n287), .ZN(new_n442));
  OR2_X1    g0242(.A1(new_n442), .A2(KEYINPUT74), .ZN(new_n443));
  XNOR2_X1  g0243(.A(KEYINPUT15), .B(G87), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n442), .A2(KEYINPUT74), .B1(new_n426), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n370), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n441), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n259), .B1(new_n223), .B2(new_n331), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  OAI22_X1  g0251(.A1(new_n273), .A2(new_n332), .B1(new_n224), .B2(new_n266), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n452), .B1(new_n269), .B2(G238), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n451), .B(new_n303), .C1(new_n453), .C2(new_n252), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n453), .A2(new_n252), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n336), .B1(new_n455), .B2(new_n450), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n449), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(G200), .B1(new_n455), .B2(new_n450), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n451), .B(G190), .C1(new_n453), .C2(new_n252), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n448), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n434), .A2(new_n439), .A3(new_n461), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n317), .A2(new_n405), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n208), .A2(new_n266), .A3(G87), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT22), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(KEYINPUT88), .ZN(new_n466));
  XNOR2_X1  g0266(.A(new_n464), .B(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(KEYINPUT23), .A2(G107), .ZN(new_n468));
  AOI21_X1  g0268(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n468), .B1(new_n469), .B2(G20), .ZN(new_n470));
  NOR2_X1   g0270(.A1(KEYINPUT23), .A2(G107), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n470), .B1(new_n364), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT24), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n370), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n475), .B1(new_n474), .B2(new_n473), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n292), .A2(new_n224), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT89), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n477), .A2(new_n478), .A3(KEYINPUT25), .ZN(new_n479));
  XOR2_X1   g0279(.A(KEYINPUT89), .B(KEYINPUT25), .Z(new_n480));
  NAND2_X1  g0280(.A1(new_n214), .A2(G33), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n293), .A2(new_n481), .ZN(new_n482));
  OAI221_X1 g0282(.A(new_n479), .B1(new_n477), .B2(new_n480), .C1(new_n482), .C2(new_n224), .ZN(new_n483));
  XOR2_X1   g0283(.A(new_n483), .B(KEYINPUT90), .Z(new_n484));
  NAND3_X1  g0284(.A1(new_n266), .A2(G257), .A3(G1698), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G33), .A2(G294), .ZN(new_n486));
  INV_X1    g0286(.A(G250), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n485), .B(new_n486), .C1(new_n273), .C2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n260), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n214), .B(G45), .C1(new_n251), .C2(KEYINPUT5), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT84), .ZN(new_n491));
  XNOR2_X1  g0291(.A(new_n490), .B(new_n491), .ZN(new_n492));
  XNOR2_X1  g0292(.A(KEYINPUT85), .B(KEYINPUT5), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n251), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n492), .A2(G274), .A3(new_n252), .A4(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n490), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n260), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G264), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n489), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  OR2_X1    g0299(.A1(new_n499), .A2(new_n398), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(G200), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n476), .A2(new_n484), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(G107), .B1(new_n355), .B2(new_n357), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n286), .A2(G77), .ZN(new_n504));
  XNOR2_X1  g0304(.A(KEYINPUT82), .B(G107), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n408), .A2(new_n224), .A3(KEYINPUT6), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n507), .B1(KEYINPUT6), .B2(new_n408), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n506), .A2(new_n508), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n503), .B(new_n504), .C1(new_n208), .C2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n280), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n297), .A2(G97), .ZN(new_n514));
  INV_X1    g0314(.A(new_n482), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n514), .B1(new_n515), .B2(G97), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n497), .A2(G257), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n495), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n266), .A2(G244), .A3(new_n272), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT4), .ZN(new_n522));
  OR2_X1    g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n266), .A2(G250), .A3(G1698), .ZN(new_n524));
  NAND2_X1  g0324(.A1(G33), .A2(G283), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n521), .A2(new_n522), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT83), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n521), .A2(KEYINPUT83), .A3(new_n522), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n527), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n303), .B(new_n520), .C1(new_n532), .C2(new_n252), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n530), .A2(new_n531), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n534), .A2(new_n523), .A3(new_n526), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n519), .B1(new_n535), .B2(new_n260), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n517), .B(new_n533), .C1(G169), .C2(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(G190), .B(new_n520), .C1(new_n532), .C2(new_n252), .ZN(new_n538));
  INV_X1    g0338(.A(new_n516), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n539), .B1(new_n512), .B2(new_n280), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n538), .B(new_n540), .C1(new_n536), .C2(new_n307), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n502), .A2(new_n537), .A3(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n422), .A2(G116), .A3(new_n370), .A4(new_n481), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n208), .B(new_n525), .C1(G33), .C2(new_n408), .ZN(new_n544));
  INV_X1    g0344(.A(G116), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n279), .A2(new_n209), .B1(G20), .B2(new_n545), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n544), .A2(KEYINPUT20), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(KEYINPUT20), .B1(new_n544), .B2(new_n546), .ZN(new_n548));
  OAI221_X1 g0348(.A(new_n543), .B1(G116), .B2(new_n422), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n266), .A2(G257), .A3(new_n272), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n324), .A2(G303), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n550), .B(new_n551), .C1(new_n267), .C2(new_n225), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n260), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n497), .A2(G270), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(new_n495), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n549), .B1(G200), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(new_n398), .B2(new_n555), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n549), .A2(KEYINPUT21), .A3(G169), .A4(new_n555), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n553), .A2(new_n495), .A3(G179), .A4(new_n554), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n549), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n549), .A2(G169), .A3(new_n555), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT21), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AND3_X1   g0365(.A1(new_n557), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n499), .A2(new_n336), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(G179), .B2(new_n499), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n568), .B1(new_n476), .B2(new_n484), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n266), .A2(G238), .A3(new_n272), .ZN(new_n570));
  NAND2_X1  g0370(.A1(G33), .A2(G116), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n570), .B(new_n571), .C1(new_n267), .C2(new_n223), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n260), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n214), .A2(G45), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n574), .A2(G274), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(KEYINPUT86), .B2(new_n487), .ZN(new_n576));
  NAND2_X1  g0376(.A1(KEYINPUT86), .A2(G250), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n252), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n573), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n336), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(G179), .B2(new_n580), .ZN(new_n582));
  NAND3_X1  g0382(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n348), .A2(new_n349), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n325), .A2(new_n408), .A3(new_n224), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(KEYINPUT87), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n208), .A2(new_n266), .A3(G68), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n348), .A2(G33), .A3(G97), .A4(new_n349), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT19), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT87), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n584), .A2(new_n592), .A3(new_n585), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n587), .A2(new_n588), .A3(new_n591), .A4(new_n593), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n594), .A2(new_n280), .B1(new_n423), .B2(new_n444), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n515), .A2(new_n445), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n582), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n580), .A2(G200), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n573), .A2(G190), .A3(new_n579), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n423), .A2(new_n444), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n515), .A2(G87), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n591), .A2(new_n588), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n584), .A2(new_n592), .A3(new_n585), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n592), .B1(new_n584), .B2(new_n585), .ZN(new_n607));
  NOR3_X1   g0407(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n603), .B(new_n604), .C1(new_n608), .C2(new_n370), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n602), .A2(new_n609), .ZN(new_n610));
  NOR3_X1   g0410(.A1(new_n569), .A2(new_n599), .A3(new_n610), .ZN(new_n611));
  AND4_X1   g0411(.A1(new_n463), .A2(new_n542), .A3(new_n566), .A4(new_n611), .ZN(G372));
  NAND2_X1  g0412(.A1(new_n386), .A2(new_n394), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT95), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n386), .A2(new_n394), .A3(KEYINPUT95), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n439), .A2(new_n457), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n403), .A2(new_n404), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n619), .A2(new_n621), .A3(new_n434), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n315), .B(new_n316), .C1(new_n618), .C2(new_n622), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n623), .A2(new_n306), .ZN(new_n624));
  INV_X1    g0424(.A(new_n463), .ZN(new_n625));
  OR3_X1    g0425(.A1(new_n537), .A2(new_n610), .A3(new_n599), .ZN(new_n626));
  XOR2_X1   g0426(.A(KEYINPUT94), .B(KEYINPUT26), .Z(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n599), .ZN(new_n630));
  INV_X1    g0430(.A(new_n600), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n609), .A2(KEYINPUT91), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT91), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n595), .A2(new_n633), .A3(new_n604), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n631), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT92), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n601), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AOI211_X1 g0437(.A(KEYINPUT92), .B(new_n631), .C1(new_n632), .C2(new_n634), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n630), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT93), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n609), .A2(KEYINPUT91), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n633), .B1(new_n595), .B2(new_n604), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n600), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(KEYINPUT92), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n635), .A2(new_n636), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(new_n601), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT93), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n646), .A2(new_n647), .A3(new_n630), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n537), .B1(new_n640), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n629), .B1(new_n649), .B2(KEYINPUT26), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n640), .A2(new_n648), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n562), .A2(new_n565), .ZN(new_n652));
  INV_X1    g0452(.A(new_n569), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n654), .A2(new_n542), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n599), .B1(new_n651), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n650), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n624), .B1(new_n625), .B2(new_n658), .ZN(G369));
  NAND2_X1  g0459(.A1(new_n562), .A2(new_n565), .ZN(new_n660));
  OR3_X1    g0460(.A1(new_n364), .A2(new_n417), .A3(KEYINPUT27), .ZN(new_n661));
  OAI21_X1  g0461(.A(KEYINPUT27), .B1(new_n364), .B2(new_n417), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n661), .A2(G213), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(G343), .ZN(new_n664));
  XNOR2_X1  g0464(.A(new_n664), .B(KEYINPUT96), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT97), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n666), .B(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n502), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n665), .B1(new_n484), .B2(new_n476), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n653), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n569), .A2(new_n665), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n668), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n672), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n665), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n549), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n566), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n652), .B2(new_n678), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(G330), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n673), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n676), .A2(new_n683), .ZN(G399));
  INV_X1    g0484(.A(new_n218), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(G41), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n585), .A2(G116), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G1), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n212), .B2(new_n687), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT28), .ZN(new_n691));
  INV_X1    g0491(.A(new_n537), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n651), .A2(KEYINPUT26), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n626), .A2(new_n627), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(KEYINPUT99), .B1(new_n651), .B2(new_n655), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n651), .A2(KEYINPUT99), .A3(new_n655), .ZN(new_n697));
  OAI211_X1 g0497(.A(new_n695), .B(new_n630), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n698), .A2(KEYINPUT29), .A3(new_n665), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n657), .A2(new_n665), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT29), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT98), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n489), .A2(new_n498), .ZN(new_n705));
  NOR3_X1   g0505(.A1(new_n559), .A2(new_n705), .A3(new_n580), .ZN(new_n706));
  AOI21_X1  g0506(.A(KEYINPUT30), .B1(new_n706), .B2(new_n536), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n499), .A2(new_n555), .A3(new_n303), .A4(new_n580), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n536), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n706), .A2(new_n536), .A3(KEYINPUT30), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n665), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n704), .B1(new_n712), .B2(KEYINPUT31), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n542), .A2(new_n611), .A3(new_n566), .A4(new_n665), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT31), .ZN(new_n715));
  INV_X1    g0515(.A(new_n711), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n716), .A2(new_n707), .A3(new_n709), .ZN(new_n717));
  OAI211_X1 g0517(.A(KEYINPUT98), .B(new_n715), .C1(new_n717), .C2(new_n665), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n712), .A2(KEYINPUT31), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n713), .A2(new_n714), .A3(new_n718), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(G330), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n703), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n691), .B1(new_n723), .B2(G1), .ZN(G364));
  NOR2_X1   g0524(.A1(new_n364), .A2(new_n291), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G45), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G1), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n686), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n682), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(G330), .B2(new_n680), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n218), .A2(new_n266), .ZN(new_n731));
  INV_X1    g0531(.A(G355), .ZN(new_n732));
  OAI22_X1  g0532(.A1(new_n731), .A2(new_n732), .B1(G116), .B2(new_n218), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n685), .A2(new_n266), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n212), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n735), .B1(new_n253), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n248), .A2(G45), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n733), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(G13), .A2(G33), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(G20), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n209), .B1(G20), .B2(new_n336), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n728), .B1(new_n739), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n208), .A2(new_n303), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n747), .A2(new_n398), .A3(new_n307), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n748), .A2(KEYINPUT100), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(KEYINPUT100), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G77), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n307), .A2(G179), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n754), .A2(G20), .A3(G190), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n266), .B1(new_n755), .B2(new_n325), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n208), .A2(G190), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n303), .A2(new_n307), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G179), .A2(G200), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n208), .B1(G190), .B2(new_n760), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n759), .A2(new_n202), .B1(new_n761), .B2(new_n408), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n757), .A2(new_n754), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n756), .B(new_n762), .C1(G107), .C2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n747), .A2(G190), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n307), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(G200), .ZN(new_n768));
  AOI22_X1  g0568(.A1(G50), .A2(new_n767), .B1(new_n768), .B2(G58), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n757), .A2(new_n760), .ZN(new_n770));
  XOR2_X1   g0570(.A(KEYINPUT101), .B(G159), .Z(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT32), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n753), .A2(new_n765), .A3(new_n769), .A4(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n752), .A2(G311), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n768), .A2(G322), .ZN(new_n776));
  INV_X1    g0576(.A(G303), .ZN(new_n777));
  XOR2_X1   g0577(.A(KEYINPUT33), .B(G317), .Z(new_n778));
  OAI221_X1 g0578(.A(new_n324), .B1(new_n777), .B2(new_n755), .C1(new_n759), .C2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(G326), .B2(new_n767), .ZN(new_n780));
  INV_X1    g0580(.A(G283), .ZN(new_n781));
  INV_X1    g0581(.A(G329), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n781), .A2(new_n763), .B1(new_n770), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n761), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n783), .B1(G294), .B2(new_n784), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n775), .A2(new_n776), .A3(new_n780), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n774), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n746), .B1(new_n787), .B2(new_n743), .ZN(new_n788));
  INV_X1    g0588(.A(new_n742), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n788), .B1(new_n680), .B2(new_n789), .ZN(new_n790));
  AND2_X1   g0590(.A1(new_n730), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(G396));
  NAND2_X1  g0592(.A1(new_n449), .A2(new_n677), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n461), .A2(KEYINPUT103), .A3(new_n793), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n457), .A2(new_n793), .A3(new_n460), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT103), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(new_n665), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n639), .A2(KEYINPUT93), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n647), .B1(new_n646), .B2(new_n630), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n692), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT26), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n628), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n651), .A2(new_n655), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(new_n630), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n800), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(KEYINPUT104), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT104), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n657), .A2(new_n810), .A3(new_n800), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n457), .A2(new_n665), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n794), .A2(new_n797), .A3(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n700), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  OR2_X1    g0617(.A1(new_n817), .A2(new_n721), .ZN(new_n818));
  XOR2_X1   g0618(.A(new_n818), .B(KEYINPUT105), .Z(new_n819));
  AOI21_X1  g0619(.A(new_n728), .B1(new_n817), .B2(new_n721), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n743), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n741), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n728), .B1(G77), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n752), .A2(G116), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n767), .A2(G303), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n324), .B1(new_n224), .B2(new_n755), .C1(new_n761), .C2(new_n408), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(G294), .B2(new_n768), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n325), .A2(new_n763), .B1(new_n759), .B2(new_n781), .ZN(new_n829));
  INV_X1    g0629(.A(new_n770), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n829), .B1(G311), .B2(new_n830), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n825), .A2(new_n826), .A3(new_n828), .A4(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n759), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n767), .A2(G137), .B1(new_n833), .B2(G150), .ZN(new_n834));
  INV_X1    g0634(.A(new_n768), .ZN(new_n835));
  XNOR2_X1  g0635(.A(KEYINPUT102), .B(G143), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n834), .B1(new_n835), .B2(new_n836), .C1(new_n751), .C2(new_n771), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT34), .Z(new_n838));
  INV_X1    g0638(.A(G132), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n202), .A2(new_n763), .B1(new_n770), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(G50), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n266), .B1(new_n841), .B2(new_n755), .C1(new_n761), .C2(new_n201), .ZN(new_n842));
  OR2_X1    g0642(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n832), .B1(new_n838), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n824), .B1(new_n844), .B2(new_n743), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n741), .B2(new_n814), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n821), .A2(new_n846), .ZN(G384));
  INV_X1    g0647(.A(new_n511), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n545), .B(new_n211), .C1(new_n848), .C2(KEYINPUT35), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(KEYINPUT35), .B2(new_n848), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n850), .B(KEYINPUT36), .Z(new_n851));
  OAI211_X1 g0651(.A(new_n736), .B(G77), .C1(new_n201), .C2(new_n202), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n841), .A2(G68), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n214), .B(G13), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n457), .A2(new_n677), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n810), .B1(new_n657), .B2(new_n800), .ZN(new_n858));
  AOI211_X1 g0658(.A(KEYINPUT104), .B(new_n799), .C1(new_n650), .C2(new_n656), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT38), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n375), .A2(KEYINPUT16), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n344), .B1(new_n862), .B2(new_n368), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(KEYINPUT107), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n864), .A2(new_n663), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n405), .A2(KEYINPUT108), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n388), .B1(new_n392), .B2(new_n663), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n401), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT37), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n864), .B1(new_n392), .B2(new_n663), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n869), .B1(new_n385), .B2(new_n400), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n868), .A2(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n866), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT108), .B1(new_n405), .B2(new_n865), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n861), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n405), .A2(new_n865), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT108), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n878), .A2(KEYINPUT38), .A3(new_n866), .A4(new_n872), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n433), .A2(new_n677), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT106), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n881), .B(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n883), .A2(new_n439), .A3(new_n434), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n434), .A2(new_n439), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n881), .B(KEYINPUT106), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n860), .A2(new_n880), .A3(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n617), .A2(new_n663), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n615), .A2(new_n621), .A3(new_n616), .ZN(new_n892));
  INV_X1    g0692(.A(new_n663), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n385), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT109), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n869), .B1(new_n867), .B2(new_n896), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n897), .B(new_n868), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT38), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  NOR3_X1   g0699(.A1(new_n873), .A2(new_n861), .A3(new_n874), .ZN(new_n900));
  NOR3_X1   g0700(.A1(new_n899), .A2(new_n900), .A3(KEYINPUT39), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT39), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n902), .B1(new_n875), .B2(new_n879), .ZN(new_n903));
  NOR3_X1   g0703(.A1(new_n901), .A2(KEYINPUT110), .A3(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT110), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n880), .A2(KEYINPUT39), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n897), .A2(new_n401), .A3(new_n867), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n385), .B1(new_n342), .B2(new_n893), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT37), .B1(new_n908), .B2(KEYINPUT109), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n868), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n894), .B2(new_n892), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n902), .B(new_n879), .C1(new_n912), .C2(KEYINPUT38), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n905), .B1(new_n906), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n904), .A2(new_n914), .ZN(new_n915));
  OR2_X1    g0715(.A1(new_n439), .A2(new_n677), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n889), .B(new_n891), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n699), .A2(new_n702), .A3(new_n463), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n918), .A2(new_n624), .ZN(new_n919));
  XOR2_X1   g0719(.A(new_n917), .B(new_n919), .Z(new_n920));
  INV_X1    g0720(.A(KEYINPUT111), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n712), .B2(KEYINPUT31), .ZN(new_n922));
  OAI211_X1 g0722(.A(KEYINPUT111), .B(new_n715), .C1(new_n717), .C2(new_n665), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n922), .A2(new_n714), .A3(new_n923), .A4(new_n719), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT40), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n888), .A2(new_n924), .A3(new_n925), .A4(new_n814), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(new_n879), .B2(new_n875), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n888), .A2(new_n924), .A3(new_n814), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n899), .B2(new_n900), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n927), .B1(KEYINPUT40), .B2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n924), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n930), .B1(new_n625), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n879), .B1(new_n912), .B2(KEYINPUT38), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n925), .B1(new_n933), .B2(new_n928), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n463), .B(new_n924), .C1(new_n934), .C2(new_n927), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n932), .A2(G330), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n920), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n214), .B2(new_n725), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n920), .A2(new_n936), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n855), .B1(new_n938), .B2(new_n939), .ZN(G367));
  AOI21_X1  g0740(.A(new_n745), .B1(new_n685), .B2(new_n445), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n734), .A2(new_n240), .ZN(new_n942));
  AOI211_X1 g0742(.A(new_n686), .B(new_n727), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n784), .A2(G68), .ZN(new_n944));
  INV_X1    g0744(.A(G137), .ZN(new_n945));
  OAI221_X1 g0745(.A(new_n944), .B1(new_n759), .B2(new_n771), .C1(new_n945), .C2(new_n770), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n266), .B1(new_n755), .B2(new_n201), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(new_n764), .B2(G77), .ZN(new_n948));
  INV_X1    g0748(.A(new_n767), .ZN(new_n949));
  OAI221_X1 g0749(.A(new_n948), .B1(new_n835), .B2(new_n285), .C1(new_n949), .C2(new_n836), .ZN(new_n950));
  AOI211_X1 g0750(.A(new_n946), .B(new_n950), .C1(G50), .C2(new_n752), .ZN(new_n951));
  OR3_X1    g0751(.A1(new_n755), .A2(KEYINPUT46), .A3(new_n545), .ZN(new_n952));
  OAI21_X1  g0752(.A(KEYINPUT46), .B1(new_n755), .B2(new_n545), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n266), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n835), .B2(new_n777), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(G311), .B2(new_n767), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n751), .A2(new_n781), .ZN(new_n957));
  INV_X1    g0757(.A(G294), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n408), .A2(new_n763), .B1(new_n759), .B2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(G317), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n770), .A2(new_n960), .B1(new_n761), .B2(new_n224), .ZN(new_n961));
  NOR3_X1   g0761(.A1(new_n957), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n951), .B1(new_n956), .B2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT47), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n677), .A2(new_n632), .A3(new_n634), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n651), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n630), .B2(new_n965), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n943), .B1(new_n822), .B2(new_n964), .C1(new_n967), .C2(new_n789), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n537), .B(new_n541), .C1(new_n540), .C2(new_n665), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n969), .A2(new_n653), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n677), .B1(new_n970), .B2(new_n537), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n674), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n692), .A2(new_n677), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n969), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n976), .A2(KEYINPUT112), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(KEYINPUT112), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n977), .A2(KEYINPUT42), .A3(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(KEYINPUT42), .B1(new_n977), .B2(new_n978), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n972), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n982), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  NOR3_X1   g0786(.A1(new_n982), .A2(KEYINPUT113), .A3(new_n984), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT113), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n977), .A2(new_n978), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT42), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n971), .B1(new_n991), .B2(new_n979), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n988), .B1(new_n992), .B2(new_n983), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n986), .B1(new_n987), .B2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n975), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n683), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n996), .B(new_n986), .C1(new_n987), .C2(new_n993), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT44), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n676), .B2(new_n975), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n675), .A2(KEYINPUT44), .A3(new_n995), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n676), .A2(KEYINPUT45), .A3(new_n975), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT45), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n675), .B2(new_n995), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n1002), .A2(new_n1003), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  OR3_X1    g0807(.A1(new_n1007), .A2(KEYINPUT114), .A3(new_n683), .ZN(new_n1008));
  OAI21_X1  g0808(.A(KEYINPUT114), .B1(new_n1007), .B2(new_n683), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n683), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1010), .A2(KEYINPUT116), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT116), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n1007), .B2(new_n683), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1008), .B(new_n1009), .C1(new_n1011), .C2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT115), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n668), .B2(new_n673), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(new_n681), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(new_n973), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n723), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n723), .B1(new_n1014), .B2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n686), .B(KEYINPUT41), .Z(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n727), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n968), .B1(new_n1000), .B2(new_n1023), .ZN(G387));
  AOI22_X1  g0824(.A1(new_n767), .A2(G322), .B1(new_n833), .B2(G311), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1025), .B1(new_n960), .B2(new_n835), .C1(new_n751), .C2(new_n777), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT48), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n755), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n784), .A2(G283), .B1(new_n1030), .B2(G294), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1028), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT49), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n763), .A2(new_n545), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n266), .B(new_n1036), .C1(G326), .C2(new_n830), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1034), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n752), .A2(G68), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n767), .A2(G159), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n266), .B1(new_n222), .B2(new_n755), .C1(new_n763), .C2(new_n408), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(G50), .B2(new_n768), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n285), .A2(new_n770), .B1(new_n759), .B2(new_n282), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n761), .A2(new_n444), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1039), .A2(new_n1040), .A3(new_n1042), .A4(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n822), .B1(new_n1038), .B2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n673), .A2(new_n789), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n731), .A2(new_n688), .B1(G107), .B2(new_n218), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n237), .A2(new_n253), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n688), .ZN(new_n1051));
  AOI211_X1 g0851(.A(G45), .B(new_n1051), .C1(G68), .C2(G77), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n282), .A2(G50), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT50), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n735), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1049), .B1(new_n1050), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n728), .B1(new_n1056), .B2(new_n745), .ZN(new_n1057));
  NOR3_X1   g0857(.A1(new_n1047), .A2(new_n1048), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n1018), .B2(new_n727), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1019), .A2(new_n686), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n723), .A2(new_n1018), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1059), .B1(new_n1060), .B2(new_n1061), .ZN(G393));
  NOR2_X1   g0862(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1007), .A2(new_n683), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n727), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n245), .A2(new_n734), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n744), .B1(new_n408), .B2(new_n218), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n728), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n266), .B1(new_n202), .B2(new_n755), .C1(new_n763), .C2(new_n325), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n784), .A2(G77), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n770), .B2(new_n836), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1070), .B(new_n1072), .C1(G50), .C2(new_n833), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n282), .B2(new_n751), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(G150), .A2(new_n767), .B1(new_n768), .B2(G159), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT51), .ZN(new_n1076));
  INV_X1    g0876(.A(G322), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n770), .A2(new_n1077), .B1(new_n761), .B2(new_n545), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n324), .B1(new_n781), .B2(new_n755), .C1(new_n763), .C2(new_n224), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1078), .B(new_n1079), .C1(G303), .C2(new_n833), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n958), .B2(new_n751), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(G311), .A2(new_n768), .B1(new_n767), .B2(G317), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT52), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n1074), .A2(new_n1076), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1069), .B1(new_n1084), .B2(new_n743), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n975), .B2(new_n789), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1019), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1065), .A2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n686), .B1(new_n1014), .B2(new_n1019), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1066), .B(new_n1086), .C1(new_n1088), .C2(new_n1089), .ZN(G390));
  INV_X1    g0890(.A(KEYINPUT99), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n806), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n651), .A2(KEYINPUT99), .A3(new_n655), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n599), .B1(new_n693), .B2(new_n694), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n799), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1096), .A2(new_n856), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n888), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n916), .B(new_n933), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n888), .A2(G330), .A3(new_n720), .A4(new_n814), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n916), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n860), .B2(new_n888), .ZN(new_n1102));
  OAI21_X1  g0902(.A(KEYINPUT110), .B1(new_n901), .B2(new_n903), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n906), .A2(new_n913), .A3(new_n905), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1099), .B(new_n1100), .C1(new_n1102), .C2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n933), .A2(new_n916), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n698), .A2(new_n800), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n857), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1107), .B1(new_n1109), .B2(new_n888), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n856), .B1(new_n809), .B2(new_n811), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n916), .B1(new_n1111), .B2(new_n1098), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1110), .B1(new_n1112), .B2(new_n915), .ZN(new_n1113));
  INV_X1    g0913(.A(G330), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n931), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1115), .A2(new_n814), .A3(new_n888), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1106), .B1(new_n1113), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n924), .A2(G330), .A3(new_n814), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n1098), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n1100), .ZN(new_n1120));
  NOR3_X1   g0920(.A1(new_n1096), .A2(new_n1120), .A3(new_n856), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1098), .B1(new_n721), .B2(new_n815), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1116), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1121), .B1(new_n860), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n463), .A2(new_n1115), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n918), .A2(new_n624), .A3(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1117), .A2(new_n1128), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1106), .B(new_n1127), .C1(new_n1113), .C2(new_n1116), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1129), .A2(new_n686), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n282), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n728), .B1(new_n1132), .B2(new_n823), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n752), .A2(G97), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n767), .A2(G283), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n324), .B1(new_n325), .B2(new_n755), .C1(new_n763), .C2(new_n202), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(G116), .B2(new_n768), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1071), .B1(new_n958), .B2(new_n770), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G107), .B2(new_n833), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1134), .A2(new_n1135), .A3(new_n1137), .A4(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(KEYINPUT54), .B(G143), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n752), .A2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n763), .A2(new_n841), .ZN(new_n1144));
  INV_X1    g0944(.A(G159), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n759), .A2(new_n945), .B1(new_n761), .B2(new_n1145), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n1144), .B(new_n1146), .C1(G125), .C2(new_n830), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n768), .A2(G132), .ZN(new_n1148));
  NOR3_X1   g0948(.A1(new_n755), .A2(KEYINPUT53), .A3(new_n285), .ZN(new_n1149));
  OAI21_X1  g0949(.A(KEYINPUT53), .B1(new_n755), .B2(new_n285), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n266), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1149), .B(new_n1151), .C1(new_n767), .C2(G128), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1143), .A2(new_n1147), .A3(new_n1148), .A4(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1140), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1133), .B1(new_n1154), .B2(new_n743), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n1105), .B2(new_n741), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT117), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1117), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1157), .B1(new_n1158), .B2(new_n727), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1131), .A2(new_n1159), .ZN(G378));
  OAI21_X1  g0960(.A(new_n663), .B1(new_n298), .B2(new_n299), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT119), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n317), .A2(new_n1163), .ZN(new_n1164));
  XOR2_X1   g0964(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1165));
  NAND4_X1  g0965(.A1(new_n306), .A2(new_n315), .A3(new_n316), .A4(new_n1162), .ZN(new_n1166));
  AND3_X1   g0966(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1165), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n930), .A2(new_n1114), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1170), .B(G330), .C1(new_n934), .C2(new_n927), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n917), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n890), .B1(new_n1105), .B2(new_n1101), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1174), .A2(new_n889), .A3(new_n1171), .A4(new_n1169), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT121), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1173), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1172), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1178), .A2(KEYINPUT121), .A3(new_n889), .A4(new_n1174), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1177), .A2(KEYINPUT57), .A3(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1126), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1130), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT120), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1130), .A2(KEYINPUT120), .A3(new_n1181), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1180), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(KEYINPUT122), .B1(new_n1186), .B2(new_n687), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT122), .ZN(new_n1188));
  AND3_X1   g0988(.A1(new_n1130), .A2(KEYINPUT120), .A3(new_n1181), .ZN(new_n1189));
  AOI21_X1  g0989(.A(KEYINPUT120), .B1(new_n1130), .B2(new_n1181), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1188), .B(new_n686), .C1(new_n1191), .C2(new_n1180), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT57), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1187), .A2(new_n1192), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1193), .A2(new_n727), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n728), .B1(G50), .B2(new_n823), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n324), .A2(new_n251), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n1030), .B2(G77), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n944), .B(new_n1201), .C1(new_n835), .C2(new_n224), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n830), .A2(G283), .B1(new_n764), .B2(G58), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1203), .B1(new_n408), .B2(new_n759), .C1(new_n751), .C2(new_n444), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1202), .B(new_n1204), .C1(G116), .C2(new_n767), .ZN(new_n1205));
  XOR2_X1   g1005(.A(new_n1205), .B(KEYINPUT58), .Z(new_n1206));
  OAI211_X1 g1006(.A(new_n1200), .B(new_n841), .C1(G33), .C2(G41), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n784), .A2(G150), .B1(new_n1030), .B2(new_n1142), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(G132), .B2(new_n833), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(G125), .A2(new_n767), .B1(new_n768), .B2(G128), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1210), .B(new_n1211), .C1(new_n751), .C2(new_n945), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1212), .A2(KEYINPUT59), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(KEYINPUT59), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n250), .B(new_n251), .C1(new_n763), .C2(new_n771), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G124), .B2(new_n830), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1206), .B(new_n1207), .C1(new_n1213), .C2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT118), .ZN(new_n1219));
  OR2_X1    g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n822), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1199), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n1170), .B2(new_n741), .ZN(new_n1223));
  AND2_X1   g1023(.A1(new_n1198), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1197), .A2(new_n1224), .ZN(G375));
  OAI22_X1  g1025(.A1(new_n839), .A2(new_n949), .B1(new_n835), .B2(new_n945), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n833), .A2(new_n1142), .B1(new_n784), .B2(G50), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1227), .B(new_n266), .C1(new_n201), .C2(new_n763), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1226), .B(new_n1228), .C1(G150), .C2(new_n752), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n830), .A2(G128), .B1(G159), .B2(new_n1030), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT123), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n324), .B1(new_n408), .B2(new_n755), .C1(new_n763), .C2(new_n222), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n835), .A2(new_n781), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1232), .B(new_n1233), .C1(G294), .C2(new_n767), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1044), .B1(G116), .B2(new_n833), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n777), .B2(new_n770), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(new_n752), .B2(G107), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1229), .A2(new_n1231), .B1(new_n1234), .B2(new_n1237), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n728), .B1(G68), .B2(new_n823), .C1(new_n1238), .C2(new_n822), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(new_n1098), .B2(new_n740), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1124), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1240), .B1(new_n1241), .B2(new_n727), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1128), .A2(new_n1022), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1241), .A2(new_n1181), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1242), .B1(new_n1243), .B2(new_n1244), .ZN(G381));
  INV_X1    g1045(.A(G390), .ZN(new_n1246));
  INV_X1    g1046(.A(G384), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NOR4_X1   g1048(.A1(new_n1248), .A2(G381), .A3(G396), .A4(G393), .ZN(new_n1249));
  INV_X1    g1049(.A(G387), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(G378), .B(KEYINPUT124), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  OR2_X1    g1052(.A1(new_n1252), .A2(G375), .ZN(G407));
  INV_X1    g1053(.A(G213), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1254), .A2(G343), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1251), .A2(new_n1255), .ZN(new_n1256));
  OAI211_X1 g1056(.A(G407), .B(G213), .C1(G375), .C2(new_n1256), .ZN(G409));
  NAND2_X1  g1057(.A1(G387), .A2(new_n1246), .ZN(new_n1258));
  OAI211_X1 g1058(.A(G390), .B(new_n968), .C1(new_n1000), .C2(new_n1023), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(G393), .B(G396), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT125), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n1260), .A2(new_n1261), .A3(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1261), .B1(new_n1260), .B2(new_n1262), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1197), .A2(G378), .A3(new_n1224), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1177), .A2(new_n727), .A3(new_n1179), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1223), .B(new_n1268), .C1(new_n1194), .C2(new_n1021), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1251), .A2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1255), .B1(new_n1267), .B2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT62), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1244), .B1(KEYINPUT60), .B2(new_n1128), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1124), .A2(KEYINPUT60), .A3(new_n1126), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n686), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1242), .B1(new_n1273), .B2(new_n1275), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(new_n1276), .B(G384), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1271), .A2(new_n1272), .A3(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT61), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1255), .A2(G2897), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(new_n1277), .B(new_n1280), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1278), .B(new_n1279), .C1(new_n1271), .C2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1272), .B1(new_n1271), .B2(new_n1277), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1266), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(new_n1263), .A2(new_n1264), .A3(KEYINPUT61), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1285), .B1(new_n1271), .B2(new_n1281), .ZN(new_n1286));
  AOI21_X1  g1086(.A(KEYINPUT63), .B1(new_n1271), .B2(new_n1277), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1267), .A2(new_n1270), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1255), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1277), .A2(KEYINPUT63), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1289), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(KEYINPUT126), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT126), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1271), .A2(new_n1294), .A3(new_n1291), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1293), .A2(new_n1295), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1288), .A2(new_n1296), .A3(KEYINPUT127), .ZN(new_n1297));
  AOI21_X1  g1097(.A(KEYINPUT127), .B1(new_n1288), .B2(new_n1296), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1284), .B1(new_n1297), .B2(new_n1298), .ZN(G405));
  NAND2_X1  g1099(.A1(G375), .A2(new_n1251), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1267), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1301), .B(new_n1277), .ZN(new_n1302));
  XNOR2_X1  g1102(.A(new_n1302), .B(new_n1266), .ZN(G402));
endmodule


