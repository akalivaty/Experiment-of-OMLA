//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 1 0 1 0 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 1 1 0 0 1 1 1 0 1 1 1 0 0 0 0 0 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n626, new_n627, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n793, new_n794, new_n795, new_n797, new_n798, new_n799, new_n800,
    new_n802, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n858, new_n859, new_n860,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914;
  NAND2_X1  g000(.A1(G211gat), .A2(G218gat), .ZN(new_n202));
  INV_X1    g001(.A(G211gat), .ZN(new_n203));
  INV_X1    g002(.A(G218gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT22), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n202), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G197gat), .B(G204gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT76), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n207), .A2(KEYINPUT76), .A3(new_n208), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n208), .A2(KEYINPUT22), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n214), .A2(new_n202), .A3(new_n205), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  XOR2_X1   g016(.A(G155gat), .B(G162gat), .Z(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G155gat), .ZN(new_n220));
  INV_X1    g019(.A(G162gat), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT2), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  XOR2_X1   g021(.A(G141gat), .B(G148gat), .Z(new_n223));
  NAND3_X1  g022(.A1(new_n219), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n222), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(new_n218), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n224), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT29), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n217), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT3), .B1(new_n216), .B2(new_n229), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n224), .A2(new_n226), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n231), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT82), .ZN(new_n236));
  NAND2_X1  g035(.A1(G228gat), .A2(G233gat), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT82), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n231), .B(new_n238), .C1(new_n232), .C2(new_n234), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n236), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n235), .A2(KEYINPUT82), .A3(G228gat), .A4(G233gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n240), .A2(G22gat), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT83), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(G78gat), .B(G106gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT31), .B(G50gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n240), .A2(new_n241), .ZN(new_n249));
  INV_X1    g048(.A(G22gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(new_n242), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n251), .A2(KEYINPUT83), .A3(new_n242), .A4(new_n247), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(G127gat), .A2(G134gat), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(G127gat), .A2(G134gat), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(KEYINPUT70), .A3(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n261));
  INV_X1    g060(.A(new_n259), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n261), .B1(new_n262), .B2(new_n257), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT1), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(G113gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n265), .A2(G120gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT68), .ZN(new_n267));
  INV_X1    g066(.A(G120gat), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n267), .B1(new_n268), .B2(G113gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n265), .A2(KEYINPUT68), .A3(G120gat), .ZN(new_n270));
  AOI211_X1 g069(.A(KEYINPUT69), .B(new_n266), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n269), .A2(new_n270), .ZN(new_n273));
  INV_X1    g072(.A(new_n266), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n264), .B1(new_n271), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT71), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n278), .B(new_n264), .C1(new_n271), .C2(new_n275), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G169gat), .ZN(new_n281));
  INV_X1    g080(.A(G176gat), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n281), .A2(new_n282), .A3(KEYINPUT23), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT23), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n284), .B1(G169gat), .B2(G176gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n283), .B(new_n285), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  AND3_X1   g088(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292));
  NOR3_X1   g091(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT25), .B1(new_n289), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(G183gat), .A2(G190gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT24), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G183gat), .ZN(new_n298));
  INV_X1    g097(.A(G190gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(new_n299), .A3(KEYINPUT64), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT64), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n301), .B1(G183gat), .B2(G190gat), .ZN(new_n302));
  NAND3_X1  g101(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n297), .A2(new_n300), .A3(new_n302), .A4(new_n303), .ZN(new_n304));
  AND2_X1   g103(.A1(new_n283), .A2(new_n285), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT25), .ZN(new_n306));
  INV_X1    g105(.A(new_n288), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(new_n286), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n304), .A2(new_n305), .A3(new_n306), .A4(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT28), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT27), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n312), .A2(G183gat), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n299), .B1(new_n313), .B2(KEYINPUT66), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT66), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n298), .A2(KEYINPUT27), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n312), .A2(G183gat), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n311), .B1(new_n314), .B2(new_n318), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n316), .A2(new_n317), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n320), .A2(KEYINPUT28), .A3(new_n299), .ZN(new_n321));
  AOI22_X1  g120(.A1(new_n319), .A2(new_n321), .B1(G183gat), .B2(G190gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT67), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT26), .ZN(new_n324));
  NOR2_X1   g123(.A1(G169gat), .A2(G176gat), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n308), .B(new_n323), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n324), .ZN(new_n327));
  OAI22_X1  g126(.A1(new_n287), .A2(new_n288), .B1(new_n324), .B2(new_n325), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT67), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n326), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n310), .B1(new_n322), .B2(new_n330), .ZN(new_n331));
  XOR2_X1   g130(.A(G113gat), .B(G120gat), .Z(new_n332));
  INV_X1    g131(.A(KEYINPUT1), .ZN(new_n333));
  AOI211_X1 g132(.A(new_n257), .B(new_n262), .C1(new_n332), .C2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n280), .A2(new_n331), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT72), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n280), .A2(new_n335), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n330), .ZN(new_n339));
  INV_X1    g138(.A(new_n310), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n334), .B1(new_n277), .B2(new_n279), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT72), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n343), .A2(new_n344), .A3(new_n331), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n337), .A2(new_n342), .A3(new_n345), .ZN(new_n346));
  AND2_X1   g145(.A1(G227gat), .A2(G233gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G15gat), .B(G43gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n349), .B(G71gat), .ZN(new_n350));
  INV_X1    g149(.A(G99gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n350), .B(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(KEYINPUT33), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n348), .A2(KEYINPUT32), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT74), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT32), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n356), .B1(new_n346), .B2(new_n347), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT74), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n357), .A2(new_n358), .A3(new_n353), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT33), .B1(new_n346), .B2(new_n347), .ZN(new_n361));
  INV_X1    g160(.A(new_n352), .ZN(new_n362));
  NOR4_X1   g161(.A1(new_n361), .A2(new_n357), .A3(KEYINPUT73), .A4(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT73), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n362), .B1(new_n348), .B2(KEYINPUT32), .ZN(new_n365));
  INV_X1    g164(.A(new_n361), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n360), .B1(new_n363), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n346), .A2(new_n347), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n369), .B(KEYINPUT34), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT75), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n370), .B(new_n360), .C1(new_n363), .C2(new_n367), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n368), .A2(KEYINPUT75), .A3(new_n371), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n256), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT0), .B(G57gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n378), .B(G85gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(G1gat), .B(G29gat), .ZN(new_n380));
  XOR2_X1   g179(.A(new_n379), .B(new_n380), .Z(new_n381));
  NAND2_X1  g180(.A1(G225gat), .A2(G233gat), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n343), .A2(new_n234), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n343), .A2(new_n234), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n383), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n384), .A2(new_n382), .ZN(new_n388));
  AND2_X1   g187(.A1(new_n388), .A2(KEYINPUT4), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n233), .A2(KEYINPUT3), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n228), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT4), .B1(new_n343), .B2(new_n391), .ZN(new_n392));
  AND2_X1   g191(.A1(new_n392), .A2(new_n384), .ZN(new_n393));
  OAI211_X1 g192(.A(KEYINPUT5), .B(new_n387), .C1(new_n389), .C2(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT79), .B(KEYINPUT4), .ZN(new_n395));
  OR2_X1    g194(.A1(new_n384), .A2(new_n395), .ZN(new_n396));
  OR2_X1    g195(.A1(new_n343), .A2(new_n391), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n384), .A2(new_n395), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n383), .A2(KEYINPUT5), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n396), .A2(new_n397), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n381), .B1(new_n394), .B2(new_n400), .ZN(new_n401));
  XOR2_X1   g200(.A(KEYINPUT80), .B(KEYINPUT6), .Z(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n394), .A2(new_n400), .ZN(new_n404));
  INV_X1    g203(.A(new_n381), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n387), .A2(KEYINPUT5), .ZN(new_n407));
  AOI22_X1  g206(.A1(new_n388), .A2(KEYINPUT4), .B1(new_n392), .B2(new_n384), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n381), .B(new_n400), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n402), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(KEYINPUT81), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n406), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT81), .B1(new_n409), .B2(new_n410), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n403), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(G226gat), .A2(G233gat), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n415), .B1(new_n331), .B2(KEYINPUT29), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n341), .A2(G226gat), .A3(G233gat), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n417), .A2(KEYINPUT78), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n417), .A2(KEYINPUT78), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n216), .B(new_n416), .C1(new_n418), .C2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n417), .A2(KEYINPUT77), .ZN(new_n421));
  OR3_X1    g220(.A1(new_n331), .A2(KEYINPUT77), .A3(new_n415), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(new_n416), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n217), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  XOR2_X1   g224(.A(G8gat), .B(G36gat), .Z(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(G64gat), .ZN(new_n427));
  XOR2_X1   g226(.A(new_n427), .B(G92gat), .Z(new_n428));
  NAND2_X1  g227(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n428), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n420), .A2(new_n424), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n429), .A2(KEYINPUT30), .A3(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n425), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT30), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n433), .A2(new_n434), .A3(new_n430), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n414), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n377), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT35), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT87), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n365), .A2(new_n366), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT73), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n365), .A2(new_n364), .A3(new_n366), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n370), .B1(new_n445), .B2(new_n360), .ZN(new_n446));
  INV_X1    g245(.A(new_n374), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n441), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n372), .A2(KEYINPUT87), .A3(new_n374), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT86), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n406), .A2(new_n450), .A3(new_n410), .A4(new_n409), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n409), .A2(new_n410), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT86), .B1(new_n452), .B2(new_n401), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n451), .A2(new_n403), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT35), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n255), .A2(new_n455), .A3(new_n436), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n448), .A2(new_n449), .A3(new_n454), .A4(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT88), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n457), .A2(new_n458), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n440), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n375), .A2(KEYINPUT36), .A3(new_n376), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n253), .A2(KEYINPUT84), .A3(new_n254), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT84), .B1(new_n253), .B2(new_n254), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(new_n437), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT36), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n372), .A2(new_n467), .A3(new_n374), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n462), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT85), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n451), .A2(new_n403), .A3(new_n453), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT37), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n430), .B1(new_n433), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n473), .B1(new_n472), .B2(new_n433), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT38), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT38), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n423), .A2(new_n216), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n416), .B1(new_n418), .B2(new_n419), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n477), .B(KEYINPUT37), .C1(new_n478), .C2(new_n216), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n473), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n471), .A2(new_n431), .A3(new_n475), .A4(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT40), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n383), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n484), .B(KEYINPUT39), .C1(new_n388), .C2(new_n386), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n485), .B(new_n381), .C1(KEYINPUT39), .C2(new_n484), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n436), .B1(new_n482), .B2(new_n486), .ZN(new_n487));
  OR2_X1    g286(.A1(new_n486), .A2(new_n482), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(new_n406), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n481), .A2(new_n489), .A3(new_n255), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT85), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n462), .A2(new_n466), .A3(new_n491), .A4(new_n468), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n470), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n461), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(G15gat), .B(G22gat), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT16), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n495), .B1(new_n496), .B2(G1gat), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n497), .B1(G1gat), .B2(new_n495), .ZN(new_n498));
  OR2_X1    g297(.A1(new_n498), .A2(G8gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(G8gat), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(G57gat), .B(G64gat), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n504));
  OR2_X1    g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(G71gat), .B(G78gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n505), .B(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n502), .B1(KEYINPUT21), .B2(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n508), .B(new_n298), .ZN(new_n509));
  AND2_X1   g308(.A1(G231gat), .A2(G233gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n509), .B(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(KEYINPUT92), .B(KEYINPUT93), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n507), .A2(KEYINPUT21), .ZN(new_n514));
  XNOR2_X1  g313(.A(G127gat), .B(G155gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(G211gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n514), .B(new_n516), .ZN(new_n517));
  XOR2_X1   g316(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n513), .B(new_n519), .ZN(new_n520));
  OR3_X1    g319(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n522));
  AOI22_X1  g321(.A1(new_n521), .A2(new_n522), .B1(G29gat), .B2(G36gat), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT15), .ZN(new_n524));
  XOR2_X1   g323(.A(G43gat), .B(G50gat), .Z(new_n525));
  OR3_X1    g324(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n525), .A2(new_n524), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(new_n524), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n527), .A2(new_n528), .A3(new_n523), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT90), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT17), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G85gat), .A2(G92gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT8), .ZN(new_n536));
  AND2_X1   g335(.A1(G99gat), .A2(G106gat), .ZN(new_n537));
  OAI221_X1 g336(.A(new_n535), .B1(new_n536), .B2(new_n537), .C1(G85gat), .C2(G92gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(G99gat), .B(G106gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n533), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n540), .A2(new_n530), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT41), .ZN(new_n544));
  NAND2_X1  g343(.A1(G232gat), .A2(G233gat), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n542), .B(new_n543), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n544), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  XOR2_X1   g347(.A(G190gat), .B(G218gat), .Z(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(KEYINPUT95), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n548), .B(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(KEYINPUT94), .B(G134gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(G162gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n551), .B(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n520), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n507), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n540), .B(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT10), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n541), .A2(new_n556), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT10), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G230gat), .A2(G233gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n563), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n540), .A2(new_n507), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n566), .B1(new_n560), .B2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT96), .ZN(new_n569));
  XNOR2_X1  g368(.A(G120gat), .B(G148gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G204gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT97), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(new_n282), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  OR3_X1    g373(.A1(new_n565), .A2(new_n569), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(KEYINPUT98), .B1(new_n562), .B2(new_n563), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT98), .ZN(new_n577));
  AOI211_X1 g376(.A(new_n577), .B(new_n566), .C1(new_n559), .C2(new_n561), .ZN(new_n578));
  NOR3_X1   g377(.A1(new_n569), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n575), .B1(new_n579), .B2(new_n573), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n533), .A2(new_n501), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n502), .A2(new_n530), .ZN(new_n583));
  NAND2_X1  g382(.A1(G229gat), .A2(G233gat), .ZN(new_n584));
  AND3_X1   g383(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  OR2_X1    g384(.A1(new_n585), .A2(KEYINPUT18), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n501), .B(new_n530), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n584), .B(KEYINPUT91), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT13), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n585), .A2(KEYINPUT18), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n586), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G113gat), .B(G141gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(G169gat), .B(G197gat), .Z(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(KEYINPUT12), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n593), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n586), .A2(new_n591), .A3(new_n592), .A4(new_n599), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n581), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n555), .A2(new_n604), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n494), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n414), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(KEYINPUT99), .B(G1gat), .Z(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(G1324gat));
  INV_X1    g409(.A(new_n606), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n611), .A2(new_n436), .ZN(new_n612));
  NAND2_X1  g411(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n613));
  INV_X1    g412(.A(G8gat), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n496), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n612), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT42), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n617), .B1(new_n614), .B2(new_n612), .ZN(G1325gat));
  AND3_X1   g417(.A1(new_n372), .A2(KEYINPUT87), .A3(new_n374), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT87), .B1(new_n372), .B2(new_n374), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(G15gat), .B1(new_n606), .B2(new_n621), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n462), .A2(new_n468), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n611), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n622), .B1(new_n624), .B2(G15gat), .ZN(G1326gat));
  NAND2_X1  g424(.A1(new_n606), .A2(new_n465), .ZN(new_n626));
  XNOR2_X1  g425(.A(KEYINPUT43), .B(G22gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(G1327gat));
  AOI21_X1  g427(.A(new_n554), .B1(new_n461), .B2(new_n493), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n520), .A2(new_n604), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR3_X1   g430(.A1(new_n631), .A2(G29gat), .A3(new_n414), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n632), .B(KEYINPUT45), .Z(new_n633));
  INV_X1    g432(.A(KEYINPUT44), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n551), .B(new_n553), .Z(new_n635));
  AOI21_X1  g434(.A(new_n455), .B1(new_n377), .B2(new_n438), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n621), .A2(KEYINPUT88), .A3(new_n454), .A4(new_n456), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n457), .A2(new_n458), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AND4_X1   g438(.A1(new_n490), .A2(new_n466), .A3(new_n462), .A4(new_n468), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n634), .B(new_n635), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  OAI211_X1 g440(.A(KEYINPUT100), .B(new_n641), .C1(new_n629), .C2(new_n634), .ZN(new_n642));
  AND3_X1   g441(.A1(new_n470), .A2(new_n490), .A3(new_n492), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n635), .B1(new_n643), .B2(new_n639), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT100), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n644), .A2(new_n645), .A3(KEYINPUT44), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n630), .ZN(new_n648));
  OAI21_X1  g447(.A(G29gat), .B1(new_n648), .B2(new_n414), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n649), .ZN(G1328gat));
  OAI21_X1  g449(.A(G36gat), .B1(new_n648), .B2(new_n436), .ZN(new_n651));
  NOR3_X1   g450(.A1(new_n631), .A2(G36gat), .A3(new_n436), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT46), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(G1329gat));
  INV_X1    g453(.A(new_n623), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n647), .A2(new_n655), .A3(new_n630), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(G43gat), .ZN(new_n657));
  INV_X1    g456(.A(new_n621), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n658), .A2(G43gat), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n629), .A2(new_n630), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n657), .A2(KEYINPUT47), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(KEYINPUT101), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n657), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT47), .ZN(new_n665));
  AOI21_X1  g464(.A(KEYINPUT102), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n662), .B1(new_n656), .B2(G43gat), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT102), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n667), .A2(new_n668), .A3(KEYINPUT47), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n661), .B1(new_n666), .B2(new_n669), .ZN(G1330gat));
  INV_X1    g469(.A(new_n648), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n256), .ZN(new_n672));
  AND3_X1   g471(.A1(new_n672), .A2(KEYINPUT48), .A3(G50gat), .ZN(new_n673));
  INV_X1    g472(.A(new_n465), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n631), .A2(G50gat), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n676), .B1(KEYINPUT103), .B2(KEYINPUT48), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n676), .A2(KEYINPUT103), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n671), .A2(new_n465), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n678), .B1(new_n679), .B2(G50gat), .ZN(new_n680));
  OAI22_X1  g479(.A1(new_n673), .A2(new_n677), .B1(new_n680), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g480(.A1(new_n623), .A2(new_n490), .A3(new_n466), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n581), .B1(new_n461), .B2(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n555), .A2(new_n603), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n685), .A2(new_n414), .ZN(new_n686));
  XOR2_X1   g485(.A(KEYINPUT104), .B(G57gat), .Z(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1332gat));
  NOR2_X1   g487(.A1(new_n685), .A2(new_n436), .ZN(new_n689));
  NOR2_X1   g488(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n690));
  AND2_X1   g489(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n689), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n692), .B1(new_n689), .B2(new_n690), .ZN(G1333gat));
  OAI21_X1  g492(.A(G71gat), .B1(new_n685), .B2(new_n623), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n683), .A2(new_n621), .A3(new_n684), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n694), .B1(G71gat), .B2(new_n695), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT105), .B(KEYINPUT50), .Z(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1334gat));
  NOR2_X1   g497(.A1(new_n685), .A2(new_n674), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n699), .B(G78gat), .Z(G1335gat));
  NOR3_X1   g499(.A1(new_n520), .A2(new_n581), .A3(new_n603), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n647), .A2(new_n701), .ZN(new_n702));
  OR3_X1    g501(.A1(new_n702), .A2(KEYINPUT106), .A3(new_n414), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT106), .B1(new_n702), .B2(new_n414), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(G85gat), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n461), .A2(new_n682), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n520), .A2(new_n603), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n706), .A2(KEYINPUT51), .A3(new_n635), .A4(new_n707), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n635), .B(new_n707), .C1(new_n639), .C2(new_n640), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT51), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n581), .B1(new_n708), .B2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(G85gat), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n712), .A2(new_n713), .A3(new_n607), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n705), .A2(new_n714), .ZN(G1336gat));
  OR2_X1    g514(.A1(new_n702), .A2(new_n436), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(G92gat), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n436), .A2(G92gat), .ZN(new_n718));
  AOI21_X1  g517(.A(KEYINPUT52), .B1(new_n712), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(KEYINPUT108), .B1(new_n709), .B2(KEYINPUT107), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT107), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT108), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(new_n723), .B2(new_n710), .ZN(new_n724));
  AOI22_X1  g523(.A1(new_n721), .A2(new_n710), .B1(new_n709), .B2(new_n724), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n725), .A2(new_n580), .ZN(new_n726));
  AOI22_X1  g525(.A1(new_n716), .A2(G92gat), .B1(new_n718), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT52), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n720), .B1(new_n727), .B2(new_n728), .ZN(G1337gat));
  OAI21_X1  g528(.A(G99gat), .B1(new_n702), .B2(new_n623), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n712), .A2(new_n351), .A3(new_n621), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(G1338gat));
  NAND4_X1  g531(.A1(new_n642), .A2(new_n646), .A3(new_n465), .A4(new_n701), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(G106gat), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n581), .A2(G106gat), .A3(new_n255), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n725), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(KEYINPUT53), .ZN(new_n738));
  INV_X1    g537(.A(new_n735), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n739), .B1(new_n708), .B2(new_n711), .ZN(new_n740));
  AND2_X1   g539(.A1(KEYINPUT109), .A2(KEYINPUT53), .ZN(new_n741));
  NOR2_X1   g540(.A1(KEYINPUT109), .A2(KEYINPUT53), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n642), .A2(new_n646), .A3(new_n256), .A4(new_n701), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(G106gat), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT110), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n743), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n746), .B1(new_n743), .B2(new_n745), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n738), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT111), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n738), .B(KEYINPUT111), .C1(new_n747), .C2(new_n748), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(G1339gat));
  INV_X1    g552(.A(KEYINPUT54), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n576), .B2(new_n578), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n559), .A2(new_n566), .A3(new_n561), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n564), .A2(KEYINPUT54), .A3(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n755), .A2(new_n574), .A3(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT55), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT112), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n755), .A2(new_n757), .A3(KEYINPUT55), .A4(new_n574), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n575), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n761), .A2(new_n603), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n584), .B1(new_n582), .B2(new_n583), .ZN(new_n766));
  OR2_X1    g565(.A1(new_n766), .A2(KEYINPUT113), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n587), .A2(new_n590), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n766), .A2(KEYINPUT113), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n598), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n580), .A2(new_n602), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n765), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n554), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n771), .A2(new_n602), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n761), .A2(new_n764), .A3(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n776), .A2(new_n554), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n520), .B1(new_n774), .B2(new_n778), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n555), .A2(new_n580), .A3(new_n603), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n781), .A2(new_n658), .A3(new_n465), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n607), .A2(new_n436), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n603), .ZN(new_n786));
  OAI21_X1  g585(.A(G113gat), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n781), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n788), .A2(new_n377), .A3(new_n784), .ZN(new_n789));
  XOR2_X1   g588(.A(new_n789), .B(KEYINPUT114), .Z(new_n790));
  NAND2_X1  g589(.A1(new_n603), .A2(new_n265), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n787), .B1(new_n790), .B2(new_n791), .ZN(G1340gat));
  OAI21_X1  g591(.A(G120gat), .B1(new_n785), .B2(new_n581), .ZN(new_n793));
  XOR2_X1   g592(.A(new_n793), .B(KEYINPUT115), .Z(new_n794));
  NAND2_X1  g593(.A1(new_n580), .A2(new_n268), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n794), .B1(new_n790), .B2(new_n795), .ZN(G1341gat));
  INV_X1    g595(.A(G127gat), .ZN(new_n797));
  INV_X1    g596(.A(new_n520), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n785), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(G127gat), .B1(new_n789), .B2(new_n520), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n799), .A2(new_n800), .ZN(G1342gat));
  INV_X1    g600(.A(G134gat), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n789), .A2(new_n802), .A3(new_n635), .ZN(new_n803));
  XOR2_X1   g602(.A(new_n803), .B(KEYINPUT56), .Z(new_n804));
  OAI21_X1  g603(.A(G134gat), .B1(new_n785), .B2(new_n554), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(G1343gat));
  INV_X1    g605(.A(KEYINPUT119), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n655), .A2(new_n783), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n781), .A2(new_n255), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT57), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT117), .ZN(new_n813));
  INV_X1    g612(.A(new_n760), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n814), .B2(new_n763), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n764), .A2(KEYINPUT117), .A3(new_n760), .ZN(new_n816));
  AND3_X1   g615(.A1(new_n815), .A2(new_n816), .A3(new_n603), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n772), .B(KEYINPUT116), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n554), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n778), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n780), .B1(new_n820), .B2(new_n798), .ZN(new_n821));
  OAI21_X1  g620(.A(KEYINPUT57), .B1(new_n821), .B2(new_n674), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n812), .A2(new_n603), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n807), .B1(new_n823), .B2(G141gat), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n810), .A2(new_n808), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n786), .A2(G141gat), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(KEYINPUT118), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n828), .B1(new_n823), .B2(G141gat), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n824), .A2(new_n829), .A3(KEYINPUT58), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT58), .ZN(new_n831));
  AOI221_X4 g630(.A(new_n828), .B1(new_n807), .B2(new_n831), .C1(new_n823), .C2(G141gat), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n830), .A2(new_n832), .ZN(G1344gat));
  AND2_X1   g632(.A1(new_n812), .A2(new_n822), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n580), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT59), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n835), .A2(new_n836), .A3(G148gat), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT120), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n838), .B(new_n811), .C1(new_n821), .C2(new_n674), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT116), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n772), .B(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n815), .A2(new_n816), .A3(new_n603), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n635), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n798), .B1(new_n843), .B2(new_n777), .ZN(new_n844));
  INV_X1    g643(.A(new_n780), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n674), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(KEYINPUT120), .B1(new_n846), .B2(KEYINPUT57), .ZN(new_n847));
  OAI211_X1 g646(.A(KEYINPUT57), .B(new_n256), .C1(new_n779), .C2(new_n780), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n839), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n849), .A2(new_n580), .A3(new_n808), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(G148gat), .ZN(new_n851));
  AOI21_X1  g650(.A(KEYINPUT121), .B1(new_n851), .B2(KEYINPUT59), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT121), .ZN(new_n853));
  AOI211_X1 g652(.A(new_n853), .B(new_n836), .C1(new_n850), .C2(G148gat), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n837), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  OR3_X1    g654(.A1(new_n825), .A2(G148gat), .A3(new_n581), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(G1345gat));
  INV_X1    g656(.A(new_n825), .ZN(new_n858));
  AOI21_X1  g657(.A(G155gat), .B1(new_n858), .B2(new_n520), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n834), .A2(new_n520), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n859), .B1(new_n860), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g660(.A(new_n221), .B1(new_n834), .B2(new_n635), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n825), .A2(G162gat), .A3(new_n554), .ZN(new_n863));
  OR3_X1    g662(.A1(new_n862), .A2(KEYINPUT122), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT122), .B1(new_n862), .B2(new_n863), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(G1347gat));
  NOR2_X1   g665(.A1(new_n607), .A2(new_n436), .ZN(new_n867));
  AND3_X1   g666(.A1(new_n788), .A2(new_n377), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n868), .A2(new_n281), .A3(new_n603), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n869), .B(KEYINPUT123), .ZN(new_n870));
  AND4_X1   g669(.A1(new_n621), .A2(new_n788), .A3(new_n674), .A4(new_n867), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(G169gat), .B1(new_n872), .B2(new_n786), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n870), .A2(new_n873), .ZN(G1348gat));
  AOI21_X1  g673(.A(G176gat), .B1(new_n868), .B2(new_n580), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n872), .A2(new_n581), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n875), .B1(new_n876), .B2(G176gat), .ZN(G1349gat));
  AOI21_X1  g676(.A(new_n298), .B1(new_n871), .B2(new_n520), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n520), .A2(new_n320), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n878), .B1(new_n868), .B2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT60), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n880), .B(new_n881), .ZN(G1350gat));
  NAND3_X1  g681(.A1(new_n868), .A2(new_n299), .A3(new_n635), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT61), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n871), .A2(new_n635), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n884), .B1(new_n885), .B2(G190gat), .ZN(new_n886));
  AOI211_X1 g685(.A(KEYINPUT61), .B(new_n299), .C1(new_n871), .C2(new_n635), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n883), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT124), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT124), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n890), .B(new_n883), .C1(new_n886), .C2(new_n887), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(G1351gat));
  AND2_X1   g691(.A1(new_n623), .A2(new_n867), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n849), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(G197gat), .B1(new_n894), .B2(new_n786), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n810), .A2(new_n893), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n896), .A2(G197gat), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n895), .B1(new_n786), .B2(new_n897), .ZN(G1352gat));
  NOR3_X1   g697(.A1(new_n896), .A2(G204gat), .A3(new_n581), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n899), .B(KEYINPUT62), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n849), .A2(new_n580), .A3(new_n893), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(G204gat), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(new_n902), .ZN(G1353gat));
  OAI21_X1  g702(.A(G211gat), .B1(new_n894), .B2(new_n798), .ZN(new_n904));
  NAND2_X1  g703(.A1(KEYINPUT125), .A2(KEYINPUT63), .ZN(new_n905));
  OR2_X1    g704(.A1(KEYINPUT125), .A2(KEYINPUT63), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(new_n896), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(new_n203), .A3(new_n520), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n907), .B(new_n909), .C1(new_n904), .C2(new_n906), .ZN(G1354gat));
  AOI21_X1  g709(.A(G218gat), .B1(new_n908), .B2(new_n635), .ZN(new_n911));
  XOR2_X1   g710(.A(new_n894), .B(KEYINPUT126), .Z(new_n912));
  NOR2_X1   g711(.A1(new_n554), .A2(new_n204), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT127), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n911), .B1(new_n912), .B2(new_n914), .ZN(G1355gat));
endmodule


