//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 1 1 0 0 1 1 1 1 1 0 0 1 0 0 0 0 0 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 0 0 0 0 1 0 1 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n622, new_n623,
    new_n624, new_n625, new_n627, new_n628, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n781, new_n782, new_n783, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n841, new_n842, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893;
  NOR2_X1   g000(.A1(G57gat), .A2(G64gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G71gat), .A2(G78gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT9), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  AOI21_X1  g004(.A(new_n202), .B1(new_n205), .B2(KEYINPUT90), .ZN(new_n206));
  NAND2_X1  g005(.A1(G57gat), .A2(G64gat), .ZN(new_n207));
  OAI211_X1 g006(.A(new_n206), .B(new_n207), .C1(KEYINPUT90), .C2(new_n205), .ZN(new_n208));
  INV_X1    g007(.A(new_n203), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n209), .A2(KEYINPUT89), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(G71gat), .A2(G78gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n208), .B(new_n210), .C1(new_n209), .C2(new_n212), .ZN(new_n215));
  NAND2_X1  g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216));
  INV_X1    g015(.A(G85gat), .ZN(new_n217));
  INV_X1    g016(.A(G92gat), .ZN(new_n218));
  AOI22_X1  g017(.A1(KEYINPUT8), .A2(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(new_n217), .B2(new_n218), .ZN(new_n221));
  NAND4_X1  g020(.A1(KEYINPUT94), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n219), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  XOR2_X1   g022(.A(G99gat), .B(G106gat), .Z(new_n224));
  XOR2_X1   g023(.A(new_n223), .B(new_n224), .Z(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n214), .A2(new_n215), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT10), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n214), .A2(new_n215), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(new_n225), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n227), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n231), .B1(new_n228), .B2(new_n230), .ZN(new_n232));
  NAND2_X1  g031(.A1(G230gat), .A2(G233gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n227), .A2(new_n230), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n235), .A2(G230gat), .A3(G233gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(G120gat), .B(G148gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(G176gat), .B(G204gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n234), .A2(new_n236), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT98), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n241), .B(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n234), .A2(new_n236), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(new_n239), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G15gat), .B(G22gat), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT16), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n248), .B1(new_n249), .B2(G1gat), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n250), .B1(G1gat), .B2(new_n248), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(G8gat), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(G43gat), .B(G50gat), .Z(new_n254));
  NOR2_X1   g053(.A1(G29gat), .A2(G36gat), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT14), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(G29gat), .A2(G36gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n254), .B1(new_n259), .B2(KEYINPUT15), .ZN(new_n260));
  INV_X1    g059(.A(G43gat), .ZN(new_n261));
  OR2_X1    g060(.A1(new_n261), .A2(G50gat), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT15), .B1(new_n262), .B2(KEYINPUT87), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  XOR2_X1   g063(.A(new_n258), .B(KEYINPUT88), .Z(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(new_n257), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n260), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n254), .B1(new_n266), .B2(new_n263), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n267), .A2(KEYINPUT17), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT17), .B1(new_n267), .B2(new_n268), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n253), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n252), .A2(new_n268), .A3(new_n267), .ZN(new_n272));
  NAND2_X1  g071(.A1(G229gat), .A2(G233gat), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT18), .ZN(new_n275));
  OR2_X1    g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n267), .A2(new_n268), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(new_n253), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(new_n272), .ZN(new_n279));
  XOR2_X1   g078(.A(new_n273), .B(KEYINPUT13), .Z(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n274), .A2(new_n275), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n276), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G113gat), .B(G141gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(G197gat), .ZN(new_n285));
  XOR2_X1   g084(.A(KEYINPUT11), .B(G169gat), .Z(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(KEYINPUT12), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n276), .A2(new_n288), .A3(new_n281), .A4(new_n282), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n247), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n252), .B1(new_n229), .B2(KEYINPUT21), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n294), .B(KEYINPUT93), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n229), .A2(KEYINPUT21), .ZN(new_n296));
  XOR2_X1   g095(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n295), .B(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G127gat), .B(G155gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  XOR2_X1   g100(.A(G183gat), .B(G211gat), .Z(new_n302));
  NAND2_X1  g101(.A1(G231gat), .A2(G233gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(KEYINPUT91), .B(KEYINPUT92), .ZN(new_n305));
  XOR2_X1   g104(.A(new_n304), .B(new_n305), .Z(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  OR2_X1    g106(.A1(new_n301), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n301), .A2(new_n307), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n226), .B1(new_n269), .B2(new_n270), .ZN(new_n311));
  OR2_X1    g110(.A1(new_n311), .A2(KEYINPUT95), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n267), .A2(new_n225), .A3(new_n268), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT41), .ZN(new_n314));
  INV_X1    g113(.A(G232gat), .ZN(new_n315));
  INV_X1    g114(.A(G233gat), .ZN(new_n316));
  NOR3_X1   g115(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n317), .B1(new_n311), .B2(KEYINPUT95), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n312), .A2(new_n313), .A3(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(G190gat), .B(G218gat), .ZN(new_n320));
  XOR2_X1   g119(.A(new_n320), .B(KEYINPUT96), .Z(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n312), .A2(new_n318), .A3(new_n313), .A4(new_n321), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT97), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT97), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n323), .A2(new_n327), .A3(new_n324), .ZN(new_n328));
  XNOR2_X1  g127(.A(G134gat), .B(G162gat), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n314), .B1(new_n315), .B2(new_n316), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n329), .B(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n326), .A2(new_n328), .A3(new_n331), .ZN(new_n332));
  OR2_X1    g131(.A1(new_n328), .A2(new_n331), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n310), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(G183gat), .A2(G190gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NOR2_X1   g136(.A1(G183gat), .A2(G190gat), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT24), .ZN(new_n339));
  NOR3_X1   g138(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(G169gat), .ZN(new_n341));
  INV_X1    g140(.A(G176gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n341), .A2(new_n342), .A3(KEYINPUT23), .ZN(new_n343));
  NAND2_X1  g142(.A1(G169gat), .A2(G176gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g144(.A1(G169gat), .A2(G176gat), .ZN(new_n346));
  OAI22_X1  g145(.A1(new_n346), .A2(KEYINPUT23), .B1(new_n336), .B2(KEYINPUT24), .ZN(new_n347));
  NOR3_X1   g146(.A1(new_n340), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(KEYINPUT64), .B1(new_n348), .B2(KEYINPUT25), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n340), .A2(new_n347), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT25), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n351), .B1(new_n345), .B2(KEYINPUT65), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n350), .B(new_n352), .C1(KEYINPUT65), .C2(new_n345), .ZN(new_n353));
  AND2_X1   g152(.A1(G169gat), .A2(G176gat), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n354), .B1(KEYINPUT23), .B2(new_n346), .ZN(new_n355));
  INV_X1    g154(.A(G183gat), .ZN(new_n356));
  INV_X1    g155(.A(G190gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n358), .A2(KEYINPUT24), .A3(new_n336), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT23), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n360), .B1(G169gat), .B2(G176gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n337), .A2(new_n339), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n355), .A2(new_n359), .A3(new_n361), .A4(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT64), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n363), .A2(new_n364), .A3(new_n351), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n349), .A2(new_n353), .A3(new_n365), .ZN(new_n366));
  NOR3_X1   g165(.A1(new_n354), .A2(new_n346), .A3(KEYINPUT26), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n367), .B1(KEYINPUT26), .B2(new_n346), .ZN(new_n368));
  XOR2_X1   g167(.A(KEYINPUT27), .B(G183gat), .Z(new_n369));
  OAI21_X1  g168(.A(KEYINPUT28), .B1(new_n369), .B2(G190gat), .ZN(new_n370));
  OR3_X1    g169(.A1(new_n356), .A2(KEYINPUT66), .A3(KEYINPUT27), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT28), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT27), .B1(new_n356), .B2(KEYINPUT66), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n371), .A2(new_n372), .A3(new_n357), .A4(new_n373), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n368), .A2(new_n336), .A3(new_n370), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n366), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT68), .B(G120gat), .ZN(new_n377));
  INV_X1    g176(.A(G113gat), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT69), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(G120gat), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT69), .ZN(new_n381));
  INV_X1    g180(.A(G120gat), .ZN(new_n382));
  AND2_X1   g181(.A1(new_n382), .A2(KEYINPUT68), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n382), .A2(KEYINPUT68), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n381), .B(G113gat), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n379), .A2(new_n380), .A3(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT1), .ZN(new_n387));
  XNOR2_X1  g186(.A(G127gat), .B(G134gat), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT70), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(KEYINPUT67), .ZN(new_n391));
  INV_X1    g190(.A(G134gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(G127gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(G113gat), .B(G120gat), .ZN(new_n394));
  OAI221_X1 g193(.A(new_n391), .B1(KEYINPUT67), .B2(new_n393), .C1(KEYINPUT1), .C2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n389), .A2(new_n390), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n390), .B1(new_n389), .B2(new_n395), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n376), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n389), .A2(new_n395), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT70), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n401), .A2(new_n396), .A3(new_n375), .A4(new_n366), .ZN(new_n402));
  INV_X1    g201(.A(G227gat), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n403), .A2(new_n316), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n399), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT33), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT71), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(G15gat), .B(G43gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(G71gat), .B(G99gat), .ZN(new_n411));
  XOR2_X1   g210(.A(new_n410), .B(new_n411), .Z(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n413), .B1(new_n405), .B2(KEYINPUT32), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n405), .A2(KEYINPUT71), .A3(new_n406), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n409), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n412), .A2(KEYINPUT33), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n405), .A2(KEYINPUT32), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT72), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OR2_X1    g219(.A1(new_n418), .A2(new_n419), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n416), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n399), .A2(new_n402), .ZN(new_n423));
  INV_X1    g222(.A(new_n404), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT34), .B1(new_n425), .B2(KEYINPUT73), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT73), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n423), .A2(new_n427), .A3(new_n424), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n423), .A2(new_n427), .A3(KEYINPUT34), .A4(new_n424), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n422), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n418), .B(KEYINPUT72), .ZN(new_n433));
  AOI22_X1  g232(.A1(new_n433), .A2(new_n416), .B1(new_n430), .B2(new_n429), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(G197gat), .B(G204gat), .ZN(new_n436));
  INV_X1    g235(.A(G211gat), .ZN(new_n437));
  INV_X1    g236(.A(G218gat), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n436), .B1(KEYINPUT22), .B2(new_n439), .ZN(new_n440));
  XOR2_X1   g239(.A(G211gat), .B(G218gat), .Z(new_n441));
  XNOR2_X1  g240(.A(new_n440), .B(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(G141gat), .B(G148gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT78), .B(G162gat), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(G155gat), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n443), .B1(new_n445), .B2(KEYINPUT2), .ZN(new_n446));
  AND2_X1   g245(.A1(G155gat), .A2(G162gat), .ZN(new_n447));
  NOR2_X1   g246(.A1(G155gat), .A2(G162gat), .ZN(new_n448));
  OR2_X1    g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n443), .A2(KEYINPUT2), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n450), .A2(new_n447), .ZN(new_n451));
  XOR2_X1   g250(.A(new_n448), .B(KEYINPUT77), .Z(new_n452));
  AOI22_X1  g251(.A1(new_n446), .A2(new_n449), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT3), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT29), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n442), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n456), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n453), .B1(new_n458), .B2(new_n454), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n460), .B(G22gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(G228gat), .A2(G233gat), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT84), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n462), .B1(new_n457), .B2(new_n463), .ZN(new_n464));
  OR2_X1    g263(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n461), .A2(new_n464), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  XOR2_X1   g266(.A(G78gat), .B(G106gat), .Z(new_n468));
  XNOR2_X1  g267(.A(new_n468), .B(KEYINPUT31), .ZN(new_n469));
  XOR2_X1   g268(.A(KEYINPUT83), .B(G50gat), .Z(new_n470));
  XNOR2_X1  g269(.A(new_n469), .B(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n471), .B(KEYINPUT85), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT85), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n465), .A2(new_n474), .A3(new_n471), .A4(new_n466), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n435), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(G226gat), .A2(G233gat), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n376), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n376), .A2(new_n456), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT74), .B1(new_n481), .B2(new_n478), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT29), .B1(new_n366), .B2(new_n375), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT74), .ZN(new_n484));
  NOR3_X1   g283(.A1(new_n483), .A2(new_n484), .A3(new_n479), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n480), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n442), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n486), .A2(KEYINPUT75), .A3(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT75), .ZN(new_n489));
  INV_X1    g288(.A(new_n480), .ZN(new_n490));
  INV_X1    g289(.A(new_n375), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n363), .A2(new_n364), .A3(new_n351), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n364), .B1(new_n363), .B2(new_n351), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n491), .B1(new_n494), .B2(new_n353), .ZN(new_n495));
  OAI211_X1 g294(.A(KEYINPUT74), .B(new_n478), .C1(new_n495), .C2(KEYINPUT29), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n484), .B1(new_n483), .B2(new_n479), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n490), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n489), .B1(new_n498), .B2(new_n442), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n480), .B1(new_n479), .B2(new_n483), .ZN(new_n500));
  OR2_X1    g299(.A1(new_n500), .A2(new_n487), .ZN(new_n501));
  XNOR2_X1  g300(.A(G8gat), .B(G36gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(G64gat), .B(G92gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n502), .B(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n488), .A2(new_n499), .A3(new_n501), .A4(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT30), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n488), .A2(new_n499), .A3(new_n501), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT76), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT76), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n488), .A2(new_n499), .A3(new_n511), .A4(new_n501), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n505), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n508), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT82), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n446), .A2(new_n449), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n451), .A2(new_n452), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n518), .B1(new_n401), .B2(new_n396), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT4), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n453), .A2(new_n389), .A3(new_n395), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT4), .ZN(new_n522));
  NAND2_X1  g321(.A1(G225gat), .A2(G233gat), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n521), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT79), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n526), .B1(new_n453), .B2(new_n454), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n518), .A2(KEYINPUT79), .A3(KEYINPUT3), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n527), .A2(new_n528), .A3(new_n400), .A4(new_n455), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n520), .A2(new_n525), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT5), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n400), .A2(new_n518), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(new_n521), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n531), .B1(new_n533), .B2(new_n524), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  OR2_X1    g334(.A1(new_n519), .A2(KEYINPUT4), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n524), .A2(KEYINPUT5), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n521), .A2(new_n522), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n536), .A2(new_n529), .A3(new_n537), .A4(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(G57gat), .B(G85gat), .Z(new_n541));
  XNOR2_X1  g340(.A(G1gat), .B(G29gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  XOR2_X1   g342(.A(KEYINPUT80), .B(KEYINPUT0), .Z(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(KEYINPUT81), .ZN(new_n545));
  XOR2_X1   g344(.A(new_n543), .B(new_n545), .Z(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n540), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT6), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n515), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n546), .B1(new_n535), .B2(new_n539), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n551), .A2(KEYINPUT82), .A3(KEYINPUT6), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n535), .A2(new_n539), .A3(new_n546), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n548), .A2(new_n549), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n550), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n477), .A2(new_n514), .A3(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(KEYINPUT35), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT86), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT40), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT39), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n533), .A2(new_n524), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n529), .B(new_n538), .C1(new_n519), .C2(KEYINPUT4), .ZN(new_n562));
  AOI211_X1 g361(.A(new_n560), .B(new_n561), .C1(new_n562), .C2(new_n524), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(new_n560), .A3(new_n524), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(new_n546), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n558), .B(new_n559), .C1(new_n563), .C2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(new_n548), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n561), .B1(new_n562), .B2(new_n524), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(KEYINPUT39), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n569), .A2(new_n546), .A3(new_n564), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n559), .B1(new_n570), .B2(new_n558), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n572), .B1(new_n508), .B2(new_n513), .ZN(new_n573));
  INV_X1    g372(.A(new_n476), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT38), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n510), .A2(new_n512), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT37), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT37), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n488), .A2(new_n499), .A3(new_n578), .A4(new_n501), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n579), .A2(new_n504), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n575), .B1(new_n577), .B2(new_n580), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n551), .A2(KEYINPUT82), .A3(KEYINPUT6), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT82), .B1(new_n551), .B2(KEYINPUT6), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n500), .A2(new_n442), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n585), .B1(new_n486), .B2(new_n442), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT38), .B1(new_n586), .B2(KEYINPUT37), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n587), .A2(new_n579), .A3(new_n504), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n584), .A2(new_n554), .A3(new_n506), .A4(new_n588), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n573), .B(new_n574), .C1(new_n581), .C2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT36), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n591), .B1(new_n432), .B2(new_n434), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n422), .A2(new_n431), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n433), .A2(new_n416), .A3(new_n430), .A4(new_n429), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n593), .A2(new_n594), .A3(KEYINPUT36), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n576), .A2(new_n504), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n506), .B(KEYINPUT30), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n597), .A2(new_n555), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n596), .B1(new_n476), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n590), .A2(new_n600), .ZN(new_n601));
  AOI211_X1 g400(.A(new_n293), .B(new_n335), .C1(new_n557), .C2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n555), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(G1gat), .ZN(G1324gat));
  INV_X1    g404(.A(new_n514), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  OR2_X1    g406(.A1(new_n607), .A2(KEYINPUT99), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(KEYINPUT99), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT42), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n608), .B(new_n609), .C1(new_n610), .C2(G8gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT16), .B(G8gat), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n612), .B1(new_n607), .B2(KEYINPUT42), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT100), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n613), .B1(new_n614), .B2(KEYINPUT42), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n612), .A2(KEYINPUT100), .A3(new_n610), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n611), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT101), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n611), .A2(KEYINPUT101), .A3(new_n615), .A4(new_n616), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(G1325gat));
  INV_X1    g420(.A(new_n435), .ZN(new_n622));
  AOI21_X1  g421(.A(G15gat), .B1(new_n602), .B2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT102), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n602), .A2(G15gat), .A3(new_n596), .ZN(new_n625));
  AND2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(G1326gat));
  NAND2_X1  g425(.A1(new_n602), .A2(new_n476), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT43), .B(G22gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(G1327gat));
  AOI21_X1  g428(.A(new_n334), .B1(new_n557), .B2(new_n601), .ZN(new_n630));
  INV_X1    g429(.A(G29gat), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n310), .A2(new_n293), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n630), .A2(new_n631), .A3(new_n603), .A4(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n630), .A2(KEYINPUT44), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT104), .ZN(new_n640));
  AND3_X1   g439(.A1(new_n590), .A2(new_n600), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n640), .B1(new_n590), .B2(new_n600), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n334), .B1(new_n643), .B2(new_n557), .ZN(new_n644));
  OAI211_X1 g443(.A(new_n632), .B(new_n639), .C1(new_n644), .C2(KEYINPUT44), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(KEYINPUT105), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n601), .A2(KEYINPUT104), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n590), .A2(new_n600), .A3(new_n640), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n647), .A2(new_n557), .A3(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n334), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT44), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT105), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n653), .A2(new_n654), .A3(new_n632), .A4(new_n639), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n555), .B1(new_n646), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n638), .B1(new_n656), .B2(new_n631), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT106), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n638), .B(KEYINPUT106), .C1(new_n656), .C2(new_n631), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(G1328gat));
  NAND2_X1  g460(.A1(new_n630), .A2(new_n632), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n662), .A2(G36gat), .A3(new_n514), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT107), .B(KEYINPUT46), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n514), .B1(new_n646), .B2(new_n655), .ZN(new_n666));
  INV_X1    g465(.A(G36gat), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(G1329gat));
  INV_X1    g467(.A(new_n596), .ZN(new_n669));
  OAI21_X1  g468(.A(G43gat), .B1(new_n645), .B2(new_n669), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n662), .A2(G43gat), .A3(new_n435), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n670), .A2(KEYINPUT47), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n646), .A2(new_n655), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(new_n596), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n671), .B1(new_n675), .B2(G43gat), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n673), .B1(new_n676), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g476(.A(G50gat), .B1(new_n645), .B2(new_n574), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n662), .A2(G50gat), .A3(new_n574), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n678), .A2(KEYINPUT48), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n674), .A2(new_n476), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n679), .B1(new_n682), .B2(G50gat), .ZN(new_n683));
  XOR2_X1   g482(.A(KEYINPUT108), .B(KEYINPUT48), .Z(new_n684));
  OAI21_X1  g483(.A(new_n681), .B1(new_n683), .B2(new_n684), .ZN(G1331gat));
  NOR2_X1   g484(.A1(new_n335), .A2(new_n292), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n649), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n246), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n555), .B(KEYINPUT109), .Z(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(G57gat), .ZN(G1332gat));
  XOR2_X1   g491(.A(new_n514), .B(KEYINPUT110), .Z(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n688), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n696));
  AND2_X1   g495(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n695), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n698), .B1(new_n695), .B2(new_n696), .ZN(G1333gat));
  INV_X1    g498(.A(G71gat), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n700), .B1(new_n688), .B2(new_n435), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT111), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n688), .A2(new_n700), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n702), .B1(new_n703), .B2(new_n596), .ZN(new_n704));
  NOR4_X1   g503(.A1(new_n688), .A2(KEYINPUT111), .A3(new_n700), .A4(new_n669), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n701), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(KEYINPUT50), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT50), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n708), .B(new_n701), .C1(new_n704), .C2(new_n705), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n709), .ZN(G1334gat));
  NAND2_X1  g509(.A1(new_n689), .A2(new_n476), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g511(.A1(new_n310), .A2(new_n292), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n653), .A2(new_n246), .A3(new_n639), .A4(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(G85gat), .B1(new_n714), .B2(new_n555), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n644), .A2(KEYINPUT51), .A3(new_n713), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n649), .A2(new_n650), .A3(new_n713), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT51), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n603), .A2(new_n217), .A3(new_n246), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT112), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n715), .B1(new_n721), .B2(new_n723), .ZN(G1336gat));
  OAI21_X1  g523(.A(G92gat), .B1(new_n714), .B2(new_n694), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT52), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n693), .A2(new_n218), .A3(new_n246), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n725), .B(new_n726), .C1(new_n721), .C2(new_n727), .ZN(new_n728));
  OR2_X1    g527(.A1(new_n714), .A2(new_n514), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n727), .B(KEYINPUT113), .ZN(new_n730));
  AOI22_X1  g529(.A1(new_n729), .A2(G92gat), .B1(new_n720), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n728), .B1(new_n731), .B2(new_n726), .ZN(G1337gat));
  XNOR2_X1  g531(.A(KEYINPUT114), .B(G99gat), .ZN(new_n733));
  OR4_X1    g532(.A1(new_n247), .A2(new_n721), .A3(new_n435), .A4(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n714), .B2(new_n669), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(G1338gat));
  OAI21_X1  g535(.A(G106gat), .B1(new_n714), .B2(new_n574), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n574), .A2(G106gat), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n720), .A2(new_n246), .A3(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n737), .A2(new_n739), .A3(KEYINPUT115), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g540(.A1(new_n335), .A2(new_n246), .A3(new_n292), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT116), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n232), .A2(new_n233), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT54), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n240), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(KEYINPUT54), .B1(new_n232), .B2(new_n233), .ZN(new_n747));
  OAI211_X1 g546(.A(new_n746), .B(KEYINPUT55), .C1(new_n744), .C2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT55), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n744), .A2(new_n747), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n239), .B1(new_n234), .B2(KEYINPUT54), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n243), .A2(new_n748), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n273), .B1(new_n271), .B2(new_n272), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n279), .A2(new_n280), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n287), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n291), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n650), .A2(new_n743), .A3(new_n753), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n246), .A2(new_n757), .ZN(new_n759));
  INV_X1    g558(.A(new_n292), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n243), .A2(new_n748), .A3(new_n752), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n334), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n753), .A2(new_n332), .A3(new_n333), .A4(new_n757), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(KEYINPUT116), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n758), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n310), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n742), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n477), .ZN(new_n769));
  INV_X1    g568(.A(new_n690), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n771), .A2(new_n694), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n772), .A2(new_n378), .A3(new_n292), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n768), .A2(new_n769), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n774), .A2(new_n603), .A3(new_n694), .ZN(new_n775));
  OAI21_X1  g574(.A(G113gat), .B1(new_n775), .B2(new_n760), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n773), .A2(new_n776), .ZN(G1340gat));
  OAI211_X1 g576(.A(new_n772), .B(new_n246), .C1(new_n383), .C2(new_n384), .ZN(new_n778));
  OAI21_X1  g577(.A(G120gat), .B1(new_n775), .B2(new_n247), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(G1341gat));
  INV_X1    g579(.A(G127gat), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n775), .A2(new_n781), .A3(new_n767), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n772), .A2(new_n310), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n782), .B1(new_n783), .B2(new_n781), .ZN(G1342gat));
  NOR2_X1   g583(.A1(new_n606), .A2(new_n334), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n771), .A2(new_n392), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n786), .A2(KEYINPUT56), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT117), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(KEYINPUT56), .ZN(new_n789));
  OAI21_X1  g588(.A(G134gat), .B1(new_n775), .B2(new_n334), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n788), .A2(new_n789), .A3(new_n790), .ZN(G1343gat));
  XNOR2_X1  g590(.A(new_n764), .B(new_n743), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n761), .A2(KEYINPUT118), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n243), .A2(new_n748), .A3(new_n794), .A4(new_n752), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n793), .A2(new_n292), .A3(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n650), .B1(new_n796), .B2(new_n759), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n310), .B1(new_n792), .B2(new_n798), .ZN(new_n799));
  OAI211_X1 g598(.A(KEYINPUT57), .B(new_n476), .C1(new_n799), .C2(new_n742), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT119), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n766), .A2(new_n767), .ZN(new_n803));
  INV_X1    g602(.A(new_n742), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n476), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n758), .A2(new_n765), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n767), .B1(new_n809), .B2(new_n797), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n807), .B1(new_n810), .B2(new_n804), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n811), .A2(KEYINPUT119), .A3(new_n476), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n802), .A2(new_n808), .A3(new_n812), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n693), .A2(new_n555), .A3(new_n596), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(G141gat), .B1(new_n815), .B2(new_n760), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT121), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n817), .B1(new_n768), .B2(new_n770), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n805), .A2(KEYINPUT121), .A3(new_n690), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n596), .A2(new_n574), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n818), .A2(new_n819), .A3(new_n694), .A4(new_n820), .ZN(new_n821));
  OR3_X1    g620(.A1(new_n821), .A2(G141gat), .A3(new_n760), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n816), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT58), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT120), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n824), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n816), .B(new_n822), .C1(new_n825), .C2(new_n824), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(G1344gat));
  INV_X1    g628(.A(KEYINPUT59), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n830), .B(G148gat), .C1(new_n815), .C2(new_n247), .ZN(new_n831));
  INV_X1    g630(.A(G148gat), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n806), .A2(KEYINPUT57), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n310), .B1(new_n798), .B2(new_n764), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n807), .B(new_n476), .C1(new_n834), .C2(new_n742), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n833), .A2(new_n246), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n832), .B1(new_n836), .B2(new_n814), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n831), .B1(new_n830), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n246), .A2(new_n832), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n838), .B1(new_n821), .B2(new_n839), .ZN(G1345gat));
  NAND2_X1  g639(.A1(new_n310), .A2(G155gat), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(KEYINPUT122), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n821), .A2(new_n767), .ZN(new_n843));
  OAI22_X1  g642(.A1(new_n815), .A2(new_n842), .B1(new_n843), .B2(G155gat), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT123), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n844), .B(new_n845), .ZN(G1346gat));
  OAI21_X1  g645(.A(new_n444), .B1(new_n815), .B2(new_n334), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n334), .A2(new_n606), .A3(new_n444), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n818), .A2(new_n819), .A3(new_n820), .A4(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n849), .ZN(G1347gat));
  NOR2_X1   g649(.A1(new_n694), .A2(new_n603), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n774), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n852), .A2(new_n341), .A3(new_n292), .ZN(new_n853));
  NOR4_X1   g652(.A1(new_n768), .A2(new_n514), .A3(new_n769), .A4(new_n690), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n854), .A2(new_n292), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n853), .B1(new_n855), .B2(new_n341), .ZN(G1348gat));
  AOI21_X1  g655(.A(G176gat), .B1(new_n852), .B2(new_n246), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n247), .A2(new_n342), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n857), .B1(new_n854), .B2(new_n858), .ZN(G1349gat));
  INV_X1    g658(.A(new_n369), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n852), .A2(new_n860), .A3(new_n310), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n854), .A2(new_n310), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n861), .B1(new_n862), .B2(new_n356), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g663(.A(new_n357), .B1(new_n854), .B2(new_n650), .ZN(new_n865));
  XOR2_X1   g664(.A(new_n865), .B(KEYINPUT61), .Z(new_n866));
  NAND3_X1  g665(.A1(new_n852), .A2(new_n357), .A3(new_n650), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(G1351gat));
  XNOR2_X1  g667(.A(KEYINPUT124), .B(G197gat), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n833), .A2(new_n835), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n690), .A2(new_n514), .A3(new_n596), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n869), .B1(new_n872), .B2(new_n760), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n805), .A2(new_n851), .A3(new_n820), .ZN(new_n874));
  INV_X1    g673(.A(new_n869), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n874), .A2(new_n292), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n873), .A2(new_n876), .ZN(G1352gat));
  INV_X1    g676(.A(G204gat), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n874), .A2(new_n878), .A3(new_n246), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT62), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n878), .B1(new_n836), .B2(new_n871), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n880), .A2(new_n881), .ZN(G1353gat));
  NAND3_X1  g681(.A1(new_n874), .A2(new_n437), .A3(new_n310), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n870), .A2(new_n310), .A3(new_n871), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n884), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n885));
  AOI21_X1  g684(.A(KEYINPUT63), .B1(new_n884), .B2(G211gat), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n883), .B1(new_n885), .B2(new_n886), .ZN(G1354gat));
  AOI21_X1  g686(.A(G218gat), .B1(new_n874), .B2(new_n650), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(KEYINPUT125), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT126), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n872), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(new_n334), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n438), .B1(new_n872), .B2(new_n890), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n889), .B1(new_n892), .B2(new_n893), .ZN(G1355gat));
endmodule


