//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 1 0 1 0 0 0 1 1 0 0 0 1 0 1 1 1 1 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 1 0 0 1 0 0 0 1 1 0 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:10 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT9), .B(G234), .Z(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n187), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G104), .ZN(new_n191));
  OAI21_X1  g005(.A(KEYINPUT3), .B1(new_n191), .B2(G107), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT78), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  OR3_X1    g008(.A1(new_n191), .A2(KEYINPUT3), .A3(G107), .ZN(new_n195));
  INV_X1    g009(.A(G107), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G104), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  OAI211_X1 g012(.A(KEYINPUT78), .B(KEYINPUT3), .C1(new_n191), .C2(G107), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n194), .A2(new_n195), .A3(new_n198), .A4(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G101), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT79), .ZN(new_n202));
  NOR3_X1   g016(.A1(new_n191), .A2(KEYINPUT3), .A3(G107), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(new_n197), .ZN(new_n204));
  INV_X1    g018(.A(G101), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n204), .A2(new_n205), .A3(new_n194), .A4(new_n199), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT4), .A4(new_n206), .ZN(new_n207));
  AND3_X1   g021(.A1(new_n201), .A2(KEYINPUT4), .A3(new_n206), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT4), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n200), .A2(new_n209), .A3(G101), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT79), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n207), .B1(new_n208), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G146), .ZN(new_n214));
  INV_X1    g028(.A(G146), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G143), .ZN(new_n216));
  AND3_X1   g030(.A1(new_n214), .A2(new_n216), .A3(G128), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT64), .B1(new_n213), .B2(G146), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT64), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(new_n215), .A3(G143), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n218), .A2(new_n220), .A3(new_n214), .ZN(new_n221));
  XOR2_X1   g035(.A(KEYINPUT0), .B(G128), .Z(new_n222));
  AOI22_X1  g036(.A1(KEYINPUT0), .A2(new_n217), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n212), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT11), .ZN(new_n225));
  INV_X1    g039(.A(G134), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n225), .B1(new_n226), .B2(G137), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(G137), .ZN(new_n228));
  INV_X1    g042(.A(G137), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(KEYINPUT11), .A3(G134), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n227), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G131), .ZN(new_n232));
  INV_X1    g046(.A(G131), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n227), .A2(new_n230), .A3(new_n233), .A4(new_n228), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT1), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n214), .A2(new_n216), .A3(new_n237), .A4(G128), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n214), .A2(new_n216), .ZN(new_n239));
  INV_X1    g053(.A(G128), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n240), .B1(new_n216), .B2(KEYINPUT1), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n238), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n191), .A2(G107), .ZN(new_n243));
  OAI21_X1  g057(.A(G101), .B1(new_n243), .B2(new_n197), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n206), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT10), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT80), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n245), .A2(KEYINPUT80), .A3(new_n246), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT81), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n206), .A2(new_n252), .A3(new_n244), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n252), .B1(new_n206), .B2(new_n244), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT1), .B1(new_n213), .B2(G146), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G128), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n221), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n238), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n255), .A2(KEYINPUT10), .A3(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n224), .A2(new_n236), .A3(new_n251), .A4(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n206), .A2(new_n244), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n262), .A2(new_n258), .A3(new_n238), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n236), .B1(new_n263), .B2(new_n245), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n264), .B(KEYINPUT12), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n261), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT77), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n224), .A2(new_n251), .A3(new_n260), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n235), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n261), .ZN(new_n270));
  XNOR2_X1  g084(.A(G110), .B(G140), .ZN(new_n271));
  INV_X1    g085(.A(G953), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G227), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n271), .B(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n267), .A2(new_n270), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n274), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n261), .A2(new_n265), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n276), .B1(new_n277), .B2(KEYINPUT77), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(G469), .B1(new_n279), .B2(G902), .ZN(new_n280));
  INV_X1    g094(.A(G469), .ZN(new_n281));
  XOR2_X1   g095(.A(KEYINPUT72), .B(G902), .Z(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n264), .A2(KEYINPUT12), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT82), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT12), .ZN(new_n287));
  AOI211_X1 g101(.A(new_n287), .B(new_n236), .C1(new_n263), .C2(new_n245), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n285), .A2(new_n286), .A3(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(KEYINPUT82), .B1(new_n284), .B2(new_n288), .ZN(new_n291));
  AND4_X1   g105(.A1(new_n261), .A2(new_n290), .A3(new_n291), .A4(new_n274), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n274), .B1(new_n269), .B2(new_n261), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n281), .B(new_n283), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n190), .B1(new_n280), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(G214), .B1(G237), .B2(G902), .ZN(new_n296));
  OAI21_X1  g110(.A(G210), .B1(G237), .B2(G902), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT90), .ZN(new_n299));
  INV_X1    g113(.A(G125), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT73), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT73), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G125), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n223), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT73), .B(G125), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n259), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G224), .ZN(new_n309));
  OAI21_X1  g123(.A(KEYINPUT7), .B1(new_n309), .B2(G953), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n310), .B1(new_n305), .B2(new_n307), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT88), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n262), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT5), .ZN(new_n317));
  INV_X1    g131(.A(G119), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n318), .A3(G116), .ZN(new_n319));
  XNOR2_X1  g133(.A(G116), .B(G119), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  OAI211_X1 g135(.A(G113), .B(new_n319), .C1(new_n321), .C2(new_n317), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT2), .B(G113), .ZN(new_n323));
  OR2_X1    g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n206), .A2(KEYINPUT88), .A3(new_n244), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n316), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(G110), .B(G122), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n328), .B(KEYINPUT84), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT8), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n329), .B(new_n330), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n262), .A2(new_n315), .A3(new_n324), .A4(new_n322), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n327), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT89), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n327), .A2(KEYINPUT89), .A3(new_n331), .A4(new_n332), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n314), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT85), .ZN(new_n338));
  NOR3_X1   g152(.A1(new_n253), .A2(new_n254), .A3(new_n325), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n321), .A2(new_n323), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n324), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n339), .B1(new_n212), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n329), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n338), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n341), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n201), .A2(KEYINPUT4), .A3(new_n206), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(KEYINPUT79), .A3(new_n210), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n345), .B1(new_n347), .B2(new_n207), .ZN(new_n348));
  NOR4_X1   g162(.A1(new_n348), .A2(KEYINPUT85), .A3(new_n329), .A4(new_n339), .ZN(new_n349));
  OAI22_X1  g163(.A1(new_n299), .A2(new_n337), .B1(new_n344), .B2(new_n349), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n337), .A2(new_n299), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n189), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n309), .A2(G953), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n353), .B(KEYINPUT87), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n308), .B(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n212), .A2(new_n341), .ZN(new_n356));
  INV_X1    g170(.A(new_n339), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT83), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT83), .ZN(new_n359));
  NOR3_X1   g173(.A1(new_n348), .A2(new_n359), .A3(new_n339), .ZN(new_n360));
  OAI211_X1 g174(.A(KEYINPUT86), .B(new_n329), .C1(new_n358), .C2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT6), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n344), .A2(new_n349), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n329), .B1(new_n358), .B2(new_n360), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n342), .A2(KEYINPUT83), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n359), .B1(new_n348), .B2(new_n339), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n369), .A2(KEYINPUT86), .A3(KEYINPUT6), .A4(new_n329), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n363), .A2(new_n366), .A3(new_n370), .ZN(new_n371));
  AOI211_X1 g185(.A(new_n298), .B(new_n352), .C1(new_n355), .C2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n355), .ZN(new_n373));
  INV_X1    g187(.A(new_n352), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n297), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n295), .B(new_n296), .C1(new_n372), .C2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT16), .ZN(new_n378));
  INV_X1    g192(.A(G140), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n301), .A2(new_n303), .A3(new_n378), .A4(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT75), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n306), .A2(KEYINPUT75), .A3(new_n378), .A4(new_n379), .ZN(new_n383));
  AND2_X1   g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(KEYINPUT74), .B1(new_n379), .B2(G125), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n385), .B1(new_n306), .B2(new_n379), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n304), .A2(KEYINPUT74), .A3(G140), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n378), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n215), .B1(new_n384), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT74), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n390), .B1(new_n300), .B2(G140), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n391), .B1(new_n304), .B2(G140), .ZN(new_n392));
  AOI211_X1 g206(.A(new_n390), .B(new_n379), .C1(new_n301), .C2(new_n303), .ZN(new_n393));
  OAI21_X1  g207(.A(KEYINPUT16), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n382), .A2(new_n383), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(G146), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n389), .A2(new_n396), .A3(KEYINPUT76), .ZN(new_n397));
  XOR2_X1   g211(.A(KEYINPUT24), .B(G110), .Z(new_n398));
  XNOR2_X1  g212(.A(G119), .B(G128), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NOR3_X1   g214(.A1(new_n318), .A2(KEYINPUT23), .A3(G128), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n401), .B1(new_n399), .B2(KEYINPUT23), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G110), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT76), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n404), .B(new_n215), .C1(new_n384), .C2(new_n388), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n397), .A2(new_n400), .A3(new_n403), .A4(new_n405), .ZN(new_n406));
  OAI22_X1  g220(.A1(new_n402), .A2(G110), .B1(new_n399), .B2(new_n398), .ZN(new_n407));
  XOR2_X1   g221(.A(G125), .B(G140), .Z(new_n408));
  OR2_X1    g222(.A1(new_n408), .A2(G146), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n396), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n272), .A2(G221), .A3(G234), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n412), .B(KEYINPUT22), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n413), .B(G137), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n411), .B(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n283), .ZN(new_n416));
  OR2_X1    g230(.A1(new_n416), .A2(KEYINPUT25), .ZN(new_n417));
  INV_X1    g231(.A(G217), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n418), .B1(new_n283), .B2(G234), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n416), .A2(KEYINPUT25), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n417), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n419), .A2(G902), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n415), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT67), .ZN(new_n426));
  XNOR2_X1  g240(.A(G134), .B(G137), .ZN(new_n427));
  OAI21_X1  g241(.A(KEYINPUT65), .B1(new_n427), .B2(new_n233), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT65), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n229), .A2(G134), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n226), .A2(G137), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n429), .B(G131), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n259), .A2(new_n234), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n223), .A2(new_n235), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT66), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT30), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(KEYINPUT66), .A2(KEYINPUT30), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n436), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n434), .A2(new_n435), .A3(new_n437), .A4(new_n438), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n426), .B1(new_n445), .B2(new_n341), .ZN(new_n446));
  AOI211_X1 g260(.A(KEYINPUT67), .B(new_n345), .C1(new_n443), .C2(new_n444), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n345), .A2(new_n434), .A3(new_n435), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n451), .B(G101), .ZN(new_n452));
  INV_X1    g266(.A(G237), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n453), .A2(new_n272), .A3(G210), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n452), .B(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n450), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT29), .ZN(new_n458));
  INV_X1    g272(.A(new_n449), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n345), .B1(new_n434), .B2(new_n435), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT28), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  OR2_X1    g275(.A1(new_n461), .A2(KEYINPUT69), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT28), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n449), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n461), .A2(KEYINPUT69), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n462), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n457), .B(new_n458), .C1(new_n456), .C2(new_n466), .ZN(new_n467));
  OR2_X1    g281(.A1(new_n459), .A2(new_n460), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n468), .A2(KEYINPUT70), .A3(KEYINPUT28), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n464), .B(KEYINPUT71), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT70), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n461), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n469), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n455), .A2(KEYINPUT29), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n467), .B(new_n283), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(G472), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT31), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT68), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n448), .A2(new_n478), .A3(new_n455), .A4(new_n449), .ZN(new_n479));
  AOI211_X1 g293(.A(new_n439), .B(new_n441), .C1(new_n434), .C2(new_n435), .ZN(new_n480));
  AND4_X1   g294(.A1(new_n437), .A2(new_n434), .A3(new_n438), .A4(new_n435), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n341), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT67), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n445), .A2(new_n426), .A3(new_n341), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n483), .A2(new_n455), .A3(new_n449), .A4(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(KEYINPUT68), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n477), .B1(new_n479), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n466), .A2(new_n456), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n485), .A2(KEYINPUT31), .ZN(new_n490));
  NOR3_X1   g304(.A1(new_n487), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(G472), .A2(G902), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NOR3_X1   g307(.A1(new_n491), .A2(KEYINPUT32), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT32), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n485), .A2(KEYINPUT68), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n485), .A2(KEYINPUT68), .ZN(new_n497));
  OAI21_X1  g311(.A(KEYINPUT31), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n490), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n488), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n495), .B1(new_n500), .B2(new_n492), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n476), .B1(new_n494), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(G475), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n453), .A2(new_n272), .A3(G214), .ZN(new_n504));
  NAND2_X1  g318(.A1(KEYINPUT91), .A2(G143), .ZN(new_n505));
  OR2_X1    g319(.A1(KEYINPUT91), .A2(G143), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(KEYINPUT91), .A2(G143), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n508), .A2(G214), .A3(new_n453), .A4(new_n272), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(KEYINPUT18), .A2(G131), .ZN(new_n511));
  XOR2_X1   g325(.A(new_n510), .B(new_n511), .Z(new_n512));
  NAND2_X1  g326(.A1(new_n386), .A2(new_n387), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n409), .B1(new_n513), .B2(new_n215), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n397), .A2(KEYINPUT95), .A3(new_n405), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n510), .A2(new_n233), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT17), .ZN(new_n518));
  AOI21_X1  g332(.A(G131), .B1(new_n507), .B2(new_n509), .ZN(new_n519));
  OR3_X1    g333(.A1(new_n517), .A2(KEYINPUT17), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n516), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(KEYINPUT95), .B1(new_n397), .B2(new_n405), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n515), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  XOR2_X1   g337(.A(G113), .B(G122), .Z(new_n524));
  XNOR2_X1  g338(.A(new_n524), .B(KEYINPUT93), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n525), .B(new_n191), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT97), .ZN(new_n527));
  OR2_X1    g341(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(G902), .B1(new_n523), .B2(new_n527), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n503), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n526), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n532), .B(new_n515), .C1(new_n521), .C2(new_n522), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n517), .A2(new_n519), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n384), .A2(new_n388), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n534), .B1(new_n535), .B2(G146), .ZN(new_n536));
  OAI21_X1  g350(.A(KEYINPUT92), .B1(new_n408), .B2(KEYINPUT19), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT19), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n537), .B1(new_n513), .B2(new_n538), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n386), .A2(new_n387), .A3(KEYINPUT92), .A4(KEYINPUT19), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n539), .A2(new_n215), .A3(new_n540), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n536), .A2(new_n541), .B1(new_n514), .B2(new_n512), .ZN(new_n542));
  OAI21_X1  g356(.A(KEYINPUT94), .B1(new_n542), .B2(new_n532), .ZN(new_n543));
  INV_X1    g357(.A(new_n541), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n396), .B1(new_n517), .B2(new_n519), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n515), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT94), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(new_n547), .A3(new_n526), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n543), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n533), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n550), .A2(new_n503), .A3(new_n189), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT96), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n552), .B1(new_n533), .B2(new_n549), .ZN(new_n553));
  NOR3_X1   g367(.A1(new_n551), .A2(KEYINPUT20), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n550), .A2(KEYINPUT96), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT20), .ZN(new_n556));
  AOI21_X1  g370(.A(G475), .B1(new_n533), .B2(new_n549), .ZN(new_n557));
  AOI22_X1  g371(.A1(new_n555), .A2(new_n556), .B1(new_n557), .B2(new_n189), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n531), .B1(new_n554), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(G952), .ZN(new_n560));
  AOI211_X1 g374(.A(G953), .B(new_n560), .C1(G234), .C2(G237), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  AOI211_X1 g376(.A(new_n272), .B(new_n283), .C1(G234), .C2(G237), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  XOR2_X1   g378(.A(KEYINPUT21), .B(G898), .Z(new_n565));
  OAI21_X1  g379(.A(new_n562), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(G128), .B(G143), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(new_n226), .ZN(new_n569));
  XNOR2_X1  g383(.A(G116), .B(G122), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT14), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(G116), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(KEYINPUT14), .A3(G122), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n572), .A2(G107), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n570), .A2(new_n196), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n569), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT98), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n568), .A2(KEYINPUT13), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n213), .A2(G128), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n580), .B(G134), .C1(KEYINPUT13), .C2(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n570), .B(new_n196), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n568), .A2(new_n226), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n579), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n188), .A2(G217), .A3(new_n272), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(KEYINPUT99), .ZN(new_n588));
  OR2_X1    g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n586), .A2(new_n588), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n282), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT100), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n591), .A2(new_n592), .ZN(new_n594));
  INV_X1    g408(.A(G478), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(KEYINPUT15), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n593), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n597), .B1(new_n596), .B2(new_n593), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n559), .A2(new_n567), .A3(new_n598), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n377), .A2(new_n425), .A3(new_n502), .A4(new_n599), .ZN(new_n600));
  XOR2_X1   g414(.A(KEYINPUT101), .B(G101), .Z(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(G3));
  OAI21_X1  g416(.A(G472), .B1(new_n491), .B2(new_n282), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n500), .A2(new_n492), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n280), .A2(new_n294), .ZN(new_n606));
  INV_X1    g420(.A(new_n190), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n605), .A2(new_n424), .A3(new_n608), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n296), .B(new_n566), .C1(new_n372), .C2(new_n375), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n551), .B1(KEYINPUT20), .B2(new_n553), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n555), .A2(new_n556), .A3(new_n189), .A4(new_n557), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n530), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n589), .A2(new_n590), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT33), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n282), .A2(new_n595), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n589), .A2(KEYINPUT103), .ZN(new_n618));
  OR3_X1    g432(.A1(new_n586), .A2(KEYINPUT103), .A3(new_n588), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n618), .A2(KEYINPUT33), .A3(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n590), .B(KEYINPUT102), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n616), .B(new_n617), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  OR2_X1    g436(.A1(new_n591), .A2(G478), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n613), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n610), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n609), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(KEYINPUT104), .B(KEYINPUT34), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(G104), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n629), .B(new_n631), .ZN(G6));
  XNOR2_X1  g446(.A(new_n551), .B(KEYINPUT20), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n633), .A2(new_n531), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n598), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n635), .A2(new_n610), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n609), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT35), .B(G107), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G9));
  INV_X1    g453(.A(new_n605), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n411), .B(KEYINPUT105), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT36), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n414), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n641), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n422), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n421), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n377), .A2(new_n640), .A3(new_n599), .A4(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(new_n647), .B(KEYINPUT37), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G110), .ZN(G12));
  OAI21_X1  g463(.A(KEYINPUT32), .B1(new_n491), .B2(new_n493), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n500), .A2(new_n495), .A3(new_n492), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n650), .A2(new_n651), .B1(G472), .B2(new_n475), .ZN(new_n652));
  INV_X1    g466(.A(new_n646), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n652), .A2(new_n376), .A3(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(G900), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n561), .B1(new_n563), .B2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n635), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G128), .ZN(G30));
  NAND2_X1  g473(.A1(new_n373), .A2(new_n374), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n298), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n373), .A2(new_n374), .A3(new_n297), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(KEYINPUT106), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n372), .A2(new_n375), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT106), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n664), .A2(new_n667), .A3(KEYINPUT38), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT38), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n372), .A2(new_n375), .A3(KEYINPUT106), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n666), .B1(new_n661), .B2(new_n662), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n669), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n559), .A2(new_n296), .A3(new_n598), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n650), .A2(new_n651), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n479), .A2(new_n486), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n468), .A2(new_n456), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT107), .ZN(new_n679));
  AOI21_X1  g493(.A(G902), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(G472), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n646), .B1(new_n676), .B2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n656), .B(KEYINPUT39), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n608), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT40), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n675), .A2(new_n683), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G143), .ZN(G45));
  INV_X1    g502(.A(new_n656), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n559), .A2(new_n624), .A3(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n654), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G146), .ZN(G48));
  INV_X1    g507(.A(KEYINPUT108), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n283), .B1(new_n292), .B2(new_n293), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(G469), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n696), .A2(new_n607), .A3(new_n294), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n502), .A2(new_n425), .A3(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n296), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n699), .B1(new_n661), .B2(new_n662), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n700), .A2(new_n566), .A3(new_n626), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n694), .B1(new_n698), .B2(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n652), .A2(new_n424), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n703), .A2(KEYINPUT108), .A3(new_n628), .A4(new_n697), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT41), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G113), .ZN(G15));
  NAND3_X1  g521(.A1(new_n703), .A2(new_n636), .A3(new_n697), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G116), .ZN(G18));
  OAI211_X1 g523(.A(new_n697), .B(new_n296), .C1(new_n372), .C2(new_n375), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT109), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n663), .A2(KEYINPUT109), .A3(new_n296), .A4(new_n697), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n653), .B1(new_n676), .B2(new_n476), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n714), .A2(new_n599), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  NAND2_X1  g531(.A1(new_n473), .A2(new_n456), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n498), .A2(new_n499), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n603), .B1(new_n493), .B2(new_n719), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n720), .A2(new_n424), .A3(new_n567), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n696), .A2(new_n294), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n607), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n674), .A2(new_n665), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G122), .ZN(G24));
  NAND2_X1  g540(.A1(new_n690), .A2(KEYINPUT110), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT110), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n559), .A2(new_n728), .A3(new_n624), .A4(new_n689), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n720), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n714), .A2(new_n730), .A3(new_n646), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G125), .ZN(G27));
  INV_X1    g546(.A(KEYINPUT42), .ZN(new_n733));
  AND4_X1   g547(.A1(new_n296), .A2(new_n295), .A3(new_n661), .A4(new_n662), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(new_n502), .A3(new_n425), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n728), .B1(new_n626), .B2(new_n689), .ZN(new_n736));
  NOR4_X1   g550(.A1(new_n613), .A2(new_n625), .A3(KEYINPUT110), .A4(new_n656), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n733), .B1(new_n735), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n727), .A2(new_n729), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n703), .A2(new_n740), .A3(KEYINPUT42), .A4(new_n734), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G131), .ZN(G33));
  NAND3_X1  g557(.A1(new_n703), .A2(new_n657), .A3(new_n734), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G134), .ZN(G36));
  NAND2_X1  g559(.A1(new_n279), .A2(KEYINPUT45), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT45), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n275), .A2(new_n278), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n746), .A2(G469), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(G469), .A2(G902), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(KEYINPUT46), .A3(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT111), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n749), .A2(new_n750), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT46), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n749), .A2(KEYINPUT111), .A3(KEYINPUT46), .A4(new_n750), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n753), .A2(new_n756), .A3(new_n294), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n607), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n759), .A2(new_n684), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n665), .A2(new_n296), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n613), .A2(new_n624), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT43), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n613), .A2(KEYINPUT43), .A3(new_n624), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n605), .A3(new_n646), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT44), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n761), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n766), .A2(KEYINPUT44), .A3(new_n605), .A4(new_n646), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n760), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(KEYINPUT112), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(new_n229), .ZN(G39));
  INV_X1    g587(.A(KEYINPUT47), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n759), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n758), .A2(KEYINPUT47), .A3(new_n607), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n502), .A2(new_n761), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n777), .A2(new_n424), .A3(new_n691), .A4(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G140), .ZN(G42));
  INV_X1    g594(.A(KEYINPUT118), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n674), .A2(new_n665), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n682), .B1(new_n494), .B2(new_n501), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n608), .A2(new_n656), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n783), .A2(new_n653), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT114), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n377), .B(new_n715), .C1(new_n657), .C2(new_n691), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n683), .A2(KEYINPUT114), .A3(new_n783), .A4(new_n785), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n731), .A2(new_n788), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT52), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n702), .A2(new_n704), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n716), .A2(new_n725), .A3(new_n708), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n761), .A2(new_n608), .A3(new_n653), .ZN(new_n796));
  INV_X1    g610(.A(new_n634), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n598), .A2(new_n656), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n652), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n796), .B1(new_n799), .B2(new_n730), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n744), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n613), .A2(new_n598), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n802), .B1(new_n610), .B2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n803), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n700), .A2(new_n805), .A3(KEYINPUT113), .A4(new_n566), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n609), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n807), .A2(new_n629), .A3(new_n647), .A4(new_n600), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n801), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n795), .A2(new_n809), .A3(new_n742), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n782), .B1(new_n792), .B2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n731), .A2(new_n789), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n788), .A2(new_n790), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n813), .A2(new_n814), .A3(KEYINPUT52), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT52), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n791), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n698), .ZN(new_n819));
  AOI22_X1  g633(.A1(new_n819), .A2(new_n636), .B1(new_n721), .B2(new_n724), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n742), .A2(new_n705), .A3(new_n716), .A4(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n801), .A2(new_n808), .A3(new_n782), .ZN(new_n824));
  INV_X1    g638(.A(new_n794), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n825), .A2(KEYINPUT115), .A3(new_n705), .A4(new_n742), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n818), .A2(new_n823), .A3(new_n824), .A4(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n811), .A2(new_n812), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT116), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT116), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n811), .A2(new_n827), .A3(new_n830), .A4(new_n812), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n821), .A2(new_n801), .A3(new_n808), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n832), .A2(new_n818), .A3(KEYINPUT53), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n811), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT54), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n829), .A2(new_n831), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT51), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n668), .A2(new_n672), .A3(new_n699), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n562), .B1(new_n764), .B2(new_n765), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n720), .A2(new_n424), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n839), .A2(new_n840), .A3(new_n697), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n838), .A2(KEYINPUT50), .A3(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT50), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n668), .A2(new_n672), .A3(new_n699), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n839), .A2(new_n840), .A3(new_n697), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n837), .B1(new_n842), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n761), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n839), .A2(new_n840), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n722), .A2(new_n190), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n848), .B(new_n849), .C1(new_n777), .C2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n848), .A2(new_n697), .ZN(new_n852));
  NOR4_X1   g666(.A1(new_n852), .A2(new_n424), .A3(new_n562), .A4(new_n784), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n559), .A2(new_n624), .ZN(new_n854));
  INV_X1    g668(.A(new_n839), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n852), .A2(new_n855), .A3(new_n720), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n853), .A2(new_n854), .B1(new_n856), .B2(new_n646), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n847), .A2(new_n851), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n560), .A2(G953), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT50), .B1(new_n838), .B2(new_n841), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n844), .A2(new_n845), .A3(new_n843), .ZN(new_n862));
  OAI21_X1  g676(.A(KEYINPUT117), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT117), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n842), .A2(new_n864), .A3(new_n846), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n863), .A2(new_n851), .A3(new_n857), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(new_n837), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n860), .A2(new_n867), .ZN(new_n868));
  NOR4_X1   g682(.A1(new_n855), .A2(new_n852), .A3(new_n424), .A4(new_n652), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(KEYINPUT48), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n849), .A2(new_n714), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n853), .A2(new_n626), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n868), .A2(new_n871), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n781), .B1(new_n836), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n560), .A2(new_n272), .ZN(new_n876));
  AOI22_X1  g690(.A1(new_n828), .A2(KEYINPUT116), .B1(new_n834), .B2(KEYINPUT54), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n860), .A2(new_n867), .A3(new_n872), .A4(new_n873), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n878), .A2(new_n870), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n877), .A2(new_n879), .A3(KEYINPUT118), .A4(new_n831), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n875), .A2(new_n876), .A3(new_n880), .ZN(new_n881));
  NOR4_X1   g695(.A1(new_n784), .A2(new_n699), .A3(new_n190), .A4(new_n762), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n722), .B(KEYINPUT49), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n673), .A2(new_n425), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n881), .A2(new_n884), .ZN(G75));
  AOI21_X1  g699(.A(new_n283), .B1(new_n811), .B2(new_n827), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n298), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT56), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n371), .B(new_n355), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(KEYINPUT55), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n890), .B1(KEYINPUT119), .B2(KEYINPUT56), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n887), .A2(new_n888), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n891), .B1(new_n887), .B2(new_n888), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n272), .A2(G952), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(G51));
  NOR2_X1   g709(.A1(new_n292), .A2(new_n293), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT120), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n811), .A2(new_n827), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(KEYINPUT54), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n899), .A2(new_n828), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n750), .B(KEYINPUT57), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n897), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n749), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n886), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n894), .B1(new_n902), .B2(new_n904), .ZN(G54));
  NAND3_X1  g719(.A1(new_n886), .A2(KEYINPUT58), .A3(G475), .ZN(new_n906));
  INV_X1    g720(.A(new_n550), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n906), .A2(new_n907), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n908), .A2(new_n909), .A3(new_n894), .ZN(G60));
  OAI21_X1  g724(.A(new_n616), .B1(new_n620), .B2(new_n621), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(G478), .A2(G902), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(KEYINPUT59), .Z(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n912), .B1(new_n836), .B2(new_n915), .ZN(new_n916));
  AOI211_X1 g730(.A(new_n911), .B(new_n914), .C1(new_n899), .C2(new_n828), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n916), .A2(new_n894), .A3(new_n917), .ZN(G63));
  NAND2_X1  g732(.A1(G217), .A2(G902), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT60), .Z(new_n920));
  NAND3_X1  g734(.A1(new_n898), .A2(new_n644), .A3(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n894), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n921), .A2(KEYINPUT121), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(KEYINPUT61), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n898), .A2(new_n920), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n922), .B(new_n921), .C1(new_n925), .C2(new_n415), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n924), .B(new_n926), .ZN(G66));
  AOI21_X1  g741(.A(new_n272), .B1(new_n565), .B2(G224), .ZN(new_n928));
  OR3_X1    g742(.A1(new_n793), .A2(new_n794), .A3(new_n808), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n928), .B1(new_n929), .B2(new_n272), .ZN(new_n930));
  MUX2_X1   g744(.A(new_n928), .B(new_n930), .S(KEYINPUT122), .Z(new_n931));
  INV_X1    g745(.A(G898), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n371), .B1(new_n932), .B2(G953), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n931), .B(new_n933), .ZN(G69));
  INV_X1    g748(.A(new_n744), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n771), .A2(new_n813), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n935), .B1(new_n936), .B2(KEYINPUT125), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n760), .A2(new_n703), .A3(new_n783), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n938), .A2(new_n742), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT125), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n771), .A2(new_n813), .A3(new_n940), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n937), .A2(new_n779), .A3(new_n939), .A4(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n272), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n655), .A2(G953), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT126), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n539), .A2(new_n540), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n445), .B(new_n948), .Z(new_n949));
  NAND3_X1  g763(.A1(new_n943), .A2(KEYINPUT126), .A3(new_n944), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n947), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n687), .A2(new_n813), .ZN(new_n952));
  OR2_X1    g766(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n684), .B1(new_n627), .B2(new_n803), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n703), .A2(new_n734), .A3(new_n955), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n771), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g771(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n687), .A2(new_n813), .A3(new_n958), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n954), .A2(new_n779), .A3(new_n957), .A4(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n272), .ZN(new_n961));
  INV_X1    g775(.A(new_n949), .ZN(new_n962));
  AOI21_X1  g776(.A(KEYINPUT124), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT124), .ZN(new_n964));
  AOI211_X1 g778(.A(new_n964), .B(new_n949), .C1(new_n960), .C2(new_n272), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n272), .B1(G227), .B2(G900), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n951), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n967), .B1(new_n951), .B2(new_n966), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n968), .A2(new_n969), .ZN(G72));
  NAND2_X1  g784(.A1(G472), .A2(G902), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT63), .Z(new_n972));
  OAI21_X1  g786(.A(new_n972), .B1(new_n942), .B2(new_n929), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n973), .A2(new_n456), .A3(new_n449), .A4(new_n448), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT127), .ZN(new_n975));
  AND3_X1   g789(.A1(new_n974), .A2(new_n975), .A3(new_n922), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n975), .B1(new_n974), .B2(new_n922), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n972), .B1(new_n960), .B2(new_n929), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n978), .A2(new_n455), .A3(new_n450), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n677), .A2(new_n457), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n834), .A2(new_n972), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n976), .A2(new_n977), .A3(new_n982), .ZN(G57));
endmodule


