//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 1 0 1 1 0 1 0 1 1 1 0 1 1 0 0 0 0 0 0 1 0 0 1 0 0 1 0 0 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1319, new_n1320, new_n1321,
    new_n1322, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1392, new_n1393, new_n1394;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(G50), .B1(G58), .B2(G68), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT65), .Z(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G226), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n217), .B1(new_n202), .B2(new_n218), .ZN(new_n219));
  XOR2_X1   g0019(.A(KEYINPUT64), .B(G244), .Z(new_n220));
  AOI21_X1  g0020(.A(new_n219), .B1(G77), .B2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT66), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n216), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(new_n206), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n209), .B1(new_n213), .B2(new_n214), .C1(new_n225), .C2(KEYINPUT1), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n231), .B(new_n234), .Z(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XOR2_X1   g0036(.A(G107), .B(G116), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G58), .B(G77), .Z(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G351));
  NOR2_X1   g0042(.A1(G20), .A2(G33), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G50), .ZN(new_n244));
  INV_X1    g0044(.A(G77), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n211), .A2(G33), .ZN(new_n246));
  OAI221_X1 g0046(.A(new_n244), .B1(new_n211), .B2(G68), .C1(new_n245), .C2(new_n246), .ZN(new_n247));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n210), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(KEYINPUT11), .ZN(new_n251));
  INV_X1    g0051(.A(G1), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(KEYINPUT67), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT67), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G1), .ZN(new_n255));
  NAND4_X1  g0055(.A1(new_n253), .A2(new_n255), .A3(G13), .A4(G20), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G68), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n259), .B(KEYINPUT12), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT67), .B(G1), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n249), .B1(new_n261), .B2(G20), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G68), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n251), .A2(new_n260), .A3(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT14), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n210), .B1(G33), .B2(G41), .ZN(new_n266));
  INV_X1    g0066(.A(G41), .ZN(new_n267));
  INV_X1    g0067(.A(G45), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n266), .B1(new_n261), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G238), .ZN(new_n271));
  INV_X1    g0071(.A(G274), .ZN(new_n272));
  INV_X1    g0072(.A(new_n210), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G33), .A2(G41), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(G1), .B1(new_n267), .B2(new_n268), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n271), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n274), .A2(G1), .A3(G13), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT68), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT3), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(G33), .ZN(new_n282));
  INV_X1    g0082(.A(G33), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(KEYINPUT3), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n280), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(KEYINPUT3), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n281), .A2(G33), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n286), .A2(new_n287), .A3(KEYINPUT68), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G226), .A2(G1698), .ZN(new_n289));
  INV_X1    g0089(.A(G232), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n289), .B1(new_n290), .B2(G1698), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n285), .A2(new_n288), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G97), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n279), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(KEYINPUT13), .B1(new_n278), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NOR3_X1   g0096(.A1(new_n278), .A2(new_n294), .A3(KEYINPUT13), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n265), .B(G169), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n278), .ZN(new_n299));
  INV_X1    g0099(.A(new_n294), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT13), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n302), .A2(G179), .A3(new_n295), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n298), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n295), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n265), .B1(new_n305), .B2(G169), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n264), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G190), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G200), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n310), .B1(new_n302), .B2(new_n295), .ZN(new_n311));
  OR3_X1    g0111(.A1(new_n309), .A2(new_n264), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n248), .A2(new_n210), .ZN(new_n314));
  XNOR2_X1  g0114(.A(KEYINPUT8), .B(G58), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n316), .A2(new_n243), .B1(G20), .B2(G77), .ZN(new_n317));
  INV_X1    g0117(.A(G87), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT15), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT15), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G87), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n246), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n314), .B1(new_n317), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n262), .A2(G77), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(G77), .B2(new_n256), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n270), .A2(new_n220), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n277), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT69), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n285), .A2(new_n288), .ZN(new_n334));
  INV_X1    g0134(.A(G107), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n279), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(G232), .A2(G1698), .ZN(new_n337));
  INV_X1    g0137(.A(G238), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n337), .B1(new_n338), .B2(G1698), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n336), .B1(new_n334), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n330), .A2(KEYINPUT69), .A3(new_n277), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n333), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n329), .B1(new_n343), .B2(G190), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(G200), .ZN(new_n345));
  INV_X1    g0145(.A(G179), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G169), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n328), .B1(new_n342), .B2(new_n348), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n344), .A2(new_n345), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n316), .A2(new_n323), .B1(G150), .B2(new_n243), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n203), .A2(G20), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n314), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n262), .A2(G50), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(G50), .B2(new_n256), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n279), .B1(new_n334), .B2(new_n245), .ZN(new_n357));
  MUX2_X1   g0157(.A(G222), .B(G223), .S(G1698), .Z(new_n358));
  OAI21_X1  g0158(.A(new_n357), .B1(new_n334), .B2(new_n358), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n270), .A2(G226), .B1(new_n275), .B2(new_n276), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n356), .B1(new_n361), .B2(new_n348), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(G179), .B2(new_n361), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n356), .A2(KEYINPUT9), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT9), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(new_n353), .B2(new_n355), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n361), .A2(new_n308), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n310), .B1(new_n359), .B2(new_n360), .ZN(new_n369));
  NOR3_X1   g0169(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT10), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NOR4_X1   g0172(.A1(new_n367), .A2(new_n368), .A3(new_n369), .A4(KEYINPUT10), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n350), .B(new_n363), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT70), .ZN(new_n375));
  INV_X1    g0175(.A(new_n373), .ZN(new_n376));
  INV_X1    g0176(.A(new_n368), .ZN(new_n377));
  INV_X1    g0177(.A(new_n369), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n377), .A2(new_n378), .A3(new_n366), .A4(new_n364), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT10), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT70), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n381), .A2(new_n382), .A3(new_n363), .A4(new_n350), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n313), .B1(new_n375), .B2(new_n383), .ZN(new_n384));
  XNOR2_X1  g0184(.A(KEYINPUT3), .B(G33), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n218), .A2(G1698), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n385), .B(new_n386), .C1(G223), .C2(G1698), .ZN(new_n387));
  NAND2_X1  g0187(.A1(G33), .A2(G87), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n266), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n270), .A2(G232), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n390), .A2(G179), .A3(new_n277), .A4(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n261), .A2(new_n269), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n279), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n277), .B1(new_n394), .B2(new_n290), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n279), .B1(new_n387), .B2(new_n388), .ZN(new_n396));
  OAI21_X1  g0196(.A(G169), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n392), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G58), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n400), .A2(new_n258), .ZN(new_n401));
  OAI21_X1  g0201(.A(G20), .B1(new_n401), .B2(new_n201), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n243), .A2(G159), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT7), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(new_n385), .B2(G20), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n286), .A2(new_n287), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n407), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n404), .B1(new_n409), .B2(G68), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n314), .B1(new_n410), .B2(KEYINPUT16), .ZN(new_n411));
  AOI21_X1  g0211(.A(G20), .B1(new_n285), .B2(new_n288), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n408), .B1(new_n412), .B2(KEYINPUT7), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n404), .B1(new_n413), .B2(G68), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n411), .B1(new_n414), .B2(KEYINPUT16), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n256), .A2(new_n315), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n416), .B1(new_n262), .B2(new_n315), .ZN(new_n417));
  XNOR2_X1  g0217(.A(new_n417), .B(KEYINPUT71), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n399), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT18), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT72), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n415), .A2(new_n418), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n423), .A2(KEYINPUT72), .A3(KEYINPUT18), .A4(new_n398), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT18), .ZN(new_n425));
  XOR2_X1   g0225(.A(new_n417), .B(KEYINPUT71), .Z(new_n426));
  INV_X1    g0226(.A(new_n404), .ZN(new_n427));
  AOI211_X1 g0227(.A(new_n405), .B(G20), .C1(new_n286), .C2(new_n287), .ZN(new_n428));
  AND3_X1   g0228(.A1(new_n286), .A2(new_n287), .A3(KEYINPUT68), .ZN(new_n429));
  AOI21_X1  g0229(.A(KEYINPUT68), .B1(new_n286), .B2(new_n287), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n211), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n428), .B1(new_n431), .B2(new_n405), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n427), .B1(new_n432), .B2(new_n258), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT16), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n426), .B1(new_n435), .B2(new_n411), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n425), .B1(new_n436), .B2(new_n399), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n422), .A2(new_n424), .A3(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n310), .B1(new_n395), .B2(new_n396), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n390), .A2(new_n277), .A3(new_n391), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n439), .B1(new_n440), .B2(G190), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n415), .A2(new_n418), .A3(new_n441), .ZN(new_n442));
  XNOR2_X1  g0242(.A(new_n442), .B(KEYINPUT17), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n438), .A2(KEYINPUT73), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n437), .A2(new_n424), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT72), .B1(new_n419), .B2(KEYINPUT18), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n443), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT73), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n384), .A2(new_n444), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT5), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n268), .B1(new_n452), .B2(G41), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT74), .B1(new_n452), .B2(G41), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT74), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n455), .A2(new_n267), .A3(KEYINPUT5), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n261), .A2(new_n453), .A3(new_n454), .A4(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n279), .A2(G274), .ZN(new_n458));
  OAI21_X1  g0258(.A(KEYINPUT75), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n452), .A2(G41), .ZN(new_n460));
  AND4_X1   g0260(.A1(G45), .A2(new_n253), .A3(new_n255), .A4(new_n460), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n454), .A2(new_n456), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT75), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n461), .A2(new_n462), .A3(new_n463), .A4(new_n275), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n459), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G303), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n466), .B1(new_n285), .B2(new_n288), .ZN(new_n467));
  INV_X1    g0267(.A(G257), .ZN(new_n468));
  INV_X1    g0268(.A(G1698), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OR2_X1    g0270(.A1(new_n469), .A2(G264), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n385), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n266), .B1(new_n467), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n266), .B1(new_n461), .B2(new_n462), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G270), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n465), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(G116), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n248), .A2(new_n210), .B1(G20), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G283), .ZN(new_n480));
  INV_X1    g0280(.A(G97), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n480), .B(new_n211), .C1(G33), .C2(new_n481), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n479), .A2(KEYINPUT20), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(KEYINPUT20), .B1(new_n479), .B2(new_n482), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n253), .A2(new_n255), .A3(G33), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n256), .A2(new_n486), .A3(G116), .A4(new_n314), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n261), .A2(G13), .A3(G20), .A4(new_n478), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OR2_X1    g0289(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n477), .A2(new_n490), .A3(KEYINPUT21), .A4(G169), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(KEYINPUT78), .ZN(new_n492));
  OAI21_X1  g0292(.A(G169), .B1(new_n485), .B2(new_n489), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT78), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n494), .A2(new_n477), .A3(new_n495), .A4(KEYINPUT21), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n457), .A2(G264), .A3(new_n279), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G294), .ZN(new_n499));
  INV_X1    g0299(.A(G250), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n469), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n468), .A2(G1698), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n499), .B1(new_n407), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n266), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n465), .A2(new_n498), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n346), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n506), .A2(new_n348), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n318), .A2(KEYINPUT22), .A3(G20), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n285), .A2(new_n288), .A3(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n286), .A2(new_n287), .A3(new_n211), .A4(G87), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(KEYINPUT22), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT23), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(new_n211), .B2(G107), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n335), .A2(KEYINPUT23), .A3(G20), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n323), .A2(G116), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  XOR2_X1   g0319(.A(KEYINPUT80), .B(KEYINPUT24), .Z(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n520), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n514), .A2(new_n522), .A3(new_n518), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n314), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n249), .B1(new_n261), .B2(G33), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n525), .A2(G107), .A3(new_n256), .ZN(new_n526));
  XOR2_X1   g0326(.A(KEYINPUT81), .B(KEYINPUT25), .Z(new_n527));
  NAND3_X1  g0327(.A1(new_n257), .A2(new_n335), .A3(new_n527), .ZN(new_n528));
  OAI211_X1 g0328(.A(KEYINPUT81), .B(KEYINPUT25), .C1(new_n256), .C2(G107), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n526), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n508), .B(new_n509), .C1(new_n524), .C2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n494), .A2(new_n477), .ZN(new_n532));
  XOR2_X1   g0332(.A(KEYINPUT79), .B(KEYINPUT21), .Z(new_n533));
  OAI21_X1  g0333(.A(G303), .B1(new_n429), .B2(new_n430), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n472), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n346), .B1(new_n535), .B2(new_n266), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n464), .A2(new_n459), .B1(new_n475), .B2(G270), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n532), .A2(new_n533), .B1(new_n538), .B2(new_n490), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n497), .A2(new_n531), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n507), .A2(G190), .ZN(new_n541));
  INV_X1    g0341(.A(new_n523), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n522), .B1(new_n514), .B2(new_n518), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n249), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n530), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n505), .A2(new_n498), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n310), .B1(new_n546), .B2(new_n465), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n541), .A2(new_n544), .A3(new_n545), .A4(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n490), .B1(new_n477), .B2(G200), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n537), .A2(G190), .A3(new_n474), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n525), .A2(G97), .A3(new_n256), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n257), .A2(new_n481), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n335), .A2(KEYINPUT6), .A3(G97), .ZN(new_n557));
  XOR2_X1   g0357(.A(G97), .B(G107), .Z(new_n558));
  OAI21_X1  g0358(.A(new_n557), .B1(new_n558), .B2(KEYINPUT6), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n559), .A2(G20), .B1(G77), .B2(new_n243), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n432), .B2(new_n335), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n556), .B1(new_n561), .B2(new_n249), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n469), .A2(G244), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT4), .ZN(new_n564));
  OAI22_X1  g0364(.A1(new_n563), .A2(new_n564), .B1(new_n500), .B2(new_n469), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n285), .A2(new_n288), .A3(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n480), .ZN(new_n567));
  INV_X1    g0367(.A(G244), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n568), .A2(G1698), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n569), .A2(new_n286), .A3(new_n287), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n567), .B1(new_n570), .B2(new_n564), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n266), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n475), .A2(G257), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(new_n465), .A3(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n575), .A2(G190), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n464), .A2(new_n459), .B1(new_n475), .B2(G257), .ZN(new_n577));
  AOI21_X1  g0377(.A(G200), .B1(new_n577), .B2(new_n573), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n562), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n577), .A2(new_n346), .A3(new_n573), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n575), .A2(new_n348), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n413), .A2(G107), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n314), .B1(new_n582), .B2(new_n560), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n580), .B(new_n581), .C1(new_n583), .C2(new_n556), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT76), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n579), .A2(new_n584), .A3(KEYINPUT76), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n338), .A2(new_n469), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n568), .A2(G1698), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n286), .A2(new_n589), .A3(new_n287), .A4(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n283), .A2(new_n478), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n266), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n261), .A2(new_n279), .A3(G45), .A4(G274), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n253), .A2(new_n255), .A3(G45), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n597), .A2(G250), .A3(new_n279), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n595), .A2(G190), .A3(new_n596), .A4(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n596), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n279), .B1(new_n591), .B2(new_n593), .ZN(new_n601));
  OAI21_X1  g0401(.A(G200), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT19), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n211), .B1(new_n293), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n318), .A2(new_n481), .A3(new_n335), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n286), .A2(new_n287), .A3(new_n211), .A4(G68), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n603), .B1(new_n246), .B2(new_n481), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  XNOR2_X1  g0409(.A(KEYINPUT15), .B(G87), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n609), .A2(new_n249), .B1(new_n257), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n525), .A2(G87), .A3(new_n256), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n599), .A2(new_n602), .A3(new_n611), .A4(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n609), .A2(new_n249), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n322), .A2(KEYINPUT77), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT77), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n525), .A2(new_n256), .A3(new_n615), .A4(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n257), .A2(new_n610), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n614), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n595), .A2(new_n346), .A3(new_n596), .A4(new_n598), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n348), .B1(new_n600), .B2(new_n601), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n613), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n587), .A2(new_n588), .A3(new_n625), .ZN(new_n626));
  NOR4_X1   g0426(.A1(new_n451), .A2(new_n540), .A3(new_n553), .A4(new_n626), .ZN(G372));
  INV_X1    g0427(.A(new_n363), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n420), .A2(new_n437), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n347), .A2(new_n349), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n307), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n443), .A2(new_n312), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n628), .B1(new_n633), .B2(new_n381), .ZN(new_n634));
  INV_X1    g0434(.A(new_n585), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n524), .A2(new_n530), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n547), .B1(new_n507), .B2(G190), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n624), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n540), .A2(new_n635), .A3(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT26), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(new_n584), .B2(new_n624), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n575), .A2(G179), .ZN(new_n642));
  AOI21_X1  g0442(.A(G169), .B1(new_n577), .B2(new_n573), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n562), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n644), .A2(new_n645), .A3(new_n625), .A4(KEYINPUT26), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(KEYINPUT82), .B1(new_n647), .B2(new_n623), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT82), .ZN(new_n649));
  INV_X1    g0449(.A(new_n623), .ZN(new_n650));
  AOI211_X1 g0450(.A(new_n649), .B(new_n650), .C1(new_n641), .C2(new_n646), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n639), .B1(new_n648), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n634), .B1(new_n451), .B2(new_n653), .ZN(G369));
  INV_X1    g0454(.A(G330), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n211), .A2(G13), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n261), .A2(new_n656), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n657), .A2(KEYINPUT27), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(KEYINPUT27), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(G213), .A3(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(G343), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n490), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n497), .A2(new_n539), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n663), .B1(new_n497), .B2(new_n539), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n552), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(KEYINPUT83), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT83), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n668), .B(new_n552), .C1(new_n664), .C2(new_n665), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n655), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n531), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n662), .B1(new_n524), .B2(new_n530), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT84), .ZN(new_n674));
  AOI22_X1  g0474(.A1(new_n673), .A2(new_n674), .B1(new_n636), .B2(new_n637), .ZN(new_n675));
  INV_X1    g0475(.A(new_n662), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n676), .B1(new_n544), .B2(new_n545), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(KEYINPUT84), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n672), .B1(new_n675), .B2(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n531), .A2(new_n662), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n671), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n549), .B1(new_n677), .B2(KEYINPUT84), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n673), .A2(new_n674), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n531), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n490), .A2(new_n536), .A3(new_n537), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n493), .B1(new_n537), .B2(new_n474), .ZN(new_n689));
  INV_X1    g0489(.A(new_n533), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(new_n492), .B2(new_n496), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(new_n662), .ZN(new_n693));
  AOI211_X1 g0493(.A(KEYINPUT85), .B(new_n680), .C1(new_n687), .C2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT85), .ZN(new_n695));
  INV_X1    g0495(.A(new_n680), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n687), .A2(new_n693), .A3(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n695), .B1(new_n697), .B2(new_n696), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n684), .B1(new_n694), .B2(new_n698), .ZN(G399));
  INV_X1    g0499(.A(new_n207), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G41), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n605), .A2(G116), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(G1), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n214), .B2(new_n702), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT28), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n652), .A2(new_n676), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT29), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n650), .B1(new_n641), .B2(new_n646), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n662), .B1(new_n639), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT29), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n505), .A2(new_n498), .ZN(new_n713));
  NOR2_X1   g0513(.A1(G238), .A2(G1698), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n714), .B1(new_n568), .B2(G1698), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n592), .B1(new_n715), .B2(new_n385), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n596), .B(new_n598), .C1(new_n716), .C2(new_n279), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  AND3_X1   g0518(.A1(new_n718), .A2(new_n537), .A3(new_n536), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n577), .A2(KEYINPUT30), .A3(new_n573), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT30), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n718), .A2(new_n537), .A3(new_n536), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n723), .B1(new_n724), .B2(new_n575), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n717), .A2(new_n346), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n575), .A2(new_n477), .A3(new_n506), .A4(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n722), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(KEYINPUT31), .B1(new_n728), .B2(new_n662), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n725), .A2(new_n727), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(KEYINPUT86), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT86), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n725), .A2(new_n732), .A3(new_n727), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n731), .A2(new_n722), .A3(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT31), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n676), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n729), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT87), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n736), .ZN(new_n740));
  AOI22_X1  g0540(.A1(new_n730), .A2(KEYINPUT86), .B1(new_n719), .B2(new_n721), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n740), .B1(new_n741), .B2(new_n733), .ZN(new_n742));
  OAI21_X1  g0542(.A(KEYINPUT87), .B1(new_n742), .B2(new_n729), .ZN(new_n743));
  AND3_X1   g0543(.A1(new_n579), .A2(new_n584), .A3(KEYINPUT76), .ZN(new_n744));
  AOI21_X1  g0544(.A(KEYINPUT76), .B1(new_n579), .B2(new_n584), .ZN(new_n745));
  NOR3_X1   g0545(.A1(new_n744), .A2(new_n745), .A3(new_n624), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n540), .A2(new_n553), .A3(new_n662), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n739), .A2(new_n743), .A3(new_n748), .ZN(new_n749));
  AOI22_X1  g0549(.A1(new_n709), .A2(new_n712), .B1(G330), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n706), .B1(new_n750), .B2(G1), .ZN(G364));
  NAND3_X1  g0551(.A1(new_n667), .A2(new_n655), .A3(new_n669), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n252), .B1(new_n656), .B2(G45), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n671), .B(new_n752), .C1(new_n701), .C2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G13), .A2(G33), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n666), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n210), .B1(G20), .B2(new_n348), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n211), .A2(new_n346), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT89), .ZN(new_n763));
  AOI21_X1  g0563(.A(G200), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n764), .B1(new_n763), .B2(new_n762), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n308), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G179), .A2(G200), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n211), .B1(new_n767), .B2(G190), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT91), .Z(new_n769));
  AOI22_X1  g0569(.A1(new_n766), .A2(G58), .B1(new_n769), .B2(G97), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n765), .A2(G190), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n770), .B1(new_n245), .B2(new_n772), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n762), .A2(G190), .A3(new_n310), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n762), .A2(new_n308), .A3(new_n310), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n774), .A2(G68), .B1(new_n775), .B2(G50), .ZN(new_n776));
  INV_X1    g0576(.A(new_n334), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n310), .A2(G179), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n778), .A2(G20), .A3(G190), .ZN(new_n779));
  OAI211_X1 g0579(.A(new_n776), .B(new_n777), .C1(new_n318), .C2(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n778), .A2(G20), .A3(new_n308), .ZN(new_n781));
  OR2_X1    g0581(.A1(new_n781), .A2(KEYINPUT90), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(KEYINPUT90), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G107), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n767), .A2(G20), .A3(new_n308), .ZN(new_n787));
  INV_X1    g0587(.A(G159), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT32), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n773), .A2(new_n780), .A3(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(KEYINPUT33), .A2(G317), .ZN(new_n793));
  AND2_X1   g0593(.A1(KEYINPUT33), .A2(G317), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n774), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(G311), .A2(new_n771), .B1(new_n766), .B2(G322), .ZN(new_n796));
  INV_X1    g0596(.A(new_n768), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n775), .A2(G326), .B1(new_n797), .B2(G294), .ZN(new_n798));
  INV_X1    g0598(.A(new_n787), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G329), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n334), .B(new_n800), .C1(new_n466), .C2(new_n779), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(new_n785), .B2(G283), .ZN(new_n802));
  AND4_X1   g0602(.A1(new_n795), .A2(new_n796), .A3(new_n798), .A4(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n760), .B1(new_n792), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n754), .A2(new_n701), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT88), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n777), .A2(G355), .A3(new_n207), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n241), .A2(new_n268), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n700), .A2(new_n385), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(G45), .B2(new_n214), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n808), .B1(G116), .B2(new_n207), .C1(new_n809), .C2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n758), .A2(new_n760), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n807), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n759), .A2(new_n804), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n755), .A2(new_n815), .ZN(G396));
  NAND3_X1  g0616(.A1(new_n347), .A2(new_n349), .A3(new_n676), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n344), .A2(new_n345), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n328), .B2(new_n676), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n818), .B1(new_n820), .B2(new_n630), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n707), .B(new_n821), .ZN(new_n822));
  AND2_X1   g0622(.A1(new_n749), .A2(G330), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT94), .Z(new_n825));
  OAI221_X1 g0625(.A(new_n825), .B1(new_n701), .B2(new_n754), .C1(new_n823), .C2(new_n822), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n760), .A2(new_n756), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n807), .B1(new_n245), .B2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(G132), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n385), .B1(new_n787), .B2(new_n829), .C1(new_n779), .C2(new_n202), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n784), .A2(new_n258), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n830), .B(new_n831), .C1(G58), .C2(new_n797), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT93), .Z(new_n833));
  AOI22_X1  g0633(.A1(new_n774), .A2(G150), .B1(new_n775), .B2(G137), .ZN(new_n834));
  INV_X1    g0634(.A(new_n766), .ZN(new_n835));
  XNOR2_X1  g0635(.A(KEYINPUT92), .B(G143), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n834), .B1(new_n835), .B2(new_n836), .C1(new_n788), .C2(new_n772), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT34), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n775), .A2(G303), .B1(G311), .B2(new_n799), .ZN(new_n839));
  INV_X1    g0639(.A(G283), .ZN(new_n840));
  INV_X1    g0640(.A(new_n774), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n839), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(G87), .B2(new_n785), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n334), .B1(new_n335), .B2(new_n779), .ZN(new_n844));
  INV_X1    g0644(.A(G294), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n478), .A2(new_n772), .B1(new_n835), .B2(new_n845), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n844), .B(new_n846), .C1(G97), .C2(new_n769), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n833), .A2(new_n838), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n760), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n828), .B1(new_n848), .B2(new_n849), .C1(new_n757), .C2(new_n821), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n826), .A2(new_n850), .ZN(G384));
  NOR2_X1   g0651(.A1(new_n261), .A2(new_n656), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n728), .A2(new_n736), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n636), .A2(new_n637), .B1(new_n551), .B2(new_n550), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n692), .A2(new_n854), .A3(new_n531), .A4(new_n676), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n853), .B1(new_n626), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n575), .ZN(new_n857));
  AOI21_X1  g0657(.A(KEYINPUT30), .B1(new_n719), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n477), .A2(new_n506), .A3(new_n726), .ZN(new_n859));
  OAI22_X1  g0659(.A1(new_n859), .A2(new_n857), .B1(new_n724), .B2(new_n720), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n662), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(KEYINPUT97), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT97), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n728), .A2(new_n863), .A3(new_n662), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n862), .A2(new_n735), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(KEYINPUT98), .ZN(new_n866));
  AOI21_X1  g0666(.A(KEYINPUT31), .B1(new_n861), .B2(KEYINPUT97), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT98), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n867), .A2(new_n868), .A3(new_n864), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n856), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n264), .A2(new_n662), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n313), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n307), .A2(new_n312), .A3(new_n871), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n821), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT99), .ZN(new_n877));
  NOR3_X1   g0677(.A1(new_n870), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n821), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(new_n874), .B2(new_n873), .ZN(new_n880));
  INV_X1    g0680(.A(new_n853), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n881), .B1(new_n746), .B2(new_n747), .ZN(new_n882));
  AND4_X1   g0682(.A1(new_n868), .A2(new_n862), .A3(new_n735), .A4(new_n864), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n868), .B1(new_n867), .B2(new_n864), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT99), .B1(new_n880), .B2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n878), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT95), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n442), .B1(new_n436), .B2(new_n399), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT37), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n436), .B2(new_n660), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT7), .B1(new_n407), .B2(new_n211), .ZN(new_n893));
  OAI21_X1  g0693(.A(G68), .B1(new_n893), .B2(new_n428), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n894), .A2(KEYINPUT16), .A3(new_n427), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n249), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n410), .A2(KEYINPUT16), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n417), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n392), .A2(new_n397), .A3(new_n660), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n890), .B1(new_n442), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n888), .B1(new_n892), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n423), .A2(new_n398), .ZN(new_n903));
  INV_X1    g0703(.A(new_n660), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n896), .B1(new_n434), .B2(new_n433), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n904), .B1(new_n905), .B2(new_n426), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n903), .A2(new_n906), .A3(new_n890), .A4(new_n442), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n442), .A2(new_n900), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT37), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n907), .A2(KEYINPUT95), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n902), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n898), .A2(new_n904), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n447), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT38), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n907), .A2(KEYINPUT95), .A3(new_n909), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT95), .B1(new_n907), .B2(new_n909), .ZN(new_n918));
  OAI21_X1  g0718(.A(KEYINPUT38), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n912), .B1(new_n438), .B2(new_n443), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT96), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT38), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(new_n902), .B2(new_n910), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT96), .B1(new_n924), .B2(new_n914), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n916), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT40), .B1(new_n887), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n906), .B1(new_n443), .B2(new_n629), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n903), .A2(new_n906), .A3(new_n442), .ZN(new_n929));
  AND3_X1   g0729(.A1(new_n415), .A2(new_n418), .A3(new_n441), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n930), .A2(new_n419), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT37), .B1(new_n423), .B2(new_n904), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n929), .A2(KEYINPUT37), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n923), .B1(new_n928), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT100), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n934), .B(new_n935), .C1(new_n919), .C2(new_n920), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n911), .A2(new_n914), .A3(KEYINPUT38), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n935), .B1(new_n938), .B2(new_n934), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT40), .ZN(new_n941));
  NOR3_X1   g0741(.A1(new_n870), .A2(new_n941), .A3(new_n876), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n927), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n451), .A2(new_n870), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n655), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n943), .B2(new_n944), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n629), .A2(new_n904), .ZN(new_n947));
  INV_X1    g0747(.A(new_n875), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n652), .A2(new_n676), .A3(new_n821), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n948), .B1(new_n949), .B2(new_n817), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n947), .B1(new_n926), .B2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT39), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n938), .A2(new_n952), .A3(new_n934), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n926), .B2(KEYINPUT39), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n307), .A2(new_n662), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n951), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n450), .A2(new_n709), .A3(new_n712), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n634), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n957), .B(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n852), .B1(new_n946), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n960), .B2(new_n946), .ZN(new_n962));
  AOI211_X1 g0762(.A(new_n478), .B(new_n213), .C1(new_n559), .C2(KEYINPUT35), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(KEYINPUT35), .B2(new_n559), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT36), .Z(new_n965));
  OAI21_X1  g0765(.A(G77), .B1(new_n400), .B2(new_n258), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n966), .A2(new_n214), .B1(G50), .B2(new_n258), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n261), .A2(G13), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n965), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n962), .A2(new_n969), .ZN(G367));
  NOR2_X1   g0770(.A1(new_n768), .A2(new_n335), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n779), .A2(new_n478), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT46), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n971), .B(new_n973), .C1(G311), .C2(new_n775), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n785), .A2(G97), .ZN(new_n975));
  INV_X1    g0775(.A(G317), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n407), .B1(new_n787), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(new_n774), .B2(G294), .ZN(new_n978));
  AOI22_X1  g0778(.A1(G283), .A2(new_n771), .B1(new_n766), .B2(G303), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n974), .A2(new_n975), .A3(new_n978), .A4(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n784), .A2(new_n245), .ZN(new_n981));
  INV_X1    g0781(.A(G137), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n777), .B1(new_n400), .B2(new_n779), .C1(new_n982), .C2(new_n787), .ZN(new_n983));
  INV_X1    g0783(.A(new_n836), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n981), .B(new_n983), .C1(new_n775), .C2(new_n984), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n772), .A2(new_n202), .B1(new_n788), .B2(new_n841), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT106), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n766), .A2(G150), .B1(new_n769), .B2(G68), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n985), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n986), .A2(new_n987), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n980), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT47), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n760), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n234), .A2(new_n810), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n760), .B(new_n758), .C1(new_n700), .C2(new_n322), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n807), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n758), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n611), .A2(new_n612), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n662), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n650), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1002), .A2(KEYINPUT101), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1002), .B(KEYINPUT101), .C1(new_n624), .C2(new_n1001), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n994), .B(new_n997), .C1(new_n998), .C2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n635), .B1(new_n562), .B2(new_n676), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n644), .A2(new_n645), .A3(new_n662), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n698), .B2(new_n694), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT45), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI211_X1 g0813(.A(KEYINPUT45), .B(new_n1010), .C1(new_n698), .C2(new_n694), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n692), .A2(new_n662), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n696), .B1(new_n1016), .B2(new_n679), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(KEYINPUT85), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n697), .A2(new_n695), .A3(new_n696), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1010), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT44), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1018), .A2(new_n1019), .A3(KEYINPUT44), .A4(new_n1020), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n684), .B1(new_n1015), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n682), .A2(new_n1016), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n670), .A2(KEYINPUT104), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT104), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n1030), .B(new_n655), .C1(new_n667), .C2(new_n669), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n697), .B(new_n1028), .C1(new_n1029), .C2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1028), .A2(new_n697), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n671), .B2(new_n1030), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1032), .A2(new_n750), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT105), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1015), .A2(new_n1025), .A3(new_n684), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1032), .A2(new_n750), .A3(KEYINPUT105), .A4(new_n1034), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1027), .A2(new_n1037), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n750), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n701), .B(new_n1042), .Z(new_n1043));
  AOI21_X1  g0843(.A(new_n754), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n681), .A2(new_n693), .A3(new_n1010), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n584), .B1(new_n1008), .B2(new_n531), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n1045), .A2(KEYINPUT42), .B1(new_n676), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(KEYINPUT42), .B2(new_n1045), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT43), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1048), .B1(new_n1049), .B2(new_n1005), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1006), .A2(KEYINPUT43), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n683), .A2(new_n1010), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n1050), .A2(new_n1051), .B1(KEYINPUT102), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n1051), .B2(new_n1050), .ZN(new_n1054));
  OR2_X1    g0854(.A1(new_n1052), .A2(KEYINPUT102), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1054), .B(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1007), .B1(new_n1044), .B2(new_n1056), .ZN(G387));
  NAND3_X1  g0857(.A1(new_n1032), .A2(new_n754), .A3(new_n1034), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n385), .B1(new_n799), .B2(G326), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n779), .A2(new_n845), .B1(new_n768), .B2(new_n840), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n774), .A2(G311), .B1(new_n775), .B2(G322), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1061), .B1(new_n835), .B2(new_n976), .C1(new_n466), .C2(new_n772), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT48), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1060), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n1063), .B2(new_n1062), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT49), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1059), .B1(new_n478), .B2(new_n784), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n779), .A2(new_n245), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n407), .B(new_n1069), .C1(G150), .C2(new_n799), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G159), .A2(new_n775), .B1(new_n774), .B2(new_n316), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n975), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n615), .A2(new_n617), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n769), .A2(new_n1074), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1075), .B1(new_n835), .B2(new_n202), .C1(new_n258), .C2(new_n772), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n1067), .A2(new_n1068), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n760), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n315), .A2(G50), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT50), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n268), .B1(new_n258), .B2(new_n245), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n703), .B2(KEYINPUT107), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1080), .B(new_n1082), .C1(KEYINPUT107), .C2(new_n703), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1083), .B(new_n810), .C1(new_n231), .C2(new_n268), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n777), .A2(new_n207), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1084), .B1(G107), .B2(new_n207), .C1(new_n703), .C2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n807), .B1(new_n1086), .B2(new_n813), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1078), .B(new_n1087), .C1(new_n681), .C2(new_n998), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1035), .A2(new_n701), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n750), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1058), .B(new_n1088), .C1(new_n1089), .C2(new_n1090), .ZN(G393));
  NAND3_X1  g0891(.A1(new_n1027), .A2(new_n754), .A3(new_n1038), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n813), .B1(new_n481), .B2(new_n207), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n238), .B2(new_n810), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n766), .A2(G311), .B1(G317), .B2(new_n775), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT52), .Z(new_n1096));
  INV_X1    g0896(.A(new_n779), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1097), .A2(G283), .B1(new_n799), .B2(G322), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n774), .A2(G303), .B1(new_n797), .B2(G116), .ZN(new_n1099));
  AND4_X1   g0899(.A1(new_n334), .A2(new_n786), .A3(new_n1098), .A4(new_n1099), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1096), .B(new_n1100), .C1(new_n845), .C2(new_n772), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n766), .A2(G159), .B1(G150), .B2(new_n775), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT108), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(KEYINPUT51), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n769), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1105), .A2(new_n245), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n385), .B1(new_n836), .B2(new_n787), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(G68), .B2(new_n1097), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n1108), .B1(new_n841), .B2(new_n202), .C1(new_n784), .C2(new_n318), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1106), .B(new_n1109), .C1(new_n316), .C2(new_n771), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1104), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1103), .A2(KEYINPUT51), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1101), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n807), .B(new_n1094), .C1(new_n1113), .C2(new_n760), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n1010), .B2(new_n998), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1092), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1038), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1035), .B1(new_n1117), .B2(new_n1026), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1040), .A2(new_n701), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(KEYINPUT109), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT109), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1040), .A2(new_n1118), .A3(new_n1121), .A4(new_n701), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1116), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(G390));
  NAND2_X1  g0924(.A1(new_n949), .A2(new_n817), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n875), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT110), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1126), .A2(new_n1127), .A3(new_n956), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n926), .A2(KEYINPUT39), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n956), .ZN(new_n1130));
  OAI21_X1  g0930(.A(KEYINPUT110), .B1(new_n950), .B2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1128), .A2(new_n1129), .A3(new_n1131), .A4(new_n953), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n938), .A2(new_n934), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(KEYINPUT100), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n936), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n820), .A2(new_n630), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n818), .B1(new_n711), .B2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n956), .B1(new_n1137), .B2(new_n948), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n749), .A2(G330), .A3(new_n875), .A4(new_n821), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1132), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1127), .B1(new_n1126), .B2(new_n956), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n921), .B1(new_n919), .B2(new_n920), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n924), .A2(KEYINPUT96), .A3(new_n914), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n915), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n953), .B1(new_n1146), .B2(new_n952), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1143), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1139), .B1(new_n1148), .B2(new_n1128), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n866), .A2(new_n869), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n655), .B1(new_n1150), .B2(new_n882), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n880), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1142), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n748), .B1(new_n737), .B2(new_n738), .ZN(new_n1154));
  NOR3_X1   g0954(.A1(new_n742), .A2(KEYINPUT87), .A3(new_n729), .ZN(new_n1155));
  OAI211_X1 g0955(.A(G330), .B(new_n821), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n948), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n1152), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1137), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n885), .A2(G330), .A3(new_n821), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1159), .B1(new_n1160), .B2(new_n948), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n1158), .A2(new_n1125), .B1(new_n1161), .B2(new_n1141), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT111), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n450), .A2(new_n1151), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n958), .A2(new_n634), .A3(new_n1164), .ZN(new_n1165));
  NOR3_X1   g0965(.A1(new_n1162), .A2(new_n1163), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1160), .A2(new_n948), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1167), .A2(new_n1137), .A3(new_n1141), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1125), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n948), .A2(new_n1156), .B1(new_n1151), .B2(new_n880), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1168), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n958), .A2(new_n634), .A3(new_n1164), .ZN(new_n1172));
  AOI21_X1  g0972(.A(KEYINPUT111), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1166), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n702), .B1(new_n1153), .B2(new_n1174), .ZN(new_n1175));
  AND3_X1   g0975(.A1(new_n1132), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1152), .B1(new_n1132), .B2(new_n1140), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1163), .B1(new_n1162), .B2(new_n1165), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1171), .A2(new_n1172), .A3(KEYINPUT111), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1178), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1175), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n955), .A2(new_n756), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n827), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n775), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n841), .A2(new_n335), .B1(new_n1187), .B2(new_n840), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n779), .A2(new_n318), .B1(new_n845), .B2(new_n787), .ZN(new_n1189));
  OR4_X1    g0989(.A1(new_n777), .A2(new_n1188), .A3(new_n831), .A4(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1106), .B1(G116), .B2(new_n766), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n1191), .B(KEYINPUT112), .Z(new_n1192));
  AOI211_X1 g0992(.A(new_n1190), .B(new_n1192), .C1(G97), .C2(new_n771), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT113), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(G128), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n841), .A2(new_n982), .B1(new_n1187), .B2(new_n1196), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n334), .B(new_n1197), .C1(G125), .C2(new_n799), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT53), .ZN(new_n1199));
  INV_X1    g0999(.A(G150), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1199), .B1(new_n779), .B2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1097), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n785), .A2(G50), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n766), .A2(G132), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(KEYINPUT54), .B(G143), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n771), .A2(new_n1206), .B1(new_n769), .B2(G159), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1198), .A2(new_n1203), .A3(new_n1204), .A4(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1195), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n1194), .B2(new_n1193), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n806), .B1(new_n316), .B2(new_n1186), .C1(new_n1210), .C2(new_n849), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n1153), .A2(new_n753), .B1(new_n1185), .B2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1183), .A2(new_n1213), .ZN(G378));
  INV_X1    g1014(.A(KEYINPUT118), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n655), .B1(new_n940), .B2(new_n942), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n877), .B1(new_n870), .B2(new_n876), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n880), .A2(new_n885), .A3(KEYINPUT99), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n941), .B1(new_n1219), .B2(new_n1146), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n381), .A2(new_n363), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n356), .A2(new_n660), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1221), .B(new_n1222), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1223), .B(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n1216), .A2(new_n1220), .A3(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1226), .B1(new_n1216), .B2(new_n1220), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(new_n1227), .A2(new_n1228), .A3(new_n957), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n1126), .A2(new_n1146), .B1(new_n629), .B2(new_n904), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n1130), .B2(new_n1147), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n942), .ZN(new_n1232));
  OAI21_X1  g1032(.A(G330), .B1(new_n1135), .B2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1225), .B1(new_n927), .B2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1216), .A2(new_n1220), .A3(new_n1226), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1231), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1215), .B1(new_n1229), .B2(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n957), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1234), .A2(new_n1231), .A3(new_n1235), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1238), .A2(KEYINPUT118), .A3(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1237), .A2(new_n754), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1225), .A2(new_n756), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n805), .B1(G50), .B2(new_n1186), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n841), .A2(new_n481), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n385), .A2(G41), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n787), .A2(new_n840), .ZN(new_n1247));
  NOR4_X1   g1047(.A1(new_n1244), .A2(new_n1069), .A3(new_n1246), .A4(new_n1247), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n1248), .B1(new_n335), .B2(new_n835), .C1(new_n1073), .C2(new_n772), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n769), .A2(G68), .B1(G116), .B2(new_n775), .ZN(new_n1250));
  XOR2_X1   g1050(.A(new_n1250), .B(KEYINPUT115), .Z(new_n1251));
  NOR2_X1   g1051(.A1(new_n784), .A2(new_n400), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(new_n1252), .B(KEYINPUT114), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(new_n1249), .A2(new_n1251), .A3(new_n1253), .ZN(new_n1254));
  XOR2_X1   g1054(.A(new_n1254), .B(KEYINPUT58), .Z(new_n1255));
  OAI211_X1 g1055(.A(new_n1246), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n775), .A2(G125), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n774), .A2(G132), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1097), .A2(new_n1206), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1257), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n835), .A2(new_n1196), .B1(new_n1200), .B2(new_n1105), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n1260), .B(new_n1261), .C1(G137), .C2(new_n771), .ZN(new_n1262));
  XOR2_X1   g1062(.A(KEYINPUT116), .B(KEYINPUT59), .Z(new_n1263));
  NOR2_X1   g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1265));
  AOI211_X1 g1065(.A(G33), .B(G41), .C1(new_n799), .C2(G124), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1265), .B(new_n1266), .C1(new_n788), .C2(new_n784), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1255), .B(new_n1256), .C1(new_n1264), .C2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1243), .B1(new_n1268), .B2(new_n760), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1242), .A2(new_n1269), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(new_n1270), .B(KEYINPUT117), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1241), .A2(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1172), .B1(new_n1153), .B2(new_n1174), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1273), .A2(new_n1237), .A3(new_n1240), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT57), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n702), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT119), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1165), .B1(new_n1178), .B2(new_n1181), .ZN(new_n1278));
  OAI21_X1  g1078(.A(KEYINPUT57), .B1(new_n1229), .B2(new_n1236), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1277), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1275), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1273), .A2(KEYINPUT119), .A3(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1280), .A2(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1272), .B1(new_n1276), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(G375));
  NAND2_X1  g1085(.A1(new_n948), .A2(new_n756), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n806), .B1(G68), .B2(new_n1186), .ZN(new_n1287));
  OAI22_X1  g1087(.A1(new_n841), .A2(new_n478), .B1(new_n1187), .B2(new_n845), .ZN(new_n1288));
  OAI22_X1  g1088(.A1(new_n779), .A2(new_n481), .B1(new_n466), .B2(new_n787), .ZN(new_n1289));
  NOR4_X1   g1089(.A1(new_n1288), .A2(new_n981), .A3(new_n777), .A4(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n766), .A2(G283), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n771), .A2(G107), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1290), .A2(new_n1075), .A3(new_n1291), .A4(new_n1292), .ZN(new_n1293));
  AOI22_X1  g1093(.A1(G132), .A2(new_n775), .B1(new_n774), .B2(new_n1206), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n385), .B1(new_n787), .B2(new_n1196), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1295), .B1(G159), .B2(new_n1097), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1296), .B1(new_n1105), .B2(new_n202), .ZN(new_n1297));
  AOI211_X1 g1097(.A(new_n1297), .B(new_n1253), .C1(G150), .C2(new_n771), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT120), .ZN(new_n1299));
  OAI221_X1 g1099(.A(new_n1294), .B1(new_n982), .B2(new_n835), .C1(new_n1298), .C2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1298), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1301), .A2(KEYINPUT120), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1293), .B1(new_n1300), .B2(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1287), .B1(new_n1303), .B2(new_n760), .ZN(new_n1304));
  AOI22_X1  g1104(.A1(new_n1171), .A2(new_n754), .B1(new_n1286), .B2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1174), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1043), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1305), .B1(new_n1307), .B2(new_n1308), .ZN(G381));
  NAND2_X1  g1109(.A1(G378), .A2(KEYINPUT121), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1212), .B1(new_n1182), .B2(new_n1175), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT121), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1310), .A2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  NOR4_X1   g1115(.A1(G387), .A2(G384), .A3(G396), .A4(G393), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(G390), .A2(G381), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1315), .A2(new_n1284), .A3(new_n1316), .A4(new_n1317), .ZN(G407));
  NAND2_X1  g1118(.A1(new_n661), .A2(G213), .ZN(new_n1319));
  XNOR2_X1  g1119(.A(new_n1319), .B(KEYINPUT122), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1315), .A2(new_n1284), .A3(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(G407), .A2(G213), .A3(new_n1321), .ZN(new_n1322));
  XNOR2_X1  g1122(.A(new_n1322), .B(KEYINPUT123), .ZN(G409));
  INV_X1    g1123(.A(new_n1007), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1056), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(new_n753), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1324), .B1(new_n1325), .B2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1328), .A2(G390), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT125), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1330), .B1(G387), .B2(new_n1123), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1329), .A2(new_n1331), .ZN(new_n1332));
  XOR2_X1   g1132(.A(G393), .B(G396), .Z(new_n1333));
  NAND3_X1  g1133(.A1(new_n1328), .A2(G390), .A3(new_n1330), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1332), .A2(new_n1333), .A3(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT126), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1336), .B1(new_n1328), .B2(G390), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1333), .B1(new_n1328), .B2(G390), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(G387), .A2(KEYINPUT126), .A3(new_n1123), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1337), .A2(new_n1338), .A3(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1335), .A2(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1341), .ZN(new_n1342));
  AOI211_X1 g1142(.A(new_n1311), .B(new_n1272), .C1(new_n1276), .C2(new_n1283), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n753), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1344), .B1(new_n1242), .B2(new_n1269), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1345), .B1(new_n1274), .B2(new_n1308), .ZN(new_n1346));
  AND3_X1   g1146(.A1(new_n1310), .A2(new_n1313), .A3(new_n1346), .ZN(new_n1347));
  OAI21_X1  g1147(.A(KEYINPUT124), .B1(new_n1343), .B2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1276), .A2(new_n1283), .ZN(new_n1349));
  INV_X1    g1149(.A(new_n1272), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1349), .A2(G378), .A3(new_n1350), .ZN(new_n1351));
  INV_X1    g1151(.A(KEYINPUT124), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1310), .A2(new_n1313), .A3(new_n1346), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1351), .A2(new_n1352), .A3(new_n1353), .ZN(new_n1354));
  INV_X1    g1154(.A(KEYINPUT60), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1306), .A2(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1356), .A2(new_n701), .ZN(new_n1357));
  AOI21_X1  g1157(.A(new_n1357), .B1(new_n1307), .B2(KEYINPUT60), .ZN(new_n1358));
  INV_X1    g1158(.A(new_n1358), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1359), .A2(G384), .A3(new_n1305), .ZN(new_n1360));
  INV_X1    g1160(.A(new_n1305), .ZN(new_n1361));
  OAI211_X1 g1161(.A(new_n826), .B(new_n850), .C1(new_n1358), .C2(new_n1361), .ZN(new_n1362));
  AND2_X1   g1162(.A1(new_n1360), .A2(new_n1362), .ZN(new_n1363));
  NAND4_X1  g1163(.A1(new_n1348), .A2(new_n1319), .A3(new_n1354), .A4(new_n1363), .ZN(new_n1364));
  INV_X1    g1164(.A(KEYINPUT62), .ZN(new_n1365));
  AOI21_X1  g1165(.A(new_n1320), .B1(new_n1351), .B2(new_n1353), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1360), .A2(new_n1362), .ZN(new_n1367));
  NOR2_X1   g1167(.A1(new_n1367), .A2(new_n1365), .ZN(new_n1368));
  AOI22_X1  g1168(.A1(new_n1364), .A2(new_n1365), .B1(new_n1366), .B2(new_n1368), .ZN(new_n1369));
  INV_X1    g1169(.A(KEYINPUT61), .ZN(new_n1370));
  AOI21_X1  g1170(.A(new_n1363), .B1(G2897), .B2(new_n1320), .ZN(new_n1371));
  INV_X1    g1171(.A(G2897), .ZN(new_n1372));
  NOR3_X1   g1172(.A1(new_n1367), .A2(new_n1372), .A3(new_n1319), .ZN(new_n1373));
  NOR2_X1   g1173(.A1(new_n1371), .A2(new_n1373), .ZN(new_n1374));
  OAI21_X1  g1174(.A(new_n1370), .B1(new_n1374), .B2(new_n1366), .ZN(new_n1375));
  OAI21_X1  g1175(.A(new_n1342), .B1(new_n1369), .B2(new_n1375), .ZN(new_n1376));
  INV_X1    g1176(.A(KEYINPUT63), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(new_n1364), .A2(new_n1377), .ZN(new_n1378));
  NAND3_X1  g1178(.A1(new_n1348), .A2(new_n1319), .A3(new_n1354), .ZN(new_n1379));
  OR2_X1    g1179(.A1(new_n1371), .A2(new_n1373), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1379), .A2(new_n1380), .ZN(new_n1381));
  INV_X1    g1181(.A(new_n1320), .ZN(new_n1382));
  NOR2_X1   g1182(.A1(new_n1367), .A2(new_n1377), .ZN(new_n1383));
  OAI211_X1 g1183(.A(new_n1382), .B(new_n1383), .C1(new_n1343), .C2(new_n1347), .ZN(new_n1384));
  AOI21_X1  g1184(.A(KEYINPUT61), .B1(new_n1335), .B2(new_n1340), .ZN(new_n1385));
  NAND2_X1  g1185(.A1(new_n1384), .A2(new_n1385), .ZN(new_n1386));
  INV_X1    g1186(.A(new_n1386), .ZN(new_n1387));
  AND4_X1   g1187(.A1(KEYINPUT127), .A2(new_n1378), .A3(new_n1381), .A4(new_n1387), .ZN(new_n1388));
  AOI21_X1  g1188(.A(new_n1386), .B1(new_n1379), .B2(new_n1380), .ZN(new_n1389));
  AOI21_X1  g1189(.A(KEYINPUT127), .B1(new_n1389), .B2(new_n1378), .ZN(new_n1390));
  OAI21_X1  g1190(.A(new_n1376), .B1(new_n1388), .B2(new_n1390), .ZN(G405));
  NOR2_X1   g1191(.A1(new_n1284), .A2(new_n1314), .ZN(new_n1392));
  NOR2_X1   g1192(.A1(new_n1392), .A2(new_n1343), .ZN(new_n1393));
  XNOR2_X1  g1193(.A(new_n1393), .B(new_n1367), .ZN(new_n1394));
  XNOR2_X1  g1194(.A(new_n1394), .B(new_n1342), .ZN(G402));
endmodule


