//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 1 1 0 0 0 1 0 0 1 1 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n878, new_n879, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948;
  INV_X1    g000(.A(G478), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(KEYINPUT15), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G122), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G116), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT14), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n193), .B(KEYINPUT97), .ZN(new_n194));
  INV_X1    g008(.A(G116), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G122), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n197), .B1(new_n192), .B2(KEYINPUT14), .ZN(new_n198));
  OAI21_X1  g012(.A(G107), .B1(new_n194), .B2(new_n198), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n196), .A2(new_n191), .ZN(new_n200));
  INV_X1    g014(.A(G107), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT66), .ZN(new_n203));
  INV_X1    g017(.A(G134), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(KEYINPUT66), .A2(G134), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT94), .ZN(new_n208));
  AND2_X1   g022(.A1(KEYINPUT68), .A2(G128), .ZN(new_n209));
  NOR2_X1   g023(.A1(KEYINPUT68), .A2(G128), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n208), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT68), .B(G128), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(KEYINPUT94), .A3(G143), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G128), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(G143), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n207), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  AND2_X1   g034(.A1(KEYINPUT66), .A2(G134), .ZN(new_n221));
  NOR2_X1   g035(.A1(KEYINPUT66), .A2(G134), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI211_X1 g037(.A(new_n223), .B(new_n218), .C1(new_n213), .C2(new_n215), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n199), .B(new_n202), .C1(new_n220), .C2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(KEYINPUT96), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n216), .A2(new_n207), .A3(new_n219), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT96), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(new_n200), .B(new_n201), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n226), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT95), .ZN(new_n232));
  INV_X1    g046(.A(new_n216), .ZN(new_n233));
  XNOR2_X1  g047(.A(new_n218), .B(KEYINPUT13), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n232), .B(G134), .C1(new_n233), .C2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n234), .B1(new_n213), .B2(new_n215), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT95), .B1(new_n236), .B2(new_n204), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n225), .B1(new_n231), .B2(new_n238), .ZN(new_n239));
  XOR2_X1   g053(.A(KEYINPUT9), .B(G234), .Z(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G217), .ZN(new_n242));
  NOR3_X1   g056(.A1(new_n241), .A2(new_n242), .A3(G953), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n239), .A2(new_n244), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n225), .B(new_n243), .C1(new_n231), .C2(new_n238), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G902), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n189), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  AOI211_X1 g063(.A(G902), .B(new_n188), .C1(new_n245), .C2(new_n246), .ZN(new_n250));
  OR2_X1    g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G125), .ZN(new_n253));
  NOR3_X1   g067(.A1(new_n253), .A2(KEYINPUT16), .A3(G140), .ZN(new_n254));
  NAND2_X1  g068(.A1(KEYINPUT76), .A2(G125), .ZN(new_n255));
  INV_X1    g069(.A(G140), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(KEYINPUT76), .A2(G125), .A3(G140), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n254), .B1(new_n259), .B2(KEYINPUT16), .ZN(new_n260));
  INV_X1    g074(.A(G146), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n260), .B(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G237), .ZN(new_n263));
  INV_X1    g077(.A(G953), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n264), .A3(G214), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(KEYINPUT91), .A3(new_n212), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n212), .A2(KEYINPUT91), .ZN(new_n267));
  NOR2_X1   g081(.A1(G237), .A2(G953), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n267), .A2(G214), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(KEYINPUT17), .A3(G131), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n270), .B(G131), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n262), .B(new_n271), .C1(new_n272), .C2(KEYINPUT17), .ZN(new_n273));
  XNOR2_X1  g087(.A(G113), .B(G122), .ZN(new_n274));
  INV_X1    g088(.A(G104), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n274), .B(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n257), .A2(G146), .A3(new_n258), .ZN(new_n277));
  OR2_X1    g091(.A1(new_n277), .A2(KEYINPUT92), .ZN(new_n278));
  XNOR2_X1  g092(.A(G125), .B(G140), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n261), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n280), .A2(KEYINPUT92), .A3(new_n277), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT18), .ZN(new_n282));
  INV_X1    g096(.A(G131), .ZN(new_n283));
  NOR3_X1   g097(.A1(new_n270), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n266), .A2(new_n269), .B1(KEYINPUT18), .B2(G131), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n278), .B(new_n281), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  AND3_X1   g100(.A1(new_n273), .A2(new_n276), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n276), .B1(new_n273), .B2(new_n286), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n248), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT93), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI211_X1 g105(.A(KEYINPUT93), .B(new_n248), .C1(new_n287), .C2(new_n288), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n291), .A2(G475), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n260), .A2(G146), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n259), .A2(KEYINPUT19), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n279), .A2(KEYINPUT19), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n261), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n272), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n286), .ZN(new_n299));
  INV_X1    g113(.A(new_n276), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n273), .A2(new_n276), .A3(new_n286), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G475), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n304), .A3(new_n248), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT20), .ZN(new_n306));
  OR2_X1    g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n306), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n293), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n252), .A2(new_n309), .ZN(new_n310));
  AND2_X1   g124(.A1(new_n264), .A2(G952), .ZN(new_n311));
  NAND2_X1  g125(.A1(G234), .A2(G237), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  XOR2_X1   g128(.A(KEYINPUT21), .B(G898), .Z(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n312), .A2(G902), .A3(G953), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n314), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n310), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(G221), .B1(new_n241), .B2(G902), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n201), .A2(G104), .ZN(new_n322));
  AND2_X1   g136(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n323));
  NOR2_X1   g137(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n275), .A2(G107), .ZN(new_n326));
  NAND2_X1  g140(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT80), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n329), .B1(new_n201), .B2(G104), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n275), .A2(KEYINPUT80), .A3(G107), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n325), .A2(new_n328), .A3(new_n330), .A4(new_n331), .ZN(new_n332));
  OR2_X1    g146(.A1(new_n332), .A2(G101), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n261), .A2(G143), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n212), .A2(G146), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(new_n335), .A3(G128), .ZN(new_n336));
  OR2_X1    g150(.A1(new_n336), .A2(KEYINPUT1), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n334), .A2(new_n335), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n217), .B1(new_n334), .B2(KEYINPUT1), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n201), .A2(G104), .ZN(new_n341));
  OAI21_X1  g155(.A(G101), .B1(new_n326), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n333), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n342), .B1(new_n332), .B2(G101), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n334), .A2(KEYINPUT1), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n211), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT65), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n348), .B1(new_n261), .B2(G143), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n212), .A2(KEYINPUT65), .A3(G146), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n351), .A2(new_n334), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n337), .B1(new_n347), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n343), .B1(new_n345), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(G137), .B1(new_n221), .B2(new_n222), .ZN(new_n355));
  XNOR2_X1  g169(.A(KEYINPUT67), .B(G137), .ZN(new_n356));
  NAND2_X1  g170(.A1(KEYINPUT11), .A2(G134), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G137), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT11), .B1(new_n223), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(G131), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT11), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n362), .B1(new_n207), .B2(G137), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n359), .A2(KEYINPUT67), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT67), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G137), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n357), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n363), .A2(new_n368), .A3(new_n283), .A4(new_n355), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n361), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(KEYINPUT12), .B1(new_n354), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n354), .A2(KEYINPUT12), .A3(new_n370), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n332), .A2(G101), .ZN(new_n375));
  NAND2_X1  g189(.A1(KEYINPUT81), .A2(KEYINPUT4), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n376), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n332), .A2(G101), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(new_n333), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT0), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n336), .A2(new_n381), .ZN(new_n382));
  AOI22_X1  g196(.A1(new_n351), .A2(new_n334), .B1(new_n381), .B2(new_n217), .ZN(new_n383));
  NAND2_X1  g197(.A1(KEYINPUT0), .A2(G128), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(KEYINPUT64), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n382), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n380), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT10), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n343), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n370), .ZN(new_n390));
  AOI22_X1  g204(.A1(new_n351), .A2(new_n334), .B1(new_n211), .B2(new_n346), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n336), .A2(KEYINPUT1), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT10), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n393), .A2(new_n344), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n387), .A2(new_n389), .A3(new_n390), .A4(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT85), .ZN(new_n397));
  XNOR2_X1  g211(.A(G110), .B(G140), .ZN(new_n398));
  INV_X1    g212(.A(G227), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n399), .A2(G953), .ZN(new_n400));
  XOR2_X1   g214(.A(new_n398), .B(new_n400), .Z(new_n401));
  AND3_X1   g215(.A1(new_n396), .A2(new_n397), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n397), .B1(new_n396), .B2(new_n401), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n374), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT86), .ZN(new_n405));
  INV_X1    g219(.A(new_n401), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT83), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n394), .B1(new_n380), .B2(new_n386), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n407), .B1(new_n408), .B2(new_n389), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(new_n407), .A3(new_n389), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n390), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n396), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n406), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT86), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n374), .B(new_n415), .C1(new_n402), .C2(new_n403), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n405), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G469), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n417), .A2(new_n418), .A3(new_n248), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n408), .A2(new_n407), .A3(new_n389), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n370), .B1(new_n420), .B2(new_n409), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n396), .A2(new_n401), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT82), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n396), .A2(KEYINPUT82), .A3(new_n401), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n421), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n373), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n396), .B1(new_n427), .B2(new_n371), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n406), .ZN(new_n429));
  AND3_X1   g243(.A1(new_n426), .A2(new_n429), .A3(KEYINPUT84), .ZN(new_n430));
  AOI21_X1  g244(.A(KEYINPUT84), .B1(new_n426), .B2(new_n429), .ZN(new_n431));
  OAI21_X1  g245(.A(G469), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n418), .A2(new_n248), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n419), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n320), .A2(new_n321), .A3(new_n435), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n217), .A2(G119), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n437), .B1(new_n214), .B2(G119), .ZN(new_n438));
  XOR2_X1   g252(.A(KEYINPUT24), .B(G110), .Z(new_n439));
  AOI21_X1  g253(.A(new_n262), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(KEYINPUT23), .B1(new_n217), .B2(G119), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT23), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n442), .B1(new_n438), .B2(new_n443), .ZN(new_n444));
  OR2_X1    g258(.A1(new_n444), .A2(KEYINPUT75), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(KEYINPUT75), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(G110), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n440), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n438), .A2(new_n439), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT77), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n449), .B(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n444), .A2(G110), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n294), .B(new_n280), .C1(new_n451), .C2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n448), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n264), .A2(G221), .A3(G234), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(KEYINPUT22), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n456), .B(G137), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n448), .A2(new_n453), .A3(new_n457), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n248), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT25), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n242), .B1(G234), .B2(new_n248), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT25), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n459), .A2(new_n464), .A3(new_n248), .A4(new_n460), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n462), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n459), .A2(new_n460), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n463), .A2(G902), .ZN(new_n468));
  XOR2_X1   g282(.A(new_n468), .B(KEYINPUT78), .Z(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n332), .A2(G101), .A3(new_n378), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n378), .B1(new_n332), .B2(G101), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n332), .A2(G101), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(KEYINPUT2), .A2(G113), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT69), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT69), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n479), .B1(KEYINPUT2), .B2(G113), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n478), .A2(new_n480), .B1(KEYINPUT2), .B2(G113), .ZN(new_n481));
  XNOR2_X1  g295(.A(G116), .B(G119), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT70), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n481), .A2(KEYINPUT70), .A3(new_n482), .ZN(new_n486));
  INV_X1    g300(.A(new_n481), .ZN(new_n487));
  INV_X1    g301(.A(new_n482), .ZN(new_n488));
  AOI22_X1  g302(.A1(new_n485), .A2(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(KEYINPUT87), .B1(new_n476), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n485), .A2(new_n486), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n482), .A2(KEYINPUT5), .ZN(new_n492));
  OR2_X1    g306(.A1(new_n195), .A2(G119), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n492), .B(G113), .C1(KEYINPUT5), .C2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n491), .A2(new_n345), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n487), .A2(new_n488), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT87), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n497), .A2(new_n380), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n490), .A2(new_n495), .A3(new_n499), .ZN(new_n500));
  XOR2_X1   g314(.A(G110), .B(G122), .Z(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n501), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n490), .A2(new_n503), .A3(new_n499), .A4(new_n495), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n502), .A2(KEYINPUT6), .A3(new_n504), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n337), .B(new_n253), .C1(new_n352), .C2(new_n347), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n506), .B1(new_n386), .B2(new_n253), .ZN(new_n507));
  INV_X1    g321(.A(G224), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n508), .A2(G953), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n507), .B(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT6), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n500), .A2(new_n511), .A3(new_n501), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n505), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  XOR2_X1   g327(.A(new_n501), .B(KEYINPUT8), .Z(new_n514));
  INV_X1    g328(.A(new_n495), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n345), .B1(new_n491), .B2(new_n494), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT88), .ZN(new_n518));
  OR2_X1    g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n507), .B1(KEYINPUT89), .B2(KEYINPUT7), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT7), .B1(new_n508), .B2(G953), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n520), .B(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n517), .A2(new_n518), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n519), .A2(new_n522), .A3(new_n504), .A4(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n513), .A2(new_n248), .A3(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(G210), .B1(G237), .B2(G902), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT90), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n513), .A2(new_n248), .A3(new_n526), .A4(new_n524), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n525), .A2(KEYINPUT90), .A3(new_n527), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(G214), .B1(G237), .B2(G902), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(G472), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n356), .A2(new_n204), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n207), .A2(G137), .ZN(new_n539));
  OAI21_X1  g353(.A(G131), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n353), .A2(new_n540), .A3(new_n369), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT71), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n370), .A2(new_n542), .A3(new_n386), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n542), .B1(new_n370), .B2(new_n386), .ZN(new_n544));
  OAI211_X1 g358(.A(KEYINPUT30), .B(new_n541), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n358), .A2(new_n360), .A3(G131), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n359), .B1(new_n205), .B2(new_n206), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n367), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n283), .B1(new_n548), .B2(new_n363), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n386), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n541), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT30), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT72), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n545), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n550), .A2(KEYINPUT71), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n370), .A2(new_n542), .A3(new_n386), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n557), .A2(KEYINPUT72), .A3(KEYINPUT30), .A4(new_n541), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n497), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n557), .A2(new_n489), .A3(new_n541), .ZN(new_n561));
  XOR2_X1   g375(.A(KEYINPUT73), .B(KEYINPUT27), .Z(new_n562));
  NAND2_X1  g376(.A1(new_n268), .A2(G210), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n562), .B(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(KEYINPUT26), .B(G101), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n564), .B(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  XOR2_X1   g381(.A(KEYINPUT74), .B(KEYINPUT31), .Z(new_n568));
  NAND4_X1  g382(.A1(new_n560), .A2(new_n561), .A3(new_n567), .A4(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n551), .A2(new_n497), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT28), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n571), .B1(new_n551), .B2(new_n497), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n570), .B(new_n572), .C1(new_n561), .C2(new_n571), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n566), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT31), .ZN(new_n576));
  INV_X1    g390(.A(new_n561), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n577), .B1(new_n559), .B2(new_n497), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n576), .B1(new_n578), .B2(new_n567), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n537), .B(new_n248), .C1(new_n575), .C2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT32), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI211_X1 g396(.A(new_n566), .B(new_n577), .C1(new_n559), .C2(new_n497), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n569), .B(new_n574), .C1(new_n583), .C2(new_n576), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n584), .A2(KEYINPUT32), .A3(new_n537), .A4(new_n248), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n578), .A2(new_n566), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n573), .A2(new_n567), .ZN(new_n587));
  AOI21_X1  g401(.A(KEYINPUT29), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n541), .B1(new_n543), .B2(new_n544), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n497), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(new_n561), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT28), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n592), .A2(KEYINPUT29), .A3(new_n567), .A4(new_n572), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n248), .ZN(new_n594));
  OAI21_X1  g408(.A(G472), .B1(new_n588), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n582), .A2(new_n585), .A3(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n436), .A2(new_n472), .A3(new_n536), .A4(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(G101), .ZN(G3));
  OAI21_X1  g412(.A(new_n248), .B1(new_n575), .B2(new_n579), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n537), .A2(KEYINPUT98), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n435), .A2(new_n472), .A3(new_n321), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n535), .B1(new_n528), .B2(new_n530), .ZN(new_n604));
  INV_X1    g418(.A(new_n319), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n293), .A2(new_n307), .A3(new_n308), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n247), .A2(new_n187), .A3(new_n248), .ZN(new_n607));
  XOR2_X1   g421(.A(KEYINPUT99), .B(KEYINPUT33), .Z(new_n608));
  AND3_X1   g422(.A1(new_n245), .A2(new_n246), .A3(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT99), .ZN(new_n610));
  AOI22_X1  g424(.A1(new_n245), .A2(new_n246), .B1(new_n610), .B2(KEYINPUT33), .ZN(new_n611));
  OAI21_X1  g425(.A(G478), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(G478), .A2(G902), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n606), .A2(new_n607), .A3(new_n612), .A4(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n604), .A2(new_n605), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n603), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT34), .B(G104), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G6));
  NAND2_X1  g433(.A1(new_n309), .A2(new_n251), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n604), .A2(new_n605), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n603), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT35), .B(G107), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT100), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n623), .B(new_n625), .ZN(G9));
  INV_X1    g440(.A(new_n601), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT101), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n458), .A2(KEYINPUT36), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n454), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n469), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n466), .A2(new_n628), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n628), .B1(new_n466), .B2(new_n631), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n627), .A2(new_n436), .A3(new_n536), .A4(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(new_n635), .B(KEYINPUT37), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G110), .ZN(G12));
  OR3_X1    g451(.A1(new_n317), .A2(KEYINPUT102), .A3(G900), .ZN(new_n638));
  OAI21_X1  g452(.A(KEYINPUT102), .B1(new_n317), .B2(G900), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n638), .A2(new_n313), .A3(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n620), .A2(new_n641), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n435), .A2(new_n642), .A3(new_n321), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n643), .A2(new_n596), .A3(new_n604), .A4(new_n634), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT103), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(new_n217), .ZN(G30));
  AND2_X1   g460(.A1(new_n435), .A2(new_n321), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n640), .B(KEYINPUT39), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT40), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n251), .A2(new_n606), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n533), .B(KEYINPUT38), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n578), .A2(new_n566), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n248), .B1(new_n591), .B2(new_n567), .ZN(new_n657));
  OAI21_X1  g471(.A(G472), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n582), .A2(new_n585), .A3(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n660), .A2(new_n535), .A3(new_n634), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n651), .A2(new_n653), .A3(new_n655), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT104), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(new_n212), .ZN(G45));
  AND2_X1   g478(.A1(new_n596), .A2(new_n634), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n614), .A2(new_n641), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n665), .A2(new_n647), .A3(new_n604), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G146), .ZN(G48));
  NAND2_X1  g482(.A1(KEYINPUT105), .A2(G469), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n417), .A2(new_n248), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n669), .B1(new_n417), .B2(new_n248), .ZN(new_n671));
  INV_X1    g485(.A(new_n321), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n596), .A2(new_n616), .A3(new_n472), .A4(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT41), .B(G113), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G15));
  NAND4_X1  g490(.A1(new_n596), .A2(new_n622), .A3(new_n472), .A4(new_n673), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G116), .ZN(G18));
  NAND4_X1  g492(.A1(new_n596), .A2(new_n320), .A3(new_n604), .A4(new_n634), .ZN(new_n679));
  INV_X1    g493(.A(new_n673), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(new_n681), .B(G119), .Z(G21));
  XNOR2_X1  g496(.A(new_n471), .B(KEYINPUT107), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n599), .A2(G472), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n592), .A2(new_n685), .A3(new_n572), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n571), .B1(new_n590), .B2(new_n561), .ZN(new_n687));
  INV_X1    g501(.A(new_n572), .ZN(new_n688));
  OAI21_X1  g502(.A(KEYINPUT106), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n686), .A2(new_n566), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n569), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n537), .B(new_n248), .C1(new_n691), .C2(new_n579), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n683), .A2(new_n684), .A3(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n604), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n695), .A2(new_n319), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n694), .A2(new_n696), .A3(new_n653), .A4(new_n673), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT108), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n680), .A2(new_n693), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n700), .A2(KEYINPUT108), .A3(new_n696), .A4(new_n653), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G122), .ZN(G24));
  AND3_X1   g517(.A1(new_n692), .A2(new_n684), .A3(new_n634), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n704), .A2(new_n604), .A3(new_n666), .A4(new_n673), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G125), .ZN(G27));
  NAND2_X1  g520(.A1(new_n596), .A2(new_n683), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n672), .A2(new_n535), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n709), .B1(new_n531), .B2(new_n532), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n426), .A2(new_n429), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(G469), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n419), .A2(new_n434), .A3(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n710), .A2(new_n666), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g528(.A(KEYINPUT42), .B1(new_n707), .B2(new_n714), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n710), .A2(new_n713), .ZN(new_n716));
  INV_X1    g530(.A(new_n666), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n717), .A2(KEYINPUT42), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n716), .A2(new_n472), .A3(new_n596), .A4(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(new_n283), .ZN(G33));
  NAND4_X1  g535(.A1(new_n596), .A2(new_n472), .A3(new_n713), .A4(new_n710), .ZN(new_n722));
  INV_X1    g536(.A(new_n642), .ZN(new_n723));
  OR2_X1    g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT109), .B(G134), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G36));
  AOI21_X1  g540(.A(new_n535), .B1(new_n531), .B2(new_n532), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n601), .A2(new_n634), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT112), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n612), .A2(new_n607), .A3(new_n613), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n606), .B1(new_n732), .B2(KEYINPUT111), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT111), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n734), .A2(KEYINPUT43), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n733), .B1(new_n732), .B2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT110), .ZN(new_n737));
  OR2_X1    g551(.A1(new_n737), .A2(KEYINPUT43), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  OR2_X1    g553(.A1(new_n732), .A2(new_n606), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n737), .A3(KEYINPUT43), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n731), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n728), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n711), .A2(KEYINPUT45), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n430), .A2(new_n431), .ZN(new_n746));
  OAI211_X1 g560(.A(G469), .B(new_n745), .C1(new_n746), .C2(KEYINPUT45), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n434), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT46), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n747), .A2(KEYINPUT46), .A3(new_n434), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(new_n419), .A3(new_n751), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n752), .A2(new_n321), .A3(new_n648), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n731), .A2(KEYINPUT44), .A3(new_n739), .A4(new_n741), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n744), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G137), .ZN(G39));
  NAND2_X1  g570(.A1(new_n752), .A2(new_n321), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT47), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n752), .A2(KEYINPUT47), .A3(new_n321), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n728), .A2(new_n596), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n761), .A2(new_n471), .A3(new_n666), .A4(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G140), .ZN(G42));
  NOR2_X1   g578(.A1(new_n670), .A2(new_n671), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT49), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n683), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n767), .A2(new_n709), .A3(new_n740), .ZN(new_n768));
  XOR2_X1   g582(.A(new_n768), .B(KEYINPUT113), .Z(new_n769));
  AOI21_X1  g583(.A(new_n659), .B1(new_n766), .B2(new_n765), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(new_n654), .A3(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT50), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n741), .A2(new_n736), .A3(new_n314), .A4(new_n738), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n774), .A2(new_n673), .A3(new_n694), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n654), .A2(new_n535), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n772), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n773), .A2(new_n680), .A3(new_n693), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n778), .A2(KEYINPUT50), .A3(new_n535), .A4(new_n654), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT118), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n777), .A2(KEYINPUT118), .A3(new_n779), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n710), .A2(new_n765), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n773), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT119), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n704), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n660), .A2(new_n314), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n710), .A2(new_n472), .A3(new_n765), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(new_n309), .A3(new_n732), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n773), .A2(new_n693), .A3(new_n728), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n765), .A2(new_n672), .ZN(new_n795));
  XOR2_X1   g609(.A(new_n795), .B(KEYINPUT117), .Z(new_n796));
  OAI21_X1  g610(.A(new_n794), .B1(new_n761), .B2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n784), .A2(new_n789), .A3(new_n793), .A4(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT51), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n789), .A2(new_n780), .A3(new_n793), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n759), .A2(new_n760), .A3(new_n795), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n799), .B1(new_n802), .B2(new_n794), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n801), .A2(new_n803), .A3(KEYINPUT120), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT120), .B1(new_n801), .B2(new_n803), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n800), .B(new_n311), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n647), .A2(new_n596), .A3(new_n604), .A4(new_n634), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n705), .B(new_n644), .C1(new_n809), .C2(new_n717), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n695), .A2(new_n641), .A3(new_n652), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n713), .A2(new_n466), .A3(new_n631), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n811), .A2(new_n812), .A3(new_n321), .A4(new_n659), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n808), .B1(new_n810), .B2(new_n814), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n705), .A2(new_n644), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n816), .A2(KEYINPUT52), .A3(new_n667), .A4(new_n813), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(KEYINPUT114), .B1(new_n310), .B2(new_n641), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n596), .A2(new_n634), .A3(new_n819), .ZN(new_n820));
  OR4_X1    g634(.A1(KEYINPUT114), .A2(new_n251), .A3(new_n606), .A4(new_n641), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n727), .A2(new_n821), .A3(new_n321), .A4(new_n435), .ZN(new_n822));
  OAI22_X1  g636(.A1(new_n722), .A2(new_n723), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n716), .A2(new_n666), .A3(new_n704), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n720), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n674), .B(new_n677), .C1(new_n679), .C2(new_n680), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n826), .B1(new_n699), .B2(new_n701), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n620), .A2(new_n614), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n603), .A2(new_n536), .A3(new_n605), .A4(new_n828), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n829), .A2(new_n597), .A3(new_n635), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n825), .A2(new_n827), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n832));
  OR3_X1    g646(.A1(new_n818), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n825), .A2(new_n830), .A3(new_n827), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n815), .A2(new_n817), .A3(KEYINPUT115), .ZN(new_n835));
  OR2_X1    g649(.A1(new_n817), .A2(KEYINPUT115), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n833), .B1(new_n837), .B2(KEYINPUT53), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT54), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n774), .A2(new_n604), .A3(new_n673), .A4(new_n694), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n832), .B1(new_n818), .B2(new_n831), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n834), .A2(new_n836), .A3(KEYINPUT53), .A4(new_n835), .ZN(new_n845));
  OAI211_X1 g659(.A(KEYINPUT116), .B(new_n832), .C1(new_n818), .C2(new_n831), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n843), .A2(new_n844), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n807), .A2(new_n839), .A3(new_n840), .A4(new_n847), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n790), .A2(new_n614), .A3(new_n791), .ZN(new_n849));
  INV_X1    g663(.A(new_n707), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n788), .A2(new_n850), .ZN(new_n851));
  XOR2_X1   g665(.A(new_n851), .B(KEYINPUT48), .Z(new_n852));
  NOR3_X1   g666(.A1(new_n848), .A2(new_n849), .A3(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(G952), .A2(G953), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n771), .B1(new_n853), .B2(new_n854), .ZN(G75));
  NAND3_X1  g669(.A1(new_n843), .A2(new_n845), .A3(new_n846), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n856), .A2(G902), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(G210), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT56), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n505), .A2(new_n512), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(new_n510), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(KEYINPUT55), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n858), .A2(new_n859), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n862), .B1(new_n858), .B2(new_n859), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n264), .A2(G952), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(G51));
  INV_X1    g680(.A(KEYINPUT121), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n856), .A2(KEYINPUT54), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(new_n847), .ZN(new_n869));
  XOR2_X1   g683(.A(new_n433), .B(KEYINPUT57), .Z(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n867), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  AOI211_X1 g686(.A(KEYINPUT121), .B(new_n870), .C1(new_n868), .C2(new_n847), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n417), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n747), .B(KEYINPUT122), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n857), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n865), .B1(new_n874), .B2(new_n876), .ZN(G54));
  NAND3_X1  g691(.A1(new_n857), .A2(KEYINPUT58), .A3(G475), .ZN(new_n878));
  INV_X1    g692(.A(new_n303), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n878), .A2(new_n879), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n880), .A2(new_n881), .A3(new_n865), .ZN(G60));
  OR2_X1    g696(.A1(new_n609), .A2(new_n611), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n613), .B(KEYINPUT59), .Z(new_n884));
  NOR2_X1   g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n886), .B1(new_n868), .B2(new_n847), .ZN(new_n887));
  OR3_X1    g701(.A1(new_n887), .A2(KEYINPUT123), .A3(new_n865), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n839), .A2(new_n847), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n883), .B1(new_n889), .B2(new_n884), .ZN(new_n890));
  OAI21_X1  g704(.A(KEYINPUT123), .B1(new_n887), .B2(new_n865), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n888), .A2(new_n890), .A3(new_n891), .ZN(G63));
  NAND2_X1  g706(.A1(G217), .A2(G902), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT60), .Z(new_n894));
  NAND3_X1  g708(.A1(new_n856), .A2(new_n630), .A3(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n865), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n856), .A2(new_n894), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n895), .B(new_n896), .C1(new_n467), .C2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT61), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n898), .B(new_n899), .ZN(G66));
  OAI21_X1  g714(.A(G953), .B1(new_n316), .B2(new_n508), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n827), .A2(new_n830), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n901), .B1(new_n902), .B2(G953), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n860), .B1(G898), .B2(new_n264), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n903), .B(new_n904), .ZN(G69));
  NOR2_X1   g719(.A1(new_n295), .A2(new_n296), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n559), .B(new_n906), .Z(new_n907));
  AND2_X1   g721(.A1(new_n755), .A2(new_n763), .ZN(new_n908));
  INV_X1    g722(.A(new_n810), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n662), .A2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT62), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n910), .B(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n649), .A2(new_n728), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n913), .A2(new_n472), .A3(new_n596), .A4(new_n828), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n908), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n907), .B1(new_n915), .B2(new_n264), .ZN(new_n916));
  INV_X1    g730(.A(G900), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n907), .B1(new_n917), .B2(new_n264), .ZN(new_n918));
  INV_X1    g732(.A(new_n720), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n695), .A2(new_n652), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n753), .A2(KEYINPUT124), .A3(new_n850), .A4(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT124), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n752), .A2(new_n321), .A3(new_n648), .A4(new_n920), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n922), .B1(new_n923), .B2(new_n707), .ZN(new_n924));
  AND4_X1   g738(.A1(new_n724), .A2(new_n921), .A3(new_n909), .A4(new_n924), .ZN(new_n925));
  AND4_X1   g739(.A1(new_n919), .A2(new_n925), .A3(new_n755), .A4(new_n763), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n918), .B1(new_n926), .B2(new_n264), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n916), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(G953), .B1(new_n399), .B2(new_n917), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n928), .B(new_n929), .ZN(G72));
  INV_X1    g744(.A(new_n656), .ZN(new_n931));
  NAND2_X1  g745(.A1(G472), .A2(G902), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT63), .Z(new_n933));
  NAND4_X1  g747(.A1(new_n838), .A2(new_n586), .A3(new_n931), .A4(new_n933), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT127), .Z(new_n935));
  NAND4_X1  g749(.A1(new_n908), .A2(new_n902), .A3(new_n912), .A4(new_n914), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n931), .B1(new_n936), .B2(new_n933), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT125), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n908), .A2(new_n925), .A3(new_n919), .A4(new_n902), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n586), .B1(new_n940), .B2(new_n933), .ZN(new_n941));
  OAI21_X1  g755(.A(KEYINPUT126), .B1(new_n941), .B2(new_n865), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT126), .ZN(new_n943));
  INV_X1    g757(.A(new_n933), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n926), .B2(new_n902), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n943), .B(new_n896), .C1(new_n945), .C2(new_n586), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n942), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n935), .A2(new_n939), .A3(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(G57));
endmodule


