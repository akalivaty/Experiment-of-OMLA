//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 0 0 0 1 0 0 1 1 1 1 0 1 0 1 1 0 1 0 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1 0 1 0 1 1 0 0 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996;
  INV_X1    g000(.A(KEYINPUT94), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT90), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT89), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  INV_X1    g004(.A(G237), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G214), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n189), .A2(G143), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n190), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT89), .ZN(new_n197));
  NOR2_X1   g011(.A1(G237), .A2(G953), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n197), .B1(G214), .B2(new_n198), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n188), .B1(new_n195), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n193), .A2(new_n190), .ZN(new_n201));
  AOI22_X1  g015(.A1(new_n198), .A2(G214), .B1(new_n189), .B2(G143), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n201), .B(KEYINPUT90), .C1(new_n202), .C2(new_n190), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n200), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(KEYINPUT18), .A2(G131), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  AOI21_X1  g020(.A(KEYINPUT91), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT91), .ZN(new_n208));
  AOI211_X1 g022(.A(new_n208), .B(new_n205), .C1(new_n200), .C2(new_n203), .ZN(new_n209));
  INV_X1    g023(.A(G214), .ZN(new_n210));
  NOR3_X1   g024(.A1(new_n210), .A2(G237), .A3(G953), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n196), .A2(KEYINPUT89), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n197), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(new_n205), .A3(new_n201), .ZN(new_n214));
  XNOR2_X1  g028(.A(G125), .B(G140), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G140), .ZN(new_n218));
  INV_X1    g032(.A(G125), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n218), .B1(new_n219), .B2(KEYINPUT78), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT78), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(G125), .A3(G140), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n220), .A2(G146), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n217), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n214), .A2(new_n224), .ZN(new_n225));
  NOR3_X1   g039(.A1(new_n207), .A2(new_n209), .A3(new_n225), .ZN(new_n226));
  OR2_X1    g040(.A1(new_n215), .A2(KEYINPUT19), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n220), .A2(new_n222), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT19), .ZN(new_n229));
  AOI21_X1  g043(.A(G146), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT16), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n231), .B1(new_n220), .B2(new_n222), .ZN(new_n232));
  NOR3_X1   g046(.A1(new_n219), .A2(KEYINPUT16), .A3(G140), .ZN(new_n233));
  NOR3_X1   g047(.A1(new_n232), .A2(new_n216), .A3(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(KEYINPUT93), .B1(new_n230), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n234), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT93), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n215), .A2(KEYINPUT19), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT19), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n239), .B1(new_n220), .B2(new_n222), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n216), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n236), .A2(new_n237), .A3(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n201), .B1(new_n202), .B2(new_n190), .ZN(new_n243));
  OAI21_X1  g057(.A(KEYINPUT92), .B1(new_n243), .B2(G131), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(G131), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT92), .ZN(new_n246));
  INV_X1    g060(.A(G131), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n213), .A2(new_n246), .A3(new_n247), .A4(new_n201), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n244), .A2(new_n245), .A3(new_n248), .ZN(new_n249));
  AND3_X1   g063(.A1(new_n235), .A2(new_n242), .A3(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n187), .B1(new_n226), .B2(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(G113), .B(G122), .ZN(new_n252));
  INV_X1    g066(.A(G104), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n252), .B(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n203), .ZN(new_n256));
  AOI21_X1  g070(.A(KEYINPUT90), .B1(new_n213), .B2(new_n201), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n206), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n208), .ZN(new_n259));
  INV_X1    g073(.A(new_n225), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n204), .A2(KEYINPUT91), .A3(new_n206), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n235), .A2(new_n242), .A3(new_n249), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(KEYINPUT94), .A3(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n251), .A2(new_n255), .A3(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n232), .A2(new_n233), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n266), .A2(G146), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n267), .A2(new_n234), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n243), .A2(KEYINPUT17), .A3(G131), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n268), .B(new_n269), .C1(new_n249), .C2(KEYINPUT17), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n262), .A2(new_n254), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n265), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G475), .ZN(new_n273));
  INV_X1    g087(.A(G902), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT20), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n271), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n254), .B1(new_n262), .B2(new_n270), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n274), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G475), .ZN(new_n281));
  AOI21_X1  g095(.A(G475), .B1(new_n265), .B2(new_n271), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(KEYINPUT20), .A3(new_n274), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n277), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G478), .ZN(new_n285));
  OR2_X1    g099(.A1(new_n285), .A2(KEYINPUT15), .ZN(new_n286));
  INV_X1    g100(.A(G116), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n287), .A2(G122), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n288), .B(KEYINPUT95), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(G122), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(KEYINPUT14), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n291), .A2(new_n292), .A3(G107), .ZN(new_n293));
  INV_X1    g107(.A(G128), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n294), .A2(G143), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(G143), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G134), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n298), .B(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G107), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n289), .B(new_n290), .C1(KEYINPUT14), .C2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n293), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n295), .A2(KEYINPUT96), .A3(KEYINPUT13), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n304), .B1(new_n295), .B2(KEYINPUT13), .ZN(new_n305));
  AOI22_X1  g119(.A1(KEYINPUT13), .A2(new_n295), .B1(new_n297), .B2(KEYINPUT96), .ZN(new_n306));
  OAI21_X1  g120(.A(G134), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n298), .A2(new_n299), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n289), .A2(new_n301), .A3(new_n290), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n301), .B1(new_n289), .B2(new_n290), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n307), .B(new_n308), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n303), .A2(new_n311), .ZN(new_n312));
  XOR2_X1   g126(.A(KEYINPUT9), .B(G234), .Z(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(G217), .A3(new_n192), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT97), .ZN(new_n316));
  INV_X1    g130(.A(new_n314), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n303), .A2(new_n311), .A3(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n315), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n303), .A2(new_n311), .A3(KEYINPUT97), .A4(new_n317), .ZN(new_n320));
  AND3_X1   g134(.A1(new_n319), .A2(new_n274), .A3(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n286), .B1(new_n321), .B2(KEYINPUT98), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n319), .A2(new_n320), .A3(new_n274), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n323), .B(KEYINPUT98), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n322), .B1(new_n324), .B2(new_n286), .ZN(new_n325));
  OR2_X1    g139(.A1(new_n284), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(G214), .B1(G237), .B2(G902), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(G143), .B(G146), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n294), .A2(KEYINPUT1), .ZN(new_n330));
  AOI21_X1  g144(.A(KEYINPUT69), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n216), .A2(G143), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n196), .A2(G146), .ZN(new_n333));
  AND4_X1   g147(.A1(KEYINPUT69), .A2(new_n330), .A3(new_n332), .A4(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n196), .A2(G146), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT65), .B1(new_n216), .B2(G143), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT65), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n337), .A2(new_n196), .A3(G146), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n335), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n294), .B1(new_n332), .B2(KEYINPUT1), .ZN(new_n340));
  OAI22_X1  g154(.A1(new_n331), .A2(new_n334), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n219), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT0), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n343), .A2(new_n294), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n345), .A2(new_n329), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n336), .A2(new_n338), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n332), .ZN(new_n348));
  NOR3_X1   g162(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n348), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n346), .B1(new_n352), .B2(new_n345), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n342), .B1(new_n353), .B2(new_n219), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT85), .B(G224), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT7), .B1(new_n355), .B2(G953), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n358), .B(KEYINPUT88), .ZN(new_n359));
  INV_X1    g173(.A(G119), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT70), .B1(new_n360), .B2(G116), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT70), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(new_n287), .A3(G119), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n360), .A2(G116), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(KEYINPUT5), .A3(new_n365), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n366), .B(G113), .C1(KEYINPUT5), .C2(new_n365), .ZN(new_n367));
  XOR2_X1   g181(.A(KEYINPUT2), .B(G113), .Z(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(new_n364), .A3(new_n365), .ZN(new_n369));
  OAI21_X1  g183(.A(KEYINPUT3), .B1(new_n253), .B2(G107), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT3), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n371), .A2(new_n301), .A3(G104), .ZN(new_n372));
  INV_X1    g186(.A(G101), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n253), .A2(G107), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n370), .A2(new_n372), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n301), .A2(G104), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n253), .A2(G107), .ZN(new_n377));
  OAI21_X1  g191(.A(G101), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n367), .A2(new_n369), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n364), .A2(new_n365), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n382), .B(new_n368), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n370), .A2(new_n372), .A3(new_n374), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G101), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(KEYINPUT4), .A3(new_n375), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT4), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n384), .A2(new_n387), .A3(G101), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n381), .B1(new_n383), .B2(new_n389), .ZN(new_n390));
  XOR2_X1   g204(.A(G110), .B(G122), .Z(new_n391));
  NOR2_X1   g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n354), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n392), .B1(new_n393), .B2(new_n356), .ZN(new_n394));
  XOR2_X1   g208(.A(KEYINPUT86), .B(KEYINPUT8), .Z(new_n395));
  XNOR2_X1  g209(.A(new_n391), .B(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n381), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n380), .B1(new_n367), .B2(new_n369), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT87), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OR2_X1    g215(.A1(new_n399), .A2(new_n400), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n359), .A2(new_n394), .A3(new_n401), .A4(new_n402), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n390), .A2(new_n391), .ZN(new_n404));
  OAI21_X1  g218(.A(KEYINPUT6), .B1(new_n390), .B2(new_n391), .ZN(new_n405));
  OR2_X1    g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n355), .A2(G953), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n407), .B(KEYINPUT84), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n354), .B(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n404), .A2(new_n405), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n406), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n403), .A2(new_n411), .A3(new_n274), .ZN(new_n412));
  OAI21_X1  g226(.A(G210), .B1(G237), .B2(G902), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n403), .A2(new_n411), .A3(new_n274), .A4(new_n413), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n328), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n192), .A2(G952), .ZN(new_n418));
  INV_X1    g232(.A(G234), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n418), .B1(new_n419), .B2(new_n191), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  OAI211_X1 g235(.A(G902), .B(G953), .C1(new_n419), .C2(new_n191), .ZN(new_n422));
  XOR2_X1   g236(.A(new_n422), .B(KEYINPUT99), .Z(new_n423));
  XNOR2_X1  g237(.A(KEYINPUT21), .B(G898), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n421), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n417), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G469), .ZN(new_n428));
  OAI21_X1  g242(.A(KEYINPUT81), .B1(new_n331), .B2(new_n334), .ZN(new_n429));
  OR2_X1    g243(.A1(new_n340), .A2(new_n329), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n330), .A2(new_n332), .A3(new_n333), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT69), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n329), .A2(KEYINPUT69), .A3(new_n330), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT81), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n429), .A2(new_n430), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n380), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT10), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT11), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n441), .B1(new_n299), .B2(G137), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n299), .A2(G137), .ZN(new_n443));
  INV_X1    g257(.A(G137), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(KEYINPUT11), .A3(G134), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n442), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT66), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT66), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n442), .A2(new_n445), .A3(new_n448), .A4(new_n443), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n447), .A2(G131), .A3(new_n449), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n442), .A2(new_n445), .A3(new_n247), .A4(new_n443), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT67), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n447), .A2(KEYINPUT67), .A3(G131), .A4(new_n449), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n346), .ZN(new_n457));
  INV_X1    g271(.A(new_n351), .ZN(new_n458));
  NOR3_X1   g272(.A1(new_n339), .A2(new_n349), .A3(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n457), .B1(new_n459), .B2(new_n344), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(new_n388), .A3(new_n386), .ZN(new_n461));
  INV_X1    g275(.A(new_n340), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n348), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n433), .A2(new_n434), .ZN(new_n464));
  AOI211_X1 g278(.A(new_n439), .B(new_n379), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n440), .A2(new_n456), .A3(new_n461), .A4(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(G110), .B(G140), .ZN(new_n468));
  INV_X1    g282(.A(G227), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n469), .A2(G953), .ZN(new_n470));
  XOR2_X1   g284(.A(new_n468), .B(new_n470), .Z(new_n471));
  NAND2_X1  g285(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT83), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n473), .B1(new_n341), .B2(new_n380), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT83), .A4(new_n379), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n438), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT12), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n456), .A2(KEYINPUT82), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n477), .B1(new_n476), .B2(new_n478), .ZN(new_n480));
  NOR3_X1   g294(.A1(new_n472), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n440), .A2(new_n461), .A3(new_n466), .ZN(new_n482));
  INV_X1    g296(.A(new_n456), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n471), .B1(new_n484), .B2(new_n467), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n428), .B(new_n274), .C1(new_n481), .C2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(G469), .A2(G902), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n437), .A2(new_n380), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n474), .A2(new_n475), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n478), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT12), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n491), .A2(new_n467), .A3(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n471), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n484), .A2(new_n467), .A3(new_n471), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n486), .B(new_n487), .C1(new_n428), .C2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G221), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n499), .B1(new_n313), .B2(new_n274), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  NOR3_X1   g316(.A1(new_n326), .A2(new_n427), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT68), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n504), .A2(new_n444), .A3(G134), .ZN(new_n505));
  OAI21_X1  g319(.A(KEYINPUT68), .B1(new_n444), .B2(G134), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n299), .A2(G137), .ZN(new_n507));
  OAI211_X1 g321(.A(G131), .B(new_n505), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT71), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n508), .A2(new_n509), .A3(new_n451), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n509), .B1(new_n508), .B2(new_n451), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n341), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT72), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n460), .A2(new_n454), .A3(new_n455), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n341), .B(KEYINPUT72), .C1(new_n510), .C2(new_n511), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT30), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT30), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n341), .A2(new_n451), .A3(new_n508), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n515), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n383), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n514), .A2(new_n515), .A3(new_n383), .A4(new_n516), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(G101), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n198), .A2(G210), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n528), .B(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n515), .A2(new_n512), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n534), .B(KEYINPUT74), .ZN(new_n535));
  AOI21_X1  g349(.A(KEYINPUT28), .B1(new_n535), .B2(new_n383), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT28), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n515), .A2(new_n520), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n523), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n537), .B1(new_n539), .B2(new_n525), .ZN(new_n540));
  NOR3_X1   g354(.A1(new_n536), .A2(new_n540), .A3(new_n531), .ZN(new_n541));
  NOR3_X1   g355(.A1(new_n533), .A2(new_n541), .A3(KEYINPUT29), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n517), .A2(new_n523), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n537), .B1(new_n543), .B2(new_n525), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n536), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n545), .A2(KEYINPUT29), .A3(new_n530), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n274), .ZN(new_n547));
  OAI21_X1  g361(.A(G472), .B1(new_n542), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n525), .A2(new_n530), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(KEYINPUT73), .B1(new_n524), .B2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n383), .B1(new_n518), .B2(new_n521), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT73), .ZN(new_n553));
  NOR3_X1   g367(.A1(new_n552), .A2(new_n553), .A3(new_n549), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT31), .B1(new_n551), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n531), .B1(new_n536), .B2(new_n540), .ZN(new_n556));
  NOR3_X1   g370(.A1(new_n552), .A2(KEYINPUT31), .A3(new_n549), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n555), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT32), .ZN(new_n560));
  NOR2_X1   g374(.A1(G472), .A2(G902), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n560), .B1(new_n559), .B2(new_n561), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n548), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(G217), .B1(new_n419), .B2(G902), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(KEYINPUT75), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n294), .A2(KEYINPUT23), .A3(G119), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT76), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n569), .B(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(KEYINPUT23), .B1(new_n294), .B2(G119), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT77), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n294), .A2(G119), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n360), .A2(G128), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT77), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(new_n576), .A3(KEYINPUT23), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n573), .A2(new_n574), .A3(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(G110), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n571), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  OR2_X1    g394(.A1(new_n580), .A2(KEYINPUT79), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n574), .A2(new_n575), .ZN(new_n582));
  XNOR2_X1  g396(.A(KEYINPUT24), .B(G110), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n580), .A2(KEYINPUT79), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n581), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n586), .A2(new_n236), .A3(new_n217), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n579), .B1(new_n571), .B2(new_n578), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n582), .A2(new_n583), .ZN(new_n589));
  OR3_X1    g403(.A1(new_n268), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n192), .A2(G221), .A3(G234), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(KEYINPUT22), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(G137), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n587), .A2(new_n590), .A3(new_n594), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(new_n274), .A3(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT25), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n598), .A2(new_n599), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n568), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n602), .B1(new_n568), .B2(new_n598), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT80), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT80), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n602), .B(new_n605), .C1(new_n568), .C2(new_n598), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n503), .A2(new_n565), .A3(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(G101), .ZN(G3));
  NAND2_X1  g423(.A1(new_n559), .A2(new_n561), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n553), .B1(new_n552), .B2(new_n549), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n515), .A2(new_n519), .A3(new_n520), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n612), .B1(KEYINPUT30), .B2(new_n517), .ZN(new_n613));
  OAI211_X1 g427(.A(KEYINPUT73), .B(new_n550), .C1(new_n613), .C2(new_n383), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n557), .B1(new_n615), .B2(KEYINPUT31), .ZN(new_n616));
  AOI21_X1  g430(.A(G902), .B1(new_n616), .B2(new_n556), .ZN(new_n617));
  INV_X1    g431(.A(G472), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n610), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n607), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n621), .A2(new_n502), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n319), .A2(new_n320), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n315), .A2(KEYINPUT33), .A3(new_n318), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n624), .A2(G478), .A3(new_n274), .A4(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n323), .A2(new_n285), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n284), .A2(KEYINPUT100), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(KEYINPUT100), .B1(new_n284), .B2(new_n628), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n629), .A2(new_n427), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n622), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT34), .B(G104), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G6));
  AND3_X1   g448(.A1(new_n277), .A2(new_n281), .A3(new_n283), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n325), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(new_n427), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n622), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT35), .B(G107), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  NOR2_X1   g454(.A1(new_n595), .A2(KEYINPUT36), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n591), .B(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n642), .A2(new_n274), .A3(new_n567), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n602), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n326), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n427), .A2(new_n502), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n645), .A2(new_n620), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT101), .B(KEYINPUT37), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G110), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n647), .B(new_n649), .ZN(G12));
  INV_X1    g464(.A(new_n502), .ZN(new_n651));
  INV_X1    g465(.A(G900), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n421), .B1(new_n423), .B2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n636), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n415), .A2(new_n416), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n327), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n644), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n565), .A2(new_n651), .A3(new_n654), .A4(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G128), .ZN(G30));
  INV_X1    g473(.A(new_n615), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n530), .B1(new_n543), .B2(new_n525), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n274), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(G472), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n663), .B1(new_n563), .B2(new_n564), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n664), .A2(KEYINPUT102), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n284), .A2(new_n325), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n644), .A2(new_n327), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n653), .B(KEYINPUT39), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n651), .A2(KEYINPUT40), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT40), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n672), .B1(new_n502), .B2(new_n669), .ZN(new_n673));
  AOI211_X1 g487(.A(new_n667), .B(new_n668), .C1(new_n671), .C2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n655), .B(KEYINPUT38), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n664), .A2(KEYINPUT102), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n666), .A2(new_n674), .A3(new_n675), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G143), .ZN(G45));
  NAND2_X1  g492(.A1(new_n610), .A2(KEYINPUT32), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n562), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n502), .B1(new_n680), .B2(new_n548), .ZN(new_n681));
  INV_X1    g495(.A(new_n653), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n284), .A2(new_n628), .A3(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n681), .A2(new_n657), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G146), .ZN(G48));
  INV_X1    g500(.A(new_n467), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n465), .B1(new_n438), .B2(new_n439), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n456), .B1(new_n688), .B2(new_n461), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n494), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n491), .A2(new_n467), .A3(new_n471), .A4(new_n492), .ZN(new_n691));
  AOI21_X1  g505(.A(G902), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(KEYINPUT103), .B1(new_n692), .B2(new_n428), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n274), .B1(new_n481), .B2(new_n485), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(G469), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n694), .A2(KEYINPUT103), .A3(G469), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n500), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n631), .A2(new_n565), .A3(new_n607), .A4(new_n698), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT41), .B(G113), .Z(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT104), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n699), .B(new_n701), .ZN(G15));
  NAND4_X1  g516(.A1(new_n565), .A2(new_n607), .A3(new_n637), .A4(new_n698), .ZN(new_n703));
  XOR2_X1   g517(.A(KEYINPUT105), .B(G116), .Z(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G18));
  INV_X1    g519(.A(new_n427), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n565), .A2(new_n645), .A3(new_n706), .A4(new_n698), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G119), .ZN(G21));
  INV_X1    g522(.A(KEYINPUT106), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n709), .B1(new_n667), .B2(new_n656), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n417), .A2(new_n325), .A3(KEYINPUT106), .A4(new_n284), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n618), .B1(new_n559), .B2(new_n274), .ZN(new_n713));
  INV_X1    g527(.A(new_n561), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n531), .B1(new_n536), .B2(new_n544), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n714), .B1(new_n616), .B2(new_n715), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n713), .A2(new_n603), .A3(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n712), .A2(new_n426), .A3(new_n698), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G122), .ZN(G24));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT103), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n486), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n692), .A2(new_n428), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n697), .ZN(new_n725));
  OAI211_X1 g539(.A(new_n417), .B(new_n501), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n683), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n713), .A2(new_n644), .A3(new_n716), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n720), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(new_n628), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n262), .A2(new_n263), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n254), .B1(new_n731), .B2(new_n187), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n278), .B1(new_n732), .B2(new_n264), .ZN(new_n733));
  NOR4_X1   g547(.A1(new_n733), .A2(new_n276), .A3(G475), .A4(G902), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT20), .B1(new_n282), .B2(new_n274), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n730), .B1(new_n736), .B2(new_n281), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n698), .A2(new_n737), .A3(new_n417), .A4(new_n682), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n555), .A2(new_n558), .A3(new_n715), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n561), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n602), .A2(new_n643), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n740), .B(new_n741), .C1(new_n617), .C2(new_n618), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n738), .A2(new_n742), .A3(KEYINPUT107), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n729), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(KEYINPUT108), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n219), .ZN(G27));
  AND2_X1   g560(.A1(new_n565), .A2(new_n607), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n415), .A2(new_n327), .A3(new_n416), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n683), .A2(new_n502), .A3(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n750), .A2(KEYINPUT42), .ZN(new_n751));
  INV_X1    g565(.A(new_n603), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n565), .A2(new_n752), .A3(new_n749), .ZN(new_n753));
  AOI22_X1  g567(.A1(new_n747), .A2(new_n751), .B1(new_n753), .B2(KEYINPUT42), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G131), .ZN(G33));
  AOI21_X1  g569(.A(new_n748), .B1(new_n604), .B2(new_n606), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n681), .A2(new_n654), .A3(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G134), .ZN(G36));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n277), .A2(new_n281), .A3(new_n628), .A4(new_n283), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT43), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n759), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n760), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT43), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n760), .A2(new_n761), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(KEYINPUT110), .A3(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n764), .A2(new_n768), .A3(new_n619), .A4(new_n741), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT44), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n748), .B1(new_n769), .B2(new_n770), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT45), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n497), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n495), .A2(KEYINPUT45), .A3(new_n496), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n774), .A2(G469), .A3(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n776), .A2(KEYINPUT46), .A3(new_n487), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n486), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT109), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT46), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n774), .A2(new_n775), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n781), .B(G469), .C1(new_n782), .C2(G902), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n777), .A2(KEYINPUT109), .A3(new_n486), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n780), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n785), .A2(new_n501), .A3(new_n670), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n771), .A2(new_n772), .A3(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G137), .ZN(G39));
  INV_X1    g602(.A(new_n565), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n607), .A2(new_n683), .A3(new_n748), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n785), .A2(KEYINPUT47), .A3(new_n501), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT47), .B1(new_n785), .B2(new_n501), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n789), .B(new_n790), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G140), .ZN(G42));
  NAND2_X1  g608(.A1(new_n754), .A2(new_n757), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n748), .A2(new_n653), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n565), .A2(new_n645), .A3(new_n651), .A4(new_n796), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n797), .A2(KEYINPUT111), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(KEYINPUT111), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n795), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n741), .A2(new_n653), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n712), .A2(new_n664), .A3(new_n651), .A4(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT113), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n502), .B1(new_n680), .B2(new_n663), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n805), .A2(KEYINPUT113), .A3(new_n712), .A4(new_n801), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n685), .B(new_n658), .C1(new_n743), .C2(new_n729), .ZN(new_n808));
  OAI21_X1  g622(.A(KEYINPUT52), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n718), .A2(new_n699), .A3(new_n703), .A4(new_n707), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n608), .A2(new_n647), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n636), .B1(new_n635), .B2(new_n730), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n646), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n621), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n750), .A2(new_n742), .ZN(new_n815));
  NOR4_X1   g629(.A1(new_n810), .A2(new_n811), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n658), .B1(new_n729), .B2(new_n743), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n804), .A2(new_n806), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT52), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n818), .A2(new_n819), .A3(new_n820), .A4(new_n685), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n800), .A2(new_n809), .A3(new_n816), .A4(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XOR2_X1   g638(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n825));
  OAI21_X1  g639(.A(new_n825), .B1(new_n807), .B2(new_n808), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n681), .A2(new_n657), .A3(new_n684), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n827), .B1(new_n817), .B2(KEYINPUT112), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT112), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n829), .B(new_n658), .C1(new_n729), .C2(new_n743), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n819), .A2(KEYINPUT52), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n826), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n810), .ZN(new_n834));
  INV_X1    g648(.A(new_n815), .ZN(new_n835));
  INV_X1    g649(.A(new_n811), .ZN(new_n836));
  INV_X1    g650(.A(new_n814), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n834), .A2(new_n835), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n798), .A2(new_n799), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n839), .A2(new_n754), .A3(new_n757), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n833), .A2(new_n841), .A3(KEYINPUT53), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n824), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n843), .A2(KEYINPUT54), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n420), .B1(new_n766), .B2(new_n767), .ZN(new_n846));
  INV_X1    g660(.A(new_n748), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n846), .A2(new_n698), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n848), .A2(new_n565), .A3(new_n752), .ZN(new_n849));
  NAND2_X1  g663(.A1(KEYINPUT116), .A2(KEYINPUT48), .ZN(new_n850));
  OR2_X1    g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n846), .A2(new_n717), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n852), .A2(new_n417), .A3(new_n698), .ZN(new_n853));
  OR2_X1    g667(.A1(KEYINPUT116), .A2(KEYINPUT48), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n849), .A2(new_n850), .A3(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n851), .A2(new_n418), .A3(new_n853), .A4(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n501), .B1(new_n696), .B2(new_n697), .ZN(new_n857));
  OR3_X1    g671(.A1(new_n791), .A2(new_n792), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n858), .A2(new_n847), .A3(new_n852), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n675), .A2(new_n327), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n852), .A2(new_n698), .A3(new_n860), .ZN(new_n861));
  XOR2_X1   g675(.A(new_n861), .B(KEYINPUT50), .Z(new_n862));
  AND2_X1   g676(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n756), .A2(new_n698), .ZN(new_n864));
  INV_X1    g678(.A(new_n676), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n421), .B(new_n864), .C1(new_n865), .C2(new_n665), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n866), .A2(new_n284), .A3(new_n628), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n867), .B1(new_n728), .B2(new_n848), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT51), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n856), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n870), .B1(new_n868), .B2(KEYINPUT115), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n872), .B(new_n863), .C1(KEYINPUT115), .C2(new_n868), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n822), .A2(new_n823), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT53), .B1(new_n833), .B2(new_n841), .ZN(new_n875));
  OAI21_X1  g689(.A(KEYINPUT54), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n845), .A2(new_n871), .A3(new_n873), .A4(new_n876), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n866), .A2(new_n630), .A3(new_n629), .ZN(new_n878));
  OAI22_X1  g692(.A1(new_n877), .A2(new_n878), .B1(G952), .B2(G953), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n696), .A2(new_n697), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT49), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n752), .ZN(new_n882));
  NOR4_X1   g696(.A1(new_n882), .A2(new_n328), .A3(new_n500), .A4(new_n675), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n883), .B(new_n765), .C1(new_n865), .C2(new_n665), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n879), .A2(new_n884), .ZN(G75));
  NAND2_X1  g699(.A1(new_n406), .A2(new_n410), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n886), .B(new_n409), .Z(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT55), .ZN(new_n888));
  INV_X1    g702(.A(G210), .ZN(new_n889));
  AOI211_X1 g703(.A(new_n889), .B(new_n274), .C1(new_n824), .C2(new_n842), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n888), .B1(new_n890), .B2(KEYINPUT56), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n274), .B1(new_n824), .B2(new_n842), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(G210), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT56), .ZN(new_n894));
  INV_X1    g708(.A(new_n888), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n192), .A2(G952), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n891), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT117), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n891), .A2(new_n896), .A3(KEYINPUT117), .A4(new_n898), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(G51));
  NAND2_X1  g717(.A1(new_n487), .A2(KEYINPUT57), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n843), .A2(KEYINPUT54), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n904), .B1(new_n905), .B2(new_n844), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n487), .A2(KEYINPUT57), .ZN(new_n907));
  OAI22_X1  g721(.A1(new_n906), .A2(new_n907), .B1(new_n485), .B2(new_n481), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n892), .A2(G469), .A3(new_n782), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n897), .B1(new_n908), .B2(new_n909), .ZN(G54));
  NAND3_X1  g724(.A1(new_n892), .A2(KEYINPUT58), .A3(G475), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n733), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n892), .A2(KEYINPUT58), .A3(G475), .A4(new_n272), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n912), .A2(new_n898), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(KEYINPUT118), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT118), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n912), .A2(new_n916), .A3(new_n898), .A4(new_n913), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n915), .A2(new_n917), .ZN(G60));
  AND2_X1   g732(.A1(new_n624), .A2(new_n625), .ZN(new_n919));
  NAND2_X1  g733(.A1(G478), .A2(G902), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT59), .Z(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n919), .B(new_n922), .C1(new_n905), .C2(new_n844), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n921), .B1(new_n845), .B2(new_n876), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n923), .B(new_n898), .C1(new_n924), .C2(new_n919), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(G63));
  NAND2_X1  g740(.A1(G217), .A2(G902), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT60), .Z(new_n928));
  NAND3_X1  g742(.A1(new_n843), .A2(new_n642), .A3(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n929), .A2(KEYINPUT119), .A3(new_n898), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(KEYINPUT61), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n843), .A2(new_n928), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n596), .A2(new_n597), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n898), .B(new_n929), .C1(new_n932), .C2(new_n933), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n931), .B(new_n934), .ZN(G66));
  OAI21_X1  g749(.A(G953), .B1(new_n355), .B2(new_n424), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n810), .A2(new_n811), .A3(new_n814), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n936), .B1(new_n937), .B2(G953), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n886), .B1(G898), .B2(new_n192), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT120), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n938), .B(new_n940), .ZN(G69));
  NAND2_X1  g755(.A1(new_n227), .A2(new_n229), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n522), .B(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n943), .A2(G953), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT121), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n817), .A2(KEYINPUT112), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n946), .A2(new_n677), .A3(new_n685), .A4(new_n830), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT62), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n828), .A2(KEYINPUT62), .A3(new_n677), .A4(new_n830), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n747), .A2(new_n812), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n502), .A2(new_n669), .A3(new_n748), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n793), .A2(new_n787), .A3(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n945), .B1(new_n951), .B2(new_n956), .ZN(new_n957));
  AOI211_X1 g771(.A(KEYINPUT121), .B(new_n955), .C1(new_n949), .C2(new_n950), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n944), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n192), .A2(G900), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT122), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n793), .A2(new_n787), .ZN(new_n962));
  AND4_X1   g776(.A1(new_n565), .A2(new_n786), .A3(new_n752), .A4(new_n712), .ZN(new_n963));
  NOR4_X1   g777(.A1(new_n831), .A2(new_n962), .A3(new_n795), .A4(new_n963), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n943), .B(new_n961), .C1(new_n964), .C2(G953), .ZN(new_n965));
  OAI21_X1  g779(.A(G953), .B1(new_n469), .B2(new_n652), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT123), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n959), .A2(new_n965), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(KEYINPUT124), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT124), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n959), .A2(new_n971), .A3(new_n965), .A4(new_n968), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n966), .A2(new_n967), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n970), .A2(new_n974), .A3(new_n972), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(G72));
  INV_X1    g792(.A(KEYINPUT127), .ZN(new_n979));
  XNOR2_X1  g793(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n618), .A2(new_n274), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n980), .B(new_n981), .Z(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n983), .B1(new_n964), .B2(new_n937), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n526), .B(KEYINPUT126), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  NOR3_X1   g800(.A1(new_n984), .A2(new_n530), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n979), .B1(new_n987), .B2(new_n897), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n964), .A2(new_n937), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n531), .B(new_n985), .C1(new_n989), .C2(new_n983), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n990), .A2(KEYINPUT127), .A3(new_n898), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n988), .A2(new_n991), .ZN(new_n992));
  OAI221_X1 g806(.A(new_n982), .B1(new_n660), .B2(new_n533), .C1(new_n874), .C2(new_n875), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n957), .A2(new_n958), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n994), .A2(new_n937), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n530), .B(new_n986), .C1(new_n995), .C2(new_n983), .ZN(new_n996));
  AND3_X1   g810(.A1(new_n992), .A2(new_n993), .A3(new_n996), .ZN(G57));
endmodule


