

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730;

  XNOR2_X1 U368 ( .A(n432), .B(n397), .ZN(n717) );
  NOR2_X2 U369 ( .A1(G953), .A2(G237), .ZN(n485) );
  XNOR2_X1 U370 ( .A(n399), .B(G146), .ZN(n432) );
  XNOR2_X1 U371 ( .A(n364), .B(n389), .ZN(n596) );
  OR2_X1 U372 ( .A1(n598), .A2(KEYINPUT2), .ZN(n599) );
  XNOR2_X2 U373 ( .A(n480), .B(n481), .ZN(n501) );
  NOR2_X2 U374 ( .A1(n497), .A2(n496), .ZN(n347) );
  XNOR2_X2 U375 ( .A(n472), .B(G469), .ZN(n554) );
  NOR2_X1 U376 ( .A1(n619), .A2(n701), .ZN(n620) );
  NOR2_X1 U377 ( .A1(n626), .A2(n701), .ZN(n627) );
  NAND2_X1 U378 ( .A1(n596), .A2(n595), .ZN(n721) );
  XNOR2_X1 U379 ( .A(n505), .B(KEYINPUT33), .ZN(n659) );
  INV_X2 U380 ( .A(G953), .ZN(n723) );
  NAND2_X1 U381 ( .A1(n540), .A2(n539), .ZN(n542) );
  NOR2_X1 U382 ( .A1(n538), .A2(n537), .ZN(n539) );
  AND2_X1 U383 ( .A1(n580), .A2(n357), .ZN(n560) );
  NOR2_X1 U384 ( .A1(n601), .A2(G902), .ZN(n481) );
  XNOR2_X1 U385 ( .A(n347), .B(n348), .ZN(n728) );
  XOR2_X1 U386 ( .A(n404), .B(KEYINPUT32), .Z(n348) );
  AND2_X4 U387 ( .A1(n600), .A2(n599), .ZN(n697) );
  XNOR2_X1 U388 ( .A(G119), .B(KEYINPUT3), .ZN(n410) );
  XNOR2_X1 U389 ( .A(n450), .B(n375), .ZN(n370) );
  XNOR2_X1 U390 ( .A(KEYINPUT71), .B(KEYINPUT4), .ZN(n375) );
  INV_X1 U391 ( .A(G125), .ZN(n399) );
  XNOR2_X1 U392 ( .A(n416), .B(n415), .ZN(n417) );
  AND2_X1 U393 ( .A1(n632), .A2(n351), .ZN(n369) );
  XNOR2_X1 U394 ( .A(n445), .B(n396), .ZN(n474) );
  INV_X1 U395 ( .A(KEYINPUT8), .ZN(n396) );
  XNOR2_X1 U396 ( .A(n466), .B(n412), .ZN(n403) );
  XNOR2_X1 U397 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n412) );
  XNOR2_X1 U398 ( .A(n401), .B(KEYINPUT96), .ZN(n400) );
  OR2_X1 U399 ( .A1(n693), .A2(G902), .ZN(n472) );
  XNOR2_X1 U400 ( .A(n552), .B(n493), .ZN(n562) );
  XOR2_X1 U401 ( .A(KEYINPUT16), .B(G122), .Z(n409) );
  XNOR2_X1 U402 ( .A(G137), .B(KEYINPUT24), .ZN(n475) );
  NAND2_X1 U403 ( .A1(n474), .A2(G221), .ZN(n395) );
  XNOR2_X1 U404 ( .A(n350), .B(n477), .ZN(n393) );
  XNOR2_X1 U405 ( .A(KEYINPUT10), .B(G140), .ZN(n397) );
  XNOR2_X1 U406 ( .A(n721), .B(n376), .ZN(n597) );
  INV_X1 U407 ( .A(KEYINPUT77), .ZN(n376) );
  XNOR2_X1 U408 ( .A(n363), .B(KEYINPUT15), .ZN(n593) );
  XNOR2_X1 U409 ( .A(G902), .B(KEYINPUT95), .ZN(n363) );
  XNOR2_X1 U410 ( .A(n716), .B(n467), .ZN(n489) );
  NOR2_X1 U411 ( .A1(n628), .A2(KEYINPUT2), .ZN(n388) );
  XNOR2_X1 U412 ( .A(n421), .B(KEYINPUT92), .ZN(n561) );
  XOR2_X1 U413 ( .A(KEYINPUT22), .B(KEYINPUT73), .Z(n462) );
  AND2_X1 U414 ( .A1(n551), .A2(n635), .ZN(n405) );
  NOR2_X1 U415 ( .A1(n630), .A2(n383), .ZN(n382) );
  XNOR2_X1 U416 ( .A(n479), .B(KEYINPUT25), .ZN(n480) );
  INV_X1 U417 ( .A(n497), .ZN(n384) );
  NOR2_X1 U418 ( .A1(G237), .A2(G902), .ZN(n414) );
  XNOR2_X1 U419 ( .A(n482), .B(KEYINPUT5), .ZN(n483) );
  OR2_X1 U420 ( .A1(n668), .A2(n534), .ZN(n538) );
  XNOR2_X1 U421 ( .A(G134), .B(G131), .ZN(n464) );
  NAND2_X1 U422 ( .A1(G237), .A2(G234), .ZN(n423) );
  INV_X1 U423 ( .A(KEYINPUT48), .ZN(n389) );
  NOR2_X1 U424 ( .A1(n577), .A2(n368), .ZN(n367) );
  AND2_X1 U425 ( .A1(n377), .A2(n562), .ZN(n582) );
  XNOR2_X1 U426 ( .A(n457), .B(n456), .ZN(n645) );
  XNOR2_X1 U427 ( .A(n429), .B(KEYINPUT0), .ZN(n430) );
  XOR2_X1 U428 ( .A(G134), .B(G122), .Z(n449) );
  XNOR2_X1 U429 ( .A(G116), .B(G107), .ZN(n448) );
  XOR2_X1 U430 ( .A(KEYINPUT11), .B(KEYINPUT103), .Z(n434) );
  XNOR2_X1 U431 ( .A(G113), .B(G104), .ZN(n436) );
  XOR2_X1 U432 ( .A(KEYINPUT12), .B(G122), .Z(n437) );
  XNOR2_X1 U433 ( .A(G143), .B(G131), .ZN(n438) );
  XNOR2_X1 U434 ( .A(n402), .B(n398), .ZN(n413) );
  XNOR2_X1 U435 ( .A(n400), .B(n432), .ZN(n398) );
  XNOR2_X1 U436 ( .A(n370), .B(n403), .ZN(n402) );
  AND2_X1 U437 ( .A1(n527), .A2(n630), .ZN(n504) );
  XNOR2_X1 U438 ( .A(n582), .B(KEYINPUT113), .ZN(n564) );
  XNOR2_X1 U439 ( .A(n557), .B(KEYINPUT78), .ZN(n390) );
  AND2_X1 U440 ( .A1(n556), .A2(n351), .ZN(n557) );
  XNOR2_X1 U441 ( .A(n561), .B(n422), .ZN(n569) );
  OR2_X1 U442 ( .A1(n361), .A2(n360), .ZN(n568) );
  INV_X1 U443 ( .A(n554), .ZN(n360) );
  XNOR2_X1 U444 ( .A(n553), .B(n362), .ZN(n361) );
  INV_X1 U445 ( .A(KEYINPUT28), .ZN(n362) );
  AND2_X1 U446 ( .A1(n527), .A2(n554), .ZN(n556) );
  OR2_X1 U447 ( .A1(n607), .A2(G902), .ZN(n492) );
  INV_X1 U448 ( .A(n562), .ZN(n374) );
  XNOR2_X1 U449 ( .A(n394), .B(n392), .ZN(n601) );
  XNOR2_X1 U450 ( .A(n393), .B(n476), .ZN(n392) );
  XNOR2_X1 U451 ( .A(n717), .B(n395), .ZN(n394) );
  XNOR2_X1 U452 ( .A(n386), .B(n385), .ZN(n665) );
  INV_X1 U453 ( .A(KEYINPUT85), .ZN(n385) );
  INV_X1 U454 ( .A(KEYINPUT65), .ZN(n404) );
  BUF_X1 U455 ( .A(G128), .Z(n359) );
  NOR2_X1 U456 ( .A1(n568), .A2(n569), .ZN(n680) );
  NAND2_X1 U457 ( .A1(n349), .A2(n378), .ZN(n675) );
  NAND2_X1 U458 ( .A1(n384), .A2(n382), .ZN(n378) );
  AND2_X1 U459 ( .A1(n381), .A2(n405), .ZN(n380) );
  AND2_X1 U460 ( .A1(n371), .A2(n501), .ZN(n668) );
  XNOR2_X1 U461 ( .A(n372), .B(KEYINPUT89), .ZN(n371) );
  NAND2_X1 U462 ( .A1(n384), .A2(n373), .ZN(n372) );
  AND2_X1 U463 ( .A1(n585), .A2(n374), .ZN(n373) );
  AND2_X1 U464 ( .A1(n379), .A2(n380), .ZN(n349) );
  XOR2_X1 U465 ( .A(G119), .B(G110), .Z(n350) );
  OR2_X1 U466 ( .A1(n550), .A2(n549), .ZN(n351) );
  XOR2_X1 U467 ( .A(G113), .B(G116), .Z(n352) );
  XOR2_X1 U468 ( .A(KEYINPUT38), .B(n544), .Z(n353) );
  AND2_X1 U469 ( .A1(n559), .A2(n353), .ZN(n354) );
  OR2_X1 U470 ( .A1(n645), .A2(n461), .ZN(n355) );
  OR2_X1 U471 ( .A1(KEYINPUT47), .A2(n576), .ZN(n356) );
  AND2_X1 U472 ( .A1(n531), .A2(n530), .ZN(n357) );
  INV_X1 U473 ( .A(n501), .ZN(n551) );
  XOR2_X1 U474 ( .A(KEYINPUT46), .B(KEYINPUT87), .Z(n358) );
  XNOR2_X1 U475 ( .A(n709), .B(n413), .ZN(n621) );
  NOR2_X1 U476 ( .A1(n593), .A2(n621), .ZN(n418) );
  XNOR2_X1 U477 ( .A(n498), .B(KEYINPUT91), .ZN(n522) );
  AND2_X2 U478 ( .A1(n629), .A2(n593), .ZN(n600) );
  NAND2_X1 U479 ( .A1(n723), .A2(G224), .ZN(n401) );
  NAND2_X1 U480 ( .A1(n570), .A2(n680), .ZN(n576) );
  NAND2_X1 U481 ( .A1(n367), .A2(n365), .ZN(n364) );
  XNOR2_X1 U482 ( .A(n366), .B(n358), .ZN(n365) );
  NOR2_X2 U483 ( .A1(n729), .A2(n730), .ZN(n366) );
  NAND2_X1 U484 ( .A1(n578), .A2(n356), .ZN(n368) );
  AND2_X1 U485 ( .A1(n369), .A2(n551), .ZN(n563) );
  XNOR2_X1 U486 ( .A(n370), .B(n465), .ZN(n716) );
  XNOR2_X2 U487 ( .A(G143), .B(G128), .ZN(n450) );
  AND2_X1 U488 ( .A1(n563), .A2(n357), .ZN(n377) );
  NAND2_X1 U489 ( .A1(n728), .A2(n675), .ZN(n498) );
  NAND2_X1 U490 ( .A1(n497), .A2(n383), .ZN(n379) );
  NAND2_X1 U491 ( .A1(n630), .A2(n383), .ZN(n381) );
  INV_X1 U492 ( .A(KEYINPUT109), .ZN(n383) );
  NAND2_X1 U493 ( .A1(n387), .A2(n629), .ZN(n386) );
  XNOR2_X1 U494 ( .A(n388), .B(KEYINPUT83), .ZN(n387) );
  XNOR2_X2 U495 ( .A(n463), .B(n462), .ZN(n497) );
  XNOR2_X2 U496 ( .A(n513), .B(n512), .ZN(n614) );
  XNOR2_X2 U497 ( .A(n554), .B(n473), .ZN(n630) );
  NAND2_X1 U498 ( .A1(n390), .A2(n559), .ZN(n571) );
  NAND2_X1 U499 ( .A1(n390), .A2(n354), .ZN(n391) );
  XNOR2_X2 U500 ( .A(n391), .B(KEYINPUT39), .ZN(n580) );
  OR2_X2 U501 ( .A1(n702), .A2(n592), .ZN(n629) );
  XNOR2_X2 U502 ( .A(n542), .B(n541), .ZN(n702) );
  XNOR2_X2 U503 ( .A(KEYINPUT68), .B(G101), .ZN(n466) );
  OR2_X1 U504 ( .A1(n550), .A2(n427), .ZN(n406) );
  XNOR2_X1 U505 ( .A(n609), .B(n608), .ZN(n407) );
  INV_X1 U506 ( .A(n632), .ZN(n461) );
  XNOR2_X1 U507 ( .A(n484), .B(n483), .ZN(n487) );
  INV_X1 U508 ( .A(KEYINPUT108), .ZN(n456) );
  INV_X1 U509 ( .A(KEYINPUT81), .ZN(n415) );
  XNOR2_X1 U510 ( .A(n470), .B(n409), .ZN(n411) );
  XNOR2_X1 U511 ( .A(n411), .B(n484), .ZN(n709) );
  INV_X1 U512 ( .A(n701), .ZN(n611) );
  INV_X1 U513 ( .A(KEYINPUT123), .ZN(n605) );
  XNOR2_X2 U514 ( .A(G110), .B(G107), .ZN(n408) );
  XNOR2_X2 U515 ( .A(n408), .B(G104), .ZN(n470) );
  XNOR2_X1 U516 ( .A(n352), .B(n410), .ZN(n484) );
  XNOR2_X1 U517 ( .A(n414), .B(KEYINPUT75), .ZN(n419) );
  NAND2_X1 U518 ( .A1(G210), .A2(n419), .ZN(n416) );
  XNOR2_X1 U519 ( .A(n418), .B(n417), .ZN(n543) );
  NAND2_X1 U520 ( .A1(n419), .A2(G214), .ZN(n420) );
  XNOR2_X1 U521 ( .A(n420), .B(KEYINPUT97), .ZN(n583) );
  INV_X1 U522 ( .A(n583), .ZN(n642) );
  NAND2_X1 U523 ( .A1(n543), .A2(n642), .ZN(n421) );
  XNOR2_X1 U524 ( .A(KEYINPUT19), .B(KEYINPUT67), .ZN(n422) );
  INV_X1 U525 ( .A(n569), .ZN(n428) );
  XNOR2_X1 U526 ( .A(n423), .B(KEYINPUT14), .ZN(n424) );
  XNOR2_X1 U527 ( .A(KEYINPUT74), .B(n424), .ZN(n426) );
  NAND2_X1 U528 ( .A1(G952), .A2(n426), .ZN(n656) );
  NOR2_X1 U529 ( .A1(G953), .A2(n656), .ZN(n550) );
  XOR2_X1 U530 ( .A(G898), .B(KEYINPUT98), .Z(n706) );
  NAND2_X1 U531 ( .A1(n706), .A2(G953), .ZN(n425) );
  XOR2_X1 U532 ( .A(KEYINPUT99), .B(n425), .Z(n710) );
  NAND2_X1 U533 ( .A1(G902), .A2(n426), .ZN(n546) );
  NOR2_X1 U534 ( .A1(n710), .A2(n546), .ZN(n427) );
  NAND2_X1 U535 ( .A1(n428), .A2(n406), .ZN(n431) );
  INV_X1 U536 ( .A(KEYINPUT93), .ZN(n429) );
  XNOR2_X1 U537 ( .A(n431), .B(n430), .ZN(n499) );
  XNOR2_X1 U538 ( .A(KEYINPUT13), .B(G475), .ZN(n444) );
  NAND2_X1 U539 ( .A1(G214), .A2(n485), .ZN(n433) );
  XNOR2_X1 U540 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U541 ( .A(n435), .B(KEYINPUT104), .Z(n441) );
  XNOR2_X1 U542 ( .A(n437), .B(n436), .ZN(n439) );
  XNOR2_X1 U543 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U544 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U545 ( .A(n717), .B(n442), .ZN(n615) );
  NOR2_X1 U546 ( .A1(G902), .A2(n615), .ZN(n443) );
  XNOR2_X1 U547 ( .A(n444), .B(n443), .ZN(n531) );
  XOR2_X1 U548 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n447) );
  NAND2_X1 U549 ( .A1(G234), .A2(n723), .ZN(n445) );
  NAND2_X1 U550 ( .A1(G217), .A2(n474), .ZN(n446) );
  XNOR2_X1 U551 ( .A(n447), .B(n446), .ZN(n454) );
  XNOR2_X1 U552 ( .A(n449), .B(n448), .ZN(n452) );
  XOR2_X1 U553 ( .A(KEYINPUT105), .B(n450), .Z(n451) );
  XNOR2_X1 U554 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U555 ( .A(n454), .B(n453), .ZN(n698) );
  NOR2_X1 U556 ( .A1(G902), .A2(n698), .ZN(n455) );
  XNOR2_X1 U557 ( .A(G478), .B(n455), .ZN(n530) );
  INV_X1 U558 ( .A(n530), .ZN(n508) );
  NOR2_X1 U559 ( .A1(n531), .A2(n508), .ZN(n457) );
  INV_X1 U560 ( .A(n593), .ZN(n458) );
  NAND2_X1 U561 ( .A1(G234), .A2(n458), .ZN(n459) );
  XNOR2_X1 U562 ( .A(KEYINPUT20), .B(n459), .ZN(n478) );
  NAND2_X1 U563 ( .A1(n478), .A2(G221), .ZN(n460) );
  XOR2_X1 U564 ( .A(KEYINPUT21), .B(n460), .Z(n632) );
  OR2_X2 U565 ( .A1(n499), .A2(n355), .ZN(n463) );
  XNOR2_X1 U566 ( .A(n464), .B(G137), .ZN(n465) );
  XNOR2_X1 U567 ( .A(n466), .B(G146), .ZN(n467) );
  NAND2_X1 U568 ( .A1(n723), .A2(G227), .ZN(n468) );
  XNOR2_X1 U569 ( .A(n468), .B(G140), .ZN(n469) );
  XNOR2_X1 U570 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U571 ( .A(n489), .B(n471), .ZN(n693) );
  XNOR2_X1 U572 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n473) );
  XNOR2_X1 U573 ( .A(n475), .B(n359), .ZN(n476) );
  XNOR2_X1 U574 ( .A(KEYINPUT23), .B(KEYINPUT100), .ZN(n477) );
  NAND2_X1 U575 ( .A1(G217), .A2(n478), .ZN(n479) );
  XOR2_X1 U576 ( .A(KEYINPUT76), .B(KEYINPUT101), .Z(n482) );
  NAND2_X1 U577 ( .A1(n485), .A2(G210), .ZN(n486) );
  XNOR2_X1 U578 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U579 ( .A(n489), .B(n488), .ZN(n607) );
  XNOR2_X1 U580 ( .A(G472), .B(KEYINPUT72), .ZN(n490) );
  XNOR2_X1 U581 ( .A(n490), .B(KEYINPUT102), .ZN(n491) );
  XNOR2_X2 U582 ( .A(n492), .B(n491), .ZN(n552) );
  INV_X1 U583 ( .A(n552), .ZN(n635) );
  INV_X1 U584 ( .A(KEYINPUT6), .ZN(n493) );
  NAND2_X1 U585 ( .A1(n630), .A2(n551), .ZN(n494) );
  NOR2_X1 U586 ( .A1(n562), .A2(n494), .ZN(n495) );
  XOR2_X1 U587 ( .A(KEYINPUT80), .B(n495), .Z(n496) );
  BUF_X1 U588 ( .A(n499), .Z(n500) );
  INV_X1 U589 ( .A(n500), .ZN(n528) );
  NAND2_X1 U590 ( .A1(n501), .A2(n632), .ZN(n503) );
  INV_X1 U591 ( .A(KEYINPUT70), .ZN(n502) );
  XNOR2_X2 U592 ( .A(n503), .B(n502), .ZN(n527) );
  NAND2_X1 U593 ( .A1(n504), .A2(n562), .ZN(n505) );
  NAND2_X1 U594 ( .A1(n528), .A2(n659), .ZN(n507) );
  XNOR2_X1 U595 ( .A(KEYINPUT79), .B(KEYINPUT34), .ZN(n506) );
  XNOR2_X1 U596 ( .A(n507), .B(n506), .ZN(n511) );
  NAND2_X1 U597 ( .A1(n508), .A2(n531), .ZN(n509) );
  XNOR2_X1 U598 ( .A(n509), .B(KEYINPUT110), .ZN(n572) );
  INV_X1 U599 ( .A(n572), .ZN(n510) );
  NAND2_X1 U600 ( .A1(n511), .A2(n510), .ZN(n513) );
  XNOR2_X1 U601 ( .A(KEYINPUT86), .B(KEYINPUT35), .ZN(n512) );
  XNOR2_X1 U602 ( .A(n614), .B(KEYINPUT69), .ZN(n514) );
  NAND2_X1 U603 ( .A1(n522), .A2(n514), .ZN(n516) );
  INV_X1 U604 ( .A(KEYINPUT44), .ZN(n515) );
  NAND2_X1 U605 ( .A1(n516), .A2(n515), .ZN(n524) );
  INV_X1 U606 ( .A(n614), .ZN(n535) );
  INV_X1 U607 ( .A(KEYINPUT90), .ZN(n517) );
  NOR2_X1 U608 ( .A1(n535), .A2(n517), .ZN(n520) );
  INV_X1 U609 ( .A(KEYINPUT69), .ZN(n518) );
  NAND2_X1 U610 ( .A1(n518), .A2(KEYINPUT44), .ZN(n519) );
  NOR2_X1 U611 ( .A1(n520), .A2(n519), .ZN(n521) );
  NAND2_X1 U612 ( .A1(n522), .A2(n521), .ZN(n523) );
  NAND2_X1 U613 ( .A1(n524), .A2(n523), .ZN(n540) );
  AND2_X1 U614 ( .A1(n527), .A2(n552), .ZN(n525) );
  AND2_X1 U615 ( .A1(n525), .A2(n630), .ZN(n638) );
  NAND2_X1 U616 ( .A1(n528), .A2(n638), .ZN(n526) );
  XNOR2_X1 U617 ( .A(n526), .B(KEYINPUT31), .ZN(n684) );
  NAND2_X1 U618 ( .A1(n528), .A2(n556), .ZN(n529) );
  NOR2_X1 U619 ( .A1(n552), .A2(n529), .ZN(n670) );
  NOR2_X1 U620 ( .A1(n684), .A2(n670), .ZN(n533) );
  NOR2_X1 U621 ( .A1(n531), .A2(n530), .ZN(n683) );
  XNOR2_X1 U622 ( .A(KEYINPUT106), .B(n683), .ZN(n579) );
  OR2_X1 U623 ( .A1(n357), .A2(n579), .ZN(n532) );
  XOR2_X1 U624 ( .A(KEYINPUT107), .B(n532), .Z(n570) );
  INV_X1 U625 ( .A(n570), .ZN(n647) );
  NOR2_X1 U626 ( .A1(n533), .A2(n647), .ZN(n534) );
  NOR2_X1 U627 ( .A1(n535), .A2(n515), .ZN(n536) );
  NOR2_X1 U628 ( .A1(n536), .A2(KEYINPUT90), .ZN(n537) );
  XOR2_X1 U629 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n541) );
  BUF_X1 U630 ( .A(n543), .Z(n544) );
  NAND2_X1 U631 ( .A1(n353), .A2(n642), .ZN(n646) );
  NOR2_X1 U632 ( .A1(n646), .A2(n645), .ZN(n545) );
  XNOR2_X1 U633 ( .A(n545), .B(KEYINPUT41), .ZN(n658) );
  NOR2_X1 U634 ( .A1(G900), .A2(n546), .ZN(n547) );
  NAND2_X1 U635 ( .A1(G953), .A2(n547), .ZN(n548) );
  XNOR2_X1 U636 ( .A(KEYINPUT111), .B(n548), .ZN(n549) );
  AND2_X1 U637 ( .A1(n552), .A2(n563), .ZN(n553) );
  NOR2_X1 U638 ( .A1(n658), .A2(n568), .ZN(n555) );
  XNOR2_X1 U639 ( .A(n555), .B(KEYINPUT42), .ZN(n730) );
  NOR2_X1 U640 ( .A1(n583), .A2(n635), .ZN(n558) );
  XNOR2_X1 U641 ( .A(n558), .B(KEYINPUT30), .ZN(n559) );
  XNOR2_X2 U642 ( .A(n560), .B(KEYINPUT40), .ZN(n729) );
  BUF_X1 U643 ( .A(n561), .Z(n565) );
  NOR2_X1 U644 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U645 ( .A(KEYINPUT36), .B(n566), .ZN(n567) );
  NAND2_X1 U646 ( .A1(n567), .A2(n630), .ZN(n687) );
  XNOR2_X1 U647 ( .A(n687), .B(KEYINPUT88), .ZN(n578) );
  NAND2_X1 U648 ( .A1(n576), .A2(KEYINPUT47), .ZN(n574) );
  NOR2_X1 U649 ( .A1(n572), .A2(n571), .ZN(n573) );
  NAND2_X1 U650 ( .A1(n544), .A2(n573), .ZN(n679) );
  NAND2_X1 U651 ( .A1(n574), .A2(n679), .ZN(n575) );
  XNOR2_X1 U652 ( .A(n575), .B(KEYINPUT84), .ZN(n577) );
  NAND2_X1 U653 ( .A1(n580), .A2(n579), .ZN(n689) );
  NAND2_X1 U654 ( .A1(n689), .A2(KEYINPUT2), .ZN(n581) );
  XNOR2_X1 U655 ( .A(n581), .B(KEYINPUT82), .ZN(n590) );
  INV_X1 U656 ( .A(n582), .ZN(n584) );
  NOR2_X1 U657 ( .A1(n584), .A2(n583), .ZN(n586) );
  INV_X1 U658 ( .A(n630), .ZN(n585) );
  NAND2_X1 U659 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U660 ( .A(KEYINPUT43), .B(n587), .ZN(n588) );
  XOR2_X1 U661 ( .A(KEYINPUT112), .B(n588), .Z(n589) );
  NOR2_X1 U662 ( .A1(n589), .A2(n544), .ZN(n690) );
  NOR2_X1 U663 ( .A1(n590), .A2(n690), .ZN(n591) );
  NAND2_X1 U664 ( .A1(n596), .A2(n591), .ZN(n592) );
  INV_X1 U665 ( .A(n689), .ZN(n594) );
  NOR2_X1 U666 ( .A1(n594), .A2(n690), .ZN(n595) );
  NOR2_X1 U667 ( .A1(n702), .A2(n597), .ZN(n598) );
  NAND2_X1 U668 ( .A1(n697), .A2(G217), .ZN(n602) );
  XNOR2_X1 U669 ( .A(n602), .B(n601), .ZN(n604) );
  INV_X1 U670 ( .A(G952), .ZN(n603) );
  AND2_X1 U671 ( .A1(n603), .A2(G953), .ZN(n701) );
  NOR2_X2 U672 ( .A1(n604), .A2(n701), .ZN(n606) );
  XNOR2_X1 U673 ( .A(n606), .B(n605), .ZN(G66) );
  NAND2_X1 U674 ( .A1(n697), .A2(G472), .ZN(n610) );
  XOR2_X1 U675 ( .A(KEYINPUT62), .B(KEYINPUT94), .Z(n609) );
  XNOR2_X1 U676 ( .A(n607), .B(KEYINPUT114), .ZN(n608) );
  XNOR2_X1 U677 ( .A(n610), .B(n407), .ZN(n612) );
  NAND2_X1 U678 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U679 ( .A(n613), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U680 ( .A(G122), .B(n614), .Z(G24) );
  NAND2_X1 U681 ( .A1(n697), .A2(G475), .ZN(n618) );
  XOR2_X1 U682 ( .A(KEYINPUT122), .B(KEYINPUT59), .Z(n616) );
  XNOR2_X1 U683 ( .A(n615), .B(n616), .ZN(n617) );
  XNOR2_X1 U684 ( .A(n618), .B(n617), .ZN(n619) );
  XNOR2_X1 U685 ( .A(n620), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U686 ( .A1(n697), .A2(G210), .ZN(n625) );
  BUF_X1 U687 ( .A(n621), .Z(n623) );
  XOR2_X1 U688 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n622) );
  XNOR2_X1 U689 ( .A(n623), .B(n622), .ZN(n624) );
  XNOR2_X1 U690 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U691 ( .A(n627), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X1 U692 ( .A1(n702), .A2(n721), .ZN(n628) );
  NOR2_X1 U693 ( .A1(n527), .A2(n630), .ZN(n631) );
  XNOR2_X1 U694 ( .A(n631), .B(KEYINPUT50), .ZN(n637) );
  NOR2_X1 U695 ( .A1(n501), .A2(n632), .ZN(n633) );
  XNOR2_X1 U696 ( .A(n633), .B(KEYINPUT49), .ZN(n634) );
  NAND2_X1 U697 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U698 ( .A1(n637), .A2(n636), .ZN(n639) );
  NOR2_X1 U699 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U700 ( .A(KEYINPUT51), .B(n640), .Z(n641) );
  NOR2_X1 U701 ( .A1(n658), .A2(n641), .ZN(n653) );
  NOR2_X1 U702 ( .A1(n353), .A2(n642), .ZN(n643) );
  XNOR2_X1 U703 ( .A(n643), .B(KEYINPUT118), .ZN(n644) );
  NOR2_X1 U704 ( .A1(n645), .A2(n644), .ZN(n649) );
  NOR2_X1 U705 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U706 ( .A1(n649), .A2(n648), .ZN(n651) );
  INV_X1 U707 ( .A(n659), .ZN(n650) );
  NOR2_X1 U708 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U709 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U710 ( .A(KEYINPUT52), .B(n654), .Z(n655) );
  XNOR2_X1 U711 ( .A(n655), .B(KEYINPUT119), .ZN(n657) );
  NOR2_X1 U712 ( .A1(n657), .A2(n656), .ZN(n663) );
  INV_X1 U713 ( .A(n658), .ZN(n660) );
  NAND2_X1 U714 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U715 ( .A1(n661), .A2(n723), .ZN(n662) );
  NOR2_X1 U716 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U717 ( .A1(n665), .A2(n664), .ZN(n667) );
  XOR2_X1 U718 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n666) );
  XNOR2_X1 U719 ( .A(n667), .B(n666), .ZN(G75) );
  XOR2_X1 U720 ( .A(G101), .B(n668), .Z(G3) );
  NAND2_X1 U721 ( .A1(n670), .A2(n357), .ZN(n669) );
  XNOR2_X1 U722 ( .A(n669), .B(G104), .ZN(G6) );
  XOR2_X1 U723 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n672) );
  NAND2_X1 U724 ( .A1(n670), .A2(n683), .ZN(n671) );
  XNOR2_X1 U725 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U726 ( .A(G107), .B(n673), .ZN(G9) );
  XOR2_X1 U727 ( .A(G110), .B(KEYINPUT115), .Z(n674) );
  XNOR2_X1 U728 ( .A(n675), .B(n674), .ZN(G12) );
  XOR2_X1 U729 ( .A(KEYINPUT116), .B(KEYINPUT29), .Z(n677) );
  NAND2_X1 U730 ( .A1(n680), .A2(n683), .ZN(n676) );
  XNOR2_X1 U731 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U732 ( .A(n359), .B(n678), .ZN(G30) );
  XNOR2_X1 U733 ( .A(G143), .B(n679), .ZN(G45) );
  NAND2_X1 U734 ( .A1(n680), .A2(n357), .ZN(n681) );
  XNOR2_X1 U735 ( .A(n681), .B(G146), .ZN(G48) );
  NAND2_X1 U736 ( .A1(n357), .A2(n684), .ZN(n682) );
  XNOR2_X1 U737 ( .A(G113), .B(n682), .ZN(G15) );
  NAND2_X1 U738 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U739 ( .A(n685), .B(G116), .ZN(G18) );
  XNOR2_X1 U740 ( .A(KEYINPUT37), .B(KEYINPUT117), .ZN(n686) );
  XNOR2_X1 U741 ( .A(n687), .B(n686), .ZN(n688) );
  XNOR2_X1 U742 ( .A(G125), .B(n688), .ZN(G27) );
  XNOR2_X1 U743 ( .A(G134), .B(n689), .ZN(G36) );
  XOR2_X1 U744 ( .A(G140), .B(n690), .Z(G42) );
  NAND2_X1 U745 ( .A1(n697), .A2(G469), .ZN(n695) );
  XNOR2_X1 U746 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n691) );
  XNOR2_X1 U747 ( .A(n691), .B(KEYINPUT57), .ZN(n692) );
  XNOR2_X1 U748 ( .A(n693), .B(n692), .ZN(n694) );
  XNOR2_X1 U749 ( .A(n695), .B(n694), .ZN(n696) );
  NOR2_X1 U750 ( .A1(n701), .A2(n696), .ZN(G54) );
  NAND2_X1 U751 ( .A1(n697), .A2(G478), .ZN(n699) );
  XNOR2_X1 U752 ( .A(n699), .B(n698), .ZN(n700) );
  NOR2_X1 U753 ( .A1(n701), .A2(n700), .ZN(G63) );
  BUF_X1 U754 ( .A(n702), .Z(n703) );
  NOR2_X1 U755 ( .A1(n703), .A2(G953), .ZN(n708) );
  NAND2_X1 U756 ( .A1(G953), .A2(G224), .ZN(n704) );
  XOR2_X1 U757 ( .A(KEYINPUT61), .B(n704), .Z(n705) );
  NOR2_X1 U758 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U759 ( .A1(n708), .A2(n707), .ZN(n715) );
  XOR2_X1 U760 ( .A(KEYINPUT125), .B(KEYINPUT124), .Z(n713) );
  XOR2_X1 U761 ( .A(n709), .B(G101), .Z(n711) );
  NAND2_X1 U762 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U763 ( .A(n713), .B(n712), .ZN(n714) );
  XNOR2_X1 U764 ( .A(n715), .B(n714), .ZN(G69) );
  XNOR2_X1 U765 ( .A(n717), .B(n716), .ZN(n720) );
  XNOR2_X1 U766 ( .A(n720), .B(G227), .ZN(n718) );
  NOR2_X1 U767 ( .A1(n723), .A2(n718), .ZN(n719) );
  NAND2_X1 U768 ( .A1(n719), .A2(G900), .ZN(n726) );
  XNOR2_X1 U769 ( .A(n721), .B(n720), .ZN(n722) );
  XNOR2_X1 U770 ( .A(n722), .B(KEYINPUT126), .ZN(n724) );
  NAND2_X1 U771 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U772 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U773 ( .A(n727), .B(KEYINPUT127), .ZN(G72) );
  XNOR2_X1 U774 ( .A(n728), .B(G119), .ZN(G21) );
  XOR2_X1 U775 ( .A(n729), .B(G131), .Z(G33) );
  XOR2_X1 U776 ( .A(G137), .B(n730), .Z(G39) );
endmodule

