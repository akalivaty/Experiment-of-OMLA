//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 1 1 1 0 1 1 0 0 1 0 0 0 0 1 0 1 1 1 0 1 1 0 1 1 0 0 1 1 0 0 1 1 0 0 0 1 1 0 1 0 1 0 0 1 0 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1283, new_n1284, new_n1285,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(KEYINPUT64), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT64), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G68), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G58), .A2(G232), .ZN(new_n224));
  NAND4_X1  g0024(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n209), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n227), .A2(new_n207), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(new_n201), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n212), .B1(KEYINPUT1), .B2(new_n226), .C1(new_n229), .C2(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT65), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G250), .B(G257), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT66), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n238), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n202), .A2(G68), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n213), .A2(G50), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n246), .B(new_n251), .ZN(G351));
  NOR2_X1   g0052(.A1(new_n207), .A2(G1), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(KEYINPUT70), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n227), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n254), .A2(G50), .A3(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n260), .B1(G50), .B2(new_n255), .ZN(new_n261));
  INV_X1    g0061(.A(new_n258), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT8), .B(G58), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n207), .A2(G33), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G20), .A2(G33), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n264), .A2(new_n266), .B1(G150), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n203), .A2(G20), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n262), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n261), .A2(new_n270), .ZN(new_n271));
  XOR2_X1   g0071(.A(new_n271), .B(KEYINPUT9), .Z(new_n272));
  AND2_X1   g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  OAI21_X1  g0073(.A(G274), .B1(new_n273), .B2(new_n227), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT67), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n276));
  NOR3_X1   g0076(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G274), .ZN(new_n278));
  AND2_X1   g0078(.A1(G1), .A2(G13), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G41), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G41), .ZN(new_n282));
  INV_X1    g0082(.A(G45), .ZN(new_n283));
  AOI21_X1  g0083(.A(G1), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(KEYINPUT67), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n277), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n273), .A2(new_n227), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(new_n284), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n286), .B1(G226), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT69), .ZN(new_n290));
  NOR3_X1   g0090(.A1(new_n273), .A2(new_n290), .A3(new_n227), .ZN(new_n291));
  AOI21_X1  g0091(.A(KEYINPUT69), .B1(new_n279), .B2(new_n280), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G223), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT3), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G33), .ZN(new_n296));
  INV_X1    g0096(.A(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT3), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G1698), .ZN(new_n300));
  OAI21_X1  g0100(.A(KEYINPUT68), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  XNOR2_X1  g0101(.A(KEYINPUT3), .B(G33), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT68), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n302), .A2(new_n303), .A3(G1698), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n294), .B1(new_n301), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n302), .A2(new_n300), .ZN(new_n306));
  INV_X1    g0106(.A(G222), .ZN(new_n307));
  INV_X1    g0107(.A(G77), .ZN(new_n308));
  OAI22_X1  g0108(.A1(new_n306), .A2(new_n307), .B1(new_n308), .B2(new_n302), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n293), .B1(new_n305), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n289), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G200), .ZN(new_n312));
  INV_X1    g0112(.A(G190), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n272), .B(new_n312), .C1(new_n313), .C2(new_n311), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n314), .B(KEYINPUT10), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n311), .A2(G179), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n316), .B(KEYINPUT71), .ZN(new_n317));
  INV_X1    g0117(.A(G169), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n271), .B1(new_n311), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n254), .A2(new_n264), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n322), .A2(new_n259), .B1(new_n256), .B2(new_n263), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n201), .B1(new_n217), .B2(G58), .ZN(new_n325));
  INV_X1    g0125(.A(G159), .ZN(new_n326));
  INV_X1    g0126(.A(new_n267), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n325), .A2(new_n207), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n297), .A2(KEYINPUT3), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n295), .A2(G33), .ZN(new_n330));
  OAI211_X1 g0130(.A(KEYINPUT7), .B(new_n207), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT76), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT7), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n334), .B1(new_n302), .B2(G20), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n299), .A2(KEYINPUT76), .A3(KEYINPUT7), .A4(new_n207), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n333), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n328), .B1(new_n337), .B2(G68), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n262), .B1(new_n338), .B2(KEYINPUT16), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT16), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT77), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n296), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n295), .A2(KEYINPUT77), .A3(G33), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n342), .A2(new_n298), .A3(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n334), .A2(G20), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n218), .B1(new_n346), .B2(new_n335), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n340), .B1(new_n347), .B2(new_n328), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n324), .B1(new_n339), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n279), .A2(new_n280), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n290), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n279), .A2(KEYINPUT69), .A3(new_n280), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(G33), .A2(G87), .ZN(new_n354));
  OR2_X1    g0154(.A1(new_n300), .A2(G226), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n302), .B(new_n355), .C1(G223), .C2(G1698), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n353), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n357), .A2(G179), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n288), .A2(G232), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n277), .B2(new_n285), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT78), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n275), .B1(new_n274), .B2(new_n276), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n281), .A2(KEYINPUT67), .A3(new_n284), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n365), .A2(KEYINPUT78), .A3(new_n359), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n358), .A2(new_n362), .A3(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n318), .B1(new_n360), .B2(new_n357), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(KEYINPUT18), .B1(new_n349), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n356), .A2(new_n354), .ZN(new_n371));
  AOI21_X1  g0171(.A(G190), .B1(new_n371), .B2(new_n293), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n362), .A2(new_n366), .A3(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G200), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n360), .B2(new_n357), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n336), .A2(new_n335), .ZN(new_n377));
  AOI21_X1  g0177(.A(G20), .B1(new_n296), .B2(new_n298), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT76), .B1(new_n378), .B2(KEYINPUT7), .ZN(new_n379));
  OAI21_X1  g0179(.A(G68), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n328), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n380), .A2(new_n381), .A3(KEYINPUT16), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n382), .A2(new_n348), .A3(new_n258), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n376), .A2(new_n383), .A3(new_n323), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT17), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n369), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n383), .A2(new_n323), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT18), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n376), .A2(new_n383), .A3(KEYINPUT17), .A4(new_n323), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n370), .A2(new_n386), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n217), .A2(new_n207), .ZN(new_n393));
  OAI22_X1  g0193(.A1(new_n327), .A2(new_n202), .B1(new_n265), .B2(new_n308), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n258), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  XNOR2_X1  g0195(.A(new_n395), .B(KEYINPUT11), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n255), .A2(KEYINPUT74), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT74), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n398), .A2(new_n206), .A3(G13), .A4(G20), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n400), .A2(KEYINPUT12), .A3(new_n218), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n258), .B1(new_n397), .B2(new_n399), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n254), .A2(new_n402), .A3(G68), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT12), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(new_n255), .B2(G68), .ZN(new_n405));
  AND3_X1   g0205(.A1(new_n401), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n396), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n288), .A2(G238), .ZN(new_n408));
  NOR2_X1   g0208(.A1(G226), .A2(G1698), .ZN(new_n409));
  INV_X1    g0209(.A(G232), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n409), .B1(new_n410), .B2(G1698), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n411), .A2(new_n302), .B1(G33), .B2(G97), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n408), .B1(new_n412), .B2(new_n353), .ZN(new_n413));
  OAI21_X1  g0213(.A(KEYINPUT13), .B1(new_n413), .B2(new_n286), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G33), .A2(G97), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n410), .A2(G1698), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n416), .B1(G226), .B2(G1698), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n415), .B1(new_n417), .B2(new_n299), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n418), .A2(new_n293), .B1(new_n288), .B2(G238), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT13), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(new_n420), .A3(new_n365), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n414), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT14), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n422), .A2(new_n423), .A3(G169), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n414), .A2(G179), .A3(new_n421), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n423), .B1(new_n422), .B2(G169), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n407), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NOR3_X1   g0228(.A1(new_n413), .A2(new_n286), .A3(KEYINPUT13), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n420), .B1(new_n419), .B2(new_n365), .ZN(new_n430));
  OAI21_X1  g0230(.A(G200), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n431), .A2(new_n396), .A3(new_n406), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT75), .B1(new_n422), .B2(new_n313), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT75), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n414), .A2(new_n435), .A3(new_n421), .A4(G190), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  XNOR2_X1  g0238(.A(KEYINPUT15), .B(G87), .ZN(new_n439));
  OR3_X1    g0239(.A1(new_n439), .A2(KEYINPUT73), .A3(new_n265), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT73), .B1(new_n439), .B2(new_n265), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n264), .A2(new_n267), .B1(G20), .B2(G77), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT72), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n440), .B(new_n441), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  AND2_X1   g0244(.A1(new_n442), .A2(new_n443), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n258), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n254), .A2(G77), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n447), .A2(new_n402), .B1(new_n308), .B2(new_n400), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n286), .B1(G244), .B2(new_n288), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n219), .B1(new_n301), .B2(new_n304), .ZN(new_n450));
  INV_X1    g0250(.A(G107), .ZN(new_n451));
  OAI22_X1  g0251(.A1(new_n306), .A2(new_n410), .B1(new_n451), .B2(new_n302), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n293), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n446), .B(new_n448), .C1(new_n454), .C2(new_n313), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n374), .B1(new_n449), .B2(new_n453), .ZN(new_n456));
  OR2_X1    g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n454), .A2(new_n318), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n446), .A2(new_n448), .ZN(new_n459));
  INV_X1    g0259(.A(G179), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n449), .A2(new_n460), .A3(new_n453), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n458), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n428), .A2(new_n438), .A3(new_n457), .A4(new_n462), .ZN(new_n463));
  NOR3_X1   g0263(.A1(new_n321), .A2(new_n392), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n451), .B1(new_n346), .B2(new_n335), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT6), .ZN(new_n466));
  INV_X1    g0266(.A(G97), .ZN(new_n467));
  NOR3_X1   g0267(.A1(new_n466), .A2(new_n467), .A3(G107), .ZN(new_n468));
  XNOR2_X1  g0268(.A(G97), .B(G107), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n468), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  OAI22_X1  g0270(.A1(new_n470), .A2(new_n207), .B1(new_n308), .B2(new_n327), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n258), .B1(new_n465), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n259), .B1(G1), .B2(new_n297), .ZN(new_n473));
  MUX2_X1   g0273(.A(new_n255), .B(new_n473), .S(G97), .Z(new_n474));
  NAND2_X1  g0274(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n296), .A2(new_n298), .A3(G244), .A4(new_n300), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT4), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT79), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n302), .A2(KEYINPUT4), .A3(G244), .A4(new_n300), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT80), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n477), .A2(KEYINPUT79), .A3(new_n478), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n481), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n296), .A2(new_n298), .A3(G250), .A4(G1698), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G283), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n487), .B(new_n488), .C1(new_n482), .C2(new_n483), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n293), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n283), .A2(G1), .ZN(new_n491));
  AND2_X1   g0291(.A1(KEYINPUT5), .A2(G41), .ZN(new_n492));
  NOR2_X1   g0292(.A1(KEYINPUT5), .A2(G41), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n494), .A2(new_n274), .ZN(new_n495));
  XNOR2_X1  g0295(.A(KEYINPUT5), .B(G41), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n287), .B1(new_n491), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n495), .B1(G257), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n490), .A2(G190), .A3(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n498), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n487), .A2(new_n488), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n477), .A2(new_n478), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n501), .B1(new_n502), .B2(KEYINPUT80), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n503), .A2(new_n484), .A3(new_n481), .A4(new_n485), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n500), .B1(new_n504), .B2(new_n293), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n476), .B(new_n499), .C1(new_n374), .C2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n490), .A2(new_n460), .A3(new_n498), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n507), .B(new_n475), .C1(new_n505), .C2(G169), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n302), .A2(new_n207), .A3(G87), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT22), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT22), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n302), .A2(new_n511), .A3(new_n207), .A4(G87), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT24), .ZN(new_n514));
  INV_X1    g0314(.A(G116), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(KEYINPUT81), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT81), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G116), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n297), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT23), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n520), .B1(new_n207), .B2(G107), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n451), .A2(KEYINPUT23), .A3(G20), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n519), .A2(new_n207), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n513), .A2(new_n514), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n514), .B1(new_n513), .B2(new_n523), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n258), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n473), .A2(new_n451), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT25), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(new_n255), .B2(G107), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n256), .A2(KEYINPUT25), .A3(new_n451), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n527), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n296), .A2(new_n298), .A3(G257), .A4(G1698), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n296), .A2(new_n298), .A3(G250), .A4(new_n300), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G33), .A2(G294), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n293), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n497), .A2(G264), .ZN(new_n537));
  INV_X1    g0337(.A(new_n495), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(G190), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n293), .A2(new_n535), .B1(new_n497), .B2(G264), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n538), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(G200), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n526), .A2(new_n531), .A3(new_n540), .A4(new_n543), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n506), .A2(new_n508), .A3(new_n544), .ZN(new_n545));
  XNOR2_X1  g0345(.A(KEYINPUT81), .B(G116), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n397), .A2(new_n546), .A3(new_n399), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT87), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n397), .A2(new_n546), .A3(KEYINPUT87), .A4(new_n399), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n515), .B1(new_n206), .B2(G33), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n549), .A2(new_n550), .B1(new_n402), .B2(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n488), .B(new_n207), .C1(G33), .C2(new_n467), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT88), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n297), .A2(G97), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT88), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n555), .A2(new_n556), .A3(new_n207), .A4(new_n488), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n546), .A2(G20), .B1(new_n227), .B2(new_n257), .ZN(new_n559));
  AND3_X1   g0359(.A1(new_n558), .A2(KEYINPUT20), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(KEYINPUT20), .B1(new_n558), .B2(new_n559), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n552), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n296), .A2(new_n298), .A3(G264), .A4(G1698), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n296), .A2(new_n298), .A3(G257), .A4(new_n300), .ZN(new_n564));
  INV_X1    g0364(.A(G303), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n563), .B(new_n564), .C1(new_n565), .C2(new_n302), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n293), .ZN(new_n567));
  AOI21_X1  g0367(.A(KEYINPUT86), .B1(new_n497), .B2(G270), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n494), .A2(KEYINPUT86), .A3(G270), .A4(new_n350), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n538), .B(new_n567), .C1(new_n568), .C2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n562), .A2(G169), .A3(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(KEYINPUT89), .A2(KEYINPUT21), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT86), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n494), .A2(new_n350), .ZN(new_n576));
  INV_X1    g0376(.A(G270), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n569), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n579), .A2(G179), .A3(new_n538), .A4(new_n567), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n562), .ZN(new_n582));
  INV_X1    g0382(.A(new_n573), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n562), .A2(new_n571), .A3(G169), .A4(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n574), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n318), .B1(new_n541), .B2(new_n538), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n586), .A2(KEYINPUT90), .B1(new_n539), .B2(G179), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT90), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(new_n539), .B2(new_n318), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n587), .A2(new_n589), .B1(new_n526), .B2(new_n531), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n585), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n517), .A2(G116), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n515), .A2(KEYINPUT81), .ZN(new_n593));
  OAI21_X1  g0393(.A(G33), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n219), .A2(new_n300), .ZN(new_n595));
  INV_X1    g0395(.A(G244), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(G1698), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n296), .A2(new_n595), .A3(new_n298), .A4(new_n597), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n594), .A2(new_n598), .A3(KEYINPUT82), .ZN(new_n599));
  AOI21_X1  g0399(.A(KEYINPUT82), .B1(new_n594), .B2(new_n598), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n293), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n206), .A2(G45), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n602), .A2(G250), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n350), .A2(new_n603), .B1(new_n281), .B2(new_n491), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT19), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n207), .B1(new_n415), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(G87), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n608), .A2(new_n467), .A3(new_n451), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n296), .A2(new_n298), .A3(new_n207), .A4(G68), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n606), .B1(new_n265), .B2(new_n467), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n258), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n400), .A2(new_n439), .ZN(new_n615));
  INV_X1    g0415(.A(new_n439), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n259), .B(new_n616), .C1(G1), .C2(new_n297), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n614), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT84), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n605), .A2(new_n318), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n601), .A2(new_n460), .A3(new_n604), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT83), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n614), .A2(new_n617), .A3(new_n615), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(KEYINPUT84), .ZN(new_n625));
  INV_X1    g0425(.A(new_n604), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT82), .ZN(new_n627));
  AND4_X1   g0427(.A1(new_n296), .A2(new_n595), .A3(new_n298), .A4(new_n597), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n627), .B1(new_n628), .B2(new_n519), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n594), .A2(new_n598), .A3(KEYINPUT82), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n626), .B1(new_n631), .B2(new_n293), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n632), .A2(KEYINPUT83), .A3(new_n460), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n620), .A2(new_n623), .A3(new_n625), .A4(new_n633), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n614), .B(new_n615), .C1(new_n608), .C2(new_n473), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n635), .B1(new_n605), .B2(G200), .ZN(new_n636));
  AOI21_X1  g0436(.A(KEYINPUT85), .B1(new_n632), .B2(G190), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n353), .B1(new_n629), .B2(new_n630), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT85), .ZN(new_n639));
  NOR4_X1   g0439(.A1(new_n638), .A2(new_n639), .A3(new_n313), .A4(new_n626), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n636), .B1(new_n637), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n562), .B1(G200), .B2(new_n571), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n579), .A2(G190), .A3(new_n538), .A4(new_n567), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n634), .A2(new_n641), .A3(new_n644), .ZN(new_n645));
  AND4_X1   g0445(.A1(new_n464), .A2(new_n545), .A3(new_n591), .A4(new_n645), .ZN(new_n646));
  XNOR2_X1  g0446(.A(new_n646), .B(KEYINPUT91), .ZN(G372));
  INV_X1    g0447(.A(KEYINPUT92), .ZN(new_n648));
  OAI21_X1  g0448(.A(G200), .B1(new_n638), .B2(new_n626), .ZN(new_n649));
  INV_X1    g0449(.A(new_n635), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n639), .B1(new_n605), .B2(new_n313), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n632), .A2(KEYINPUT85), .A3(G190), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n618), .A2(new_n619), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n318), .B1(new_n638), .B2(new_n626), .ZN(new_n656));
  AND4_X1   g0456(.A1(new_n625), .A2(new_n655), .A3(new_n656), .A4(new_n621), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n648), .B1(new_n654), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n620), .A2(new_n625), .A3(new_n621), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n641), .A2(new_n659), .A3(KEYINPUT92), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT93), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n508), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n490), .A2(new_n498), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n318), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n665), .A2(KEYINPUT93), .A3(new_n475), .A4(new_n507), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT26), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n661), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n587), .A2(new_n589), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n526), .A2(new_n531), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n672), .A2(new_n574), .A3(new_n582), .A4(new_n584), .ZN(new_n673));
  INV_X1    g0473(.A(new_n660), .ZN(new_n674));
  AOI21_X1  g0474(.A(KEYINPUT92), .B1(new_n641), .B2(new_n659), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n673), .B(new_n545), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n508), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n677), .A2(new_n641), .A3(new_n634), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n657), .B1(new_n678), .B2(KEYINPUT26), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n669), .A2(new_n676), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n464), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n370), .A2(new_n390), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n462), .ZN(new_n684));
  INV_X1    g0484(.A(new_n427), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n685), .A2(new_n425), .A3(new_n424), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n438), .A2(new_n684), .B1(new_n686), .B2(new_n407), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n386), .A2(new_n391), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n683), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  AOI22_X1  g0489(.A1(new_n689), .A2(new_n315), .B1(new_n317), .B2(new_n319), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n681), .A2(new_n690), .ZN(G369));
  NAND3_X1  g0491(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n692));
  OR2_X1    g0492(.A1(new_n692), .A2(KEYINPUT27), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(KEYINPUT27), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n693), .A2(G213), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G343), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT94), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n671), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n590), .B1(new_n544), .B2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n698), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n590), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n698), .A2(new_n562), .ZN(new_n705));
  XOR2_X1   g0505(.A(new_n585), .B(new_n705), .Z(new_n706));
  NAND3_X1  g0506(.A1(new_n706), .A2(KEYINPUT95), .A3(new_n644), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(KEYINPUT95), .B1(new_n706), .B2(new_n644), .ZN(new_n709));
  OAI211_X1 g0509(.A(G330), .B(new_n704), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n699), .A2(new_n544), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n672), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n585), .A2(new_n701), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n703), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n710), .A2(new_n714), .ZN(G399));
  INV_X1    g0515(.A(new_n210), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(G41), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n609), .A2(G116), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(G1), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(new_n231), .B2(new_n718), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT28), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT99), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n668), .B1(new_n661), .B2(new_n667), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n677), .A2(new_n668), .A3(new_n641), .A4(new_n634), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n659), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n723), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  AND2_X1   g0527(.A1(new_n725), .A2(new_n659), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n663), .A2(new_n666), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n729), .B1(new_n658), .B2(new_n660), .ZN(new_n730));
  OAI211_X1 g0530(.A(new_n728), .B(KEYINPUT99), .C1(new_n730), .C2(new_n668), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n727), .A2(new_n676), .A3(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n732), .A2(KEYINPUT29), .A3(new_n701), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT98), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n680), .A2(new_n701), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT29), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AOI211_X1 g0537(.A(KEYINPUT98), .B(KEYINPUT29), .C1(new_n680), .C2(new_n701), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n733), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(KEYINPUT96), .A2(KEYINPUT30), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n536), .A2(new_n537), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n638), .A2(new_n742), .A3(new_n626), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n505), .A2(new_n581), .A3(new_n741), .A4(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(G179), .B1(new_n601), .B2(new_n604), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n664), .A2(new_n542), .A3(new_n571), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n580), .A2(new_n605), .A3(new_n742), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n741), .B1(new_n748), .B2(new_n505), .ZN(new_n749));
  OAI211_X1 g0549(.A(KEYINPUT31), .B(new_n698), .C1(new_n747), .C2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n581), .A2(new_n743), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n740), .B1(new_n752), .B2(new_n664), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n753), .A2(new_n746), .A3(new_n744), .ZN(new_n754));
  AOI21_X1  g0554(.A(KEYINPUT31), .B1(new_n754), .B2(new_n698), .ZN(new_n755));
  OAI21_X1  g0555(.A(KEYINPUT97), .B1(new_n751), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n698), .B1(new_n747), .B2(new_n749), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT31), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT97), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n759), .A2(new_n760), .A3(new_n750), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n545), .A2(new_n645), .A3(new_n591), .A4(new_n701), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n756), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G330), .ZN(new_n764));
  AND2_X1   g0564(.A1(new_n739), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n722), .B1(new_n765), .B2(G1), .ZN(G364));
  OAI21_X1  g0566(.A(G330), .B1(new_n708), .B2(new_n709), .ZN(new_n767));
  INV_X1    g0567(.A(new_n709), .ZN(new_n768));
  INV_X1    g0568(.A(G330), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n768), .A2(new_n769), .A3(new_n707), .ZN(new_n770));
  INV_X1    g0570(.A(G13), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n206), .B1(new_n772), .B2(G45), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n717), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AND3_X1   g0576(.A1(new_n767), .A2(new_n770), .A3(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n207), .A2(G179), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n778), .A2(G190), .A3(G200), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n608), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n207), .A2(new_n460), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G200), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n313), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT32), .ZN(new_n785));
  NOR2_X1   g0585(.A1(G190), .A2(G200), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n778), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n326), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n784), .A2(new_n202), .B1(new_n785), .B2(new_n788), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n780), .B(new_n789), .C1(new_n785), .C2(new_n788), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n781), .A2(G190), .A3(new_n374), .ZN(new_n791));
  INV_X1    g0591(.A(G58), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n302), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n313), .A2(G179), .A3(G200), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n207), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n778), .A2(new_n313), .A3(G200), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n795), .A2(new_n467), .B1(new_n796), .B2(new_n451), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n782), .A2(G190), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n793), .B(new_n797), .C1(G68), .C2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n781), .A2(new_n786), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AND2_X1   g0601(.A1(new_n801), .A2(KEYINPUT101), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n801), .A2(KEYINPUT101), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n790), .B(new_n799), .C1(new_n308), .C2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(G317), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(KEYINPUT33), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n806), .A2(KEYINPUT33), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n798), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(G294), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n809), .B1(new_n810), .B2(new_n795), .C1(new_n565), .C2(new_n779), .ZN(new_n811));
  INV_X1    g0611(.A(new_n787), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n302), .B1(new_n812), .B2(G329), .ZN(new_n813));
  INV_X1    g0613(.A(G311), .ZN(new_n814));
  INV_X1    g0614(.A(G322), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n813), .B1(new_n814), .B2(new_n800), .C1(new_n815), .C2(new_n791), .ZN(new_n816));
  INV_X1    g0616(.A(G326), .ZN(new_n817));
  INV_X1    g0617(.A(G283), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n784), .A2(new_n817), .B1(new_n796), .B2(new_n818), .ZN(new_n819));
  NOR3_X1   g0619(.A1(new_n811), .A2(new_n816), .A3(new_n819), .ZN(new_n820));
  OR2_X1    g0620(.A1(new_n820), .A2(KEYINPUT102), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(KEYINPUT102), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n805), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n227), .B1(G20), .B2(new_n318), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n716), .A2(new_n299), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n826), .A2(G355), .B1(new_n515), .B2(new_n716), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n210), .A2(new_n299), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT100), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(G45), .B2(new_n231), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n251), .A2(new_n283), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n827), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(G13), .A2(G33), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n834), .A2(G20), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(new_n824), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n776), .B1(new_n832), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n825), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n706), .A2(new_n644), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n838), .B1(new_n839), .B2(new_n835), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n777), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(G396));
  NAND2_X1  g0642(.A1(new_n459), .A2(new_n698), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n455), .B2(new_n456), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n462), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n684), .A2(new_n701), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n735), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n847), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n680), .A2(new_n701), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  OR2_X1    g0651(.A1(new_n851), .A2(new_n764), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n775), .B1(new_n851), .B2(new_n764), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n824), .A2(new_n833), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n608), .A2(new_n796), .B1(new_n779), .B2(new_n451), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n299), .B1(new_n787), .B2(new_n814), .ZN(new_n858));
  INV_X1    g0658(.A(new_n791), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n858), .B1(G294), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n795), .ZN(new_n861));
  AOI22_X1  g0661(.A1(G97), .A2(new_n861), .B1(new_n783), .B2(G303), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n860), .B(new_n862), .C1(new_n804), .C2(new_n546), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n857), .B(new_n863), .C1(G283), .C2(new_n798), .ZN(new_n864));
  INV_X1    g0664(.A(G132), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n302), .B1(new_n787), .B2(new_n865), .C1(new_n202), .C2(new_n779), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n795), .A2(new_n792), .B1(new_n796), .B2(new_n213), .ZN(new_n867));
  AOI22_X1  g0667(.A1(G137), .A2(new_n783), .B1(new_n859), .B2(G143), .ZN(new_n868));
  INV_X1    g0668(.A(G150), .ZN(new_n869));
  INV_X1    g0669(.A(new_n798), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n804), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n871), .B1(G159), .B2(new_n872), .ZN(new_n873));
  XOR2_X1   g0673(.A(KEYINPUT103), .B(KEYINPUT34), .Z(new_n874));
  AOI211_X1 g0674(.A(new_n866), .B(new_n867), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  OR2_X1    g0675(.A1(new_n873), .A2(new_n874), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n864), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n824), .ZN(new_n878));
  OAI221_X1 g0678(.A(new_n775), .B1(G77), .B2(new_n856), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(new_n833), .B2(new_n847), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n880), .B(KEYINPUT104), .Z(new_n881));
  NOR2_X1   g0681(.A1(new_n854), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(G384));
  INV_X1    g0683(.A(new_n470), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n515), .B(new_n229), .C1(new_n884), .C2(KEYINPUT35), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(KEYINPUT35), .B2(new_n884), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n886), .B(KEYINPUT36), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n308), .B(new_n231), .C1(new_n217), .C2(G58), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n888), .A2(KEYINPUT105), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n888), .A2(KEYINPUT105), .ZN(new_n890));
  XOR2_X1   g0690(.A(new_n247), .B(KEYINPUT106), .Z(new_n891));
  NOR3_X1   g0691(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n771), .A2(G1), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n733), .B(new_n464), .C1(new_n737), .C2(new_n738), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n690), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n850), .A2(new_n846), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n380), .A2(new_n381), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n340), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n324), .B1(new_n339), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n695), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n384), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n899), .A2(new_n369), .ZN(new_n902));
  OAI21_X1  g0702(.A(KEYINPUT37), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n387), .A2(new_n388), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n388), .A2(new_n695), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT37), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n904), .A2(new_n905), .A3(new_n906), .A4(new_n384), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n899), .A2(new_n900), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n392), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT38), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n908), .A2(new_n910), .A3(KEYINPUT38), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n432), .B1(new_n436), .B2(new_n434), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n407), .B(new_n698), .C1(new_n916), .C2(new_n686), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n698), .A2(new_n407), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n428), .A2(new_n438), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n896), .A2(new_n915), .A3(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n683), .A2(new_n695), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT39), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n908), .A2(new_n910), .A3(KEYINPUT38), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n904), .A2(new_n905), .A3(new_n384), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(KEYINPUT37), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n907), .ZN(new_n928));
  INV_X1    g0728(.A(new_n905), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n392), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT38), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n924), .B1(new_n925), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n913), .A2(KEYINPUT39), .A3(new_n914), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n686), .A2(new_n407), .A3(new_n701), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n932), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n921), .A2(new_n923), .A3(new_n936), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n895), .B(new_n937), .Z(new_n938));
  INV_X1    g0738(.A(KEYINPUT107), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n925), .A2(new_n931), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n762), .A2(new_n759), .A3(new_n750), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n847), .B1(new_n917), .B2(new_n919), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n941), .A2(new_n942), .A3(KEYINPUT40), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n939), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  AND3_X1   g0744(.A1(new_n941), .A2(new_n942), .A3(KEYINPUT40), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n907), .A2(new_n927), .B1(new_n392), .B2(new_n929), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n914), .B1(new_n946), .B2(KEYINPUT38), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n945), .A2(KEYINPUT107), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(KEYINPUT38), .B1(new_n908), .B2(new_n910), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n941), .B(new_n942), .C1(new_n925), .C2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT40), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n944), .A2(new_n948), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n464), .A2(new_n941), .ZN(new_n954));
  OAI21_X1  g0754(.A(G330), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n954), .B2(new_n953), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n938), .A2(new_n956), .B1(new_n206), .B2(new_n772), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n938), .A2(new_n956), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n887), .B1(new_n892), .B2(new_n893), .C1(new_n957), .C2(new_n958), .ZN(G367));
  OAI211_X1 g0759(.A(new_n506), .B(new_n508), .C1(new_n476), .C2(new_n701), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n677), .A2(new_n698), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT109), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n960), .A2(new_n961), .A3(KEYINPUT109), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n712), .A2(new_n702), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n585), .A2(new_n701), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(KEYINPUT110), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT110), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n966), .A2(new_n972), .A3(new_n969), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(KEYINPUT42), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT42), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n971), .A2(new_n976), .A3(new_n973), .ZN(new_n977));
  AND3_X1   g0777(.A1(new_n960), .A2(new_n961), .A3(KEYINPUT109), .ZN(new_n978));
  AOI21_X1  g0778(.A(KEYINPUT109), .B1(new_n960), .B2(new_n961), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n508), .B1(new_n980), .B2(new_n672), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n701), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n975), .A2(new_n977), .A3(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n701), .A2(new_n650), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(new_n658), .B2(new_n660), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(new_n657), .B2(new_n984), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT43), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n983), .A2(new_n988), .ZN(new_n989));
  OR3_X1    g0789(.A1(new_n710), .A2(KEYINPUT111), .A3(new_n980), .ZN(new_n990));
  OAI21_X1  g0790(.A(KEYINPUT111), .B1(new_n710), .B2(new_n980), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n986), .A2(new_n987), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT108), .Z(new_n995));
  NAND4_X1  g0795(.A1(new_n983), .A2(new_n988), .A3(new_n991), .A4(new_n990), .ZN(new_n996));
  AND3_X1   g0796(.A1(new_n993), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n995), .B1(new_n993), .B2(new_n996), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT114), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n969), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(KEYINPUT114), .B1(new_n967), .B2(new_n968), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT113), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n967), .A2(new_n1003), .A3(new_n968), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1003), .B1(new_n967), .B2(new_n968), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1001), .B(new_n1002), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n769), .B1(new_n768), .B2(new_n707), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT115), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1007), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AND2_X1   g0810(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n767), .A2(new_n1011), .A3(new_n1012), .A4(KEYINPUT115), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1014), .A2(new_n739), .A3(new_n764), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT45), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT112), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(new_n966), .B2(new_n714), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n714), .B(new_n1017), .C1(new_n978), .C2(new_n979), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1016), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n702), .B1(new_n700), .B2(new_n968), .ZN(new_n1022));
  OAI21_X1  g0822(.A(KEYINPUT112), .B1(new_n980), .B2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1023), .A2(KEYINPUT45), .A3(new_n1019), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n964), .A2(new_n1022), .A3(new_n965), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT44), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1025), .B(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1021), .A2(new_n1024), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n710), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1021), .A2(new_n1027), .A3(new_n1024), .A4(new_n710), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n765), .B1(new_n1015), .B2(new_n1032), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n717), .B(KEYINPUT41), .Z(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n773), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n999), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n829), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1039), .A2(new_n242), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n836), .B1(new_n210), .B2(new_n439), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n775), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n299), .B1(new_n787), .B2(new_n806), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n784), .A2(new_n814), .B1(new_n451), .B2(new_n795), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1043), .B(new_n1044), .C1(G303), .C2(new_n859), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n779), .A2(new_n546), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1045), .B1(KEYINPUT46), .B2(new_n1046), .C1(new_n818), .C2(new_n804), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n779), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1048), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(new_n467), .B2(new_n796), .C1(new_n870), .C2(new_n810), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n795), .A2(new_n213), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(G58), .B2(new_n1048), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n308), .B2(new_n796), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n302), .B1(new_n791), .B2(new_n869), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G137), .B2(new_n812), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(G143), .A2(new_n783), .B1(new_n798), .B2(G159), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1055), .B(new_n1056), .C1(new_n804), .C2(new_n202), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n1047), .A2(new_n1050), .B1(new_n1053), .B2(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT47), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1042), .B1(new_n1059), .B2(new_n824), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n986), .A2(new_n835), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1038), .A2(new_n1063), .ZN(G387));
  INV_X1    g0864(.A(new_n719), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n826), .A2(new_n1065), .B1(new_n451), .B2(new_n716), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n238), .A2(new_n283), .ZN(new_n1067));
  AOI21_X1  g0867(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1068));
  AND3_X1   g0868(.A1(new_n264), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n1069));
  AOI21_X1  g0869(.A(KEYINPUT50), .B1(new_n264), .B2(new_n202), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n719), .B(new_n1068), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n829), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1066), .B1(new_n1067), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n776), .B1(new_n1073), .B2(new_n836), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n616), .A2(new_n861), .B1(new_n798), .B2(new_n264), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n308), .B2(new_n779), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(G68), .A2(new_n801), .B1(new_n812), .B2(G150), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1077), .B(new_n302), .C1(new_n202), .C2(new_n791), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n784), .A2(new_n326), .B1(new_n796), .B2(new_n467), .ZN(new_n1079));
  NOR3_X1   g0879(.A1(new_n1076), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(G311), .A2(new_n798), .B1(new_n859), .B2(G317), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1081), .B1(new_n815), .B2(new_n784), .C1(new_n804), .C2(new_n565), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT48), .ZN(new_n1083));
  OR2_X1    g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n861), .A2(G283), .B1(new_n1048), .B2(G294), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n1088), .A2(KEYINPUT49), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n299), .B1(new_n787), .B2(new_n817), .C1(new_n546), .C2(new_n796), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n1088), .B2(KEYINPUT49), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1080), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1074), .B1(new_n1092), .B2(new_n878), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n967), .B2(new_n835), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(new_n1014), .B2(new_n774), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n765), .A2(new_n1014), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1015), .A2(new_n717), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1095), .B1(new_n1096), .B2(new_n1097), .ZN(G393));
  NAND3_X1  g0898(.A1(new_n1030), .A2(new_n774), .A3(new_n1031), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT116), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n980), .A2(new_n835), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G317), .A2(new_n783), .B1(new_n859), .B2(G311), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT52), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n299), .B1(new_n787), .B2(new_n815), .C1(new_n810), .C2(new_n800), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n870), .A2(new_n565), .B1(new_n796), .B2(new_n451), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n795), .A2(new_n546), .B1(new_n779), .B2(new_n818), .ZN(new_n1106));
  NOR4_X1   g0906(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n784), .A2(new_n869), .B1(new_n326), .B2(new_n791), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT51), .Z(new_n1109));
  NOR2_X1   g0909(.A1(new_n795), .A2(new_n308), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(G50), .B2(new_n798), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n218), .B2(new_n779), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n299), .B1(new_n812), .B2(G143), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1113), .B1(new_n608), .B2(new_n796), .C1(new_n804), .C2(new_n263), .ZN(new_n1114));
  NOR3_X1   g0914(.A1(new_n1109), .A2(new_n1112), .A3(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n824), .B1(new_n1107), .B2(new_n1115), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n836), .B1(new_n467), .B2(new_n210), .C1(new_n1039), .C2(new_n246), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1101), .A2(new_n775), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  AND3_X1   g0918(.A1(new_n1099), .A2(new_n1100), .A3(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1100), .B1(new_n1099), .B2(new_n1118), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n717), .B1(new_n1015), .B2(new_n1032), .ZN(new_n1121));
  AND2_X1   g0921(.A1(new_n1015), .A2(new_n1032), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n1119), .A2(new_n1120), .B1(new_n1121), .B2(new_n1122), .ZN(G390));
  NAND2_X1  g0923(.A1(new_n932), .A2(new_n933), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n833), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n775), .B1(new_n264), .B2(new_n856), .ZN(new_n1126));
  INV_X1    g0926(.A(G125), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n302), .B1(new_n787), .B2(new_n1127), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n795), .A2(new_n326), .B1(new_n796), .B2(new_n202), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n1128), .B(new_n1129), .C1(G137), .C2(new_n798), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n779), .A2(new_n869), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT53), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(KEYINPUT54), .B(G143), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1130), .B(new_n1132), .C1(new_n804), .C2(new_n1133), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(G128), .A2(new_n783), .B1(new_n859), .B2(G132), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT119), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1110), .B1(G107), .B2(new_n798), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1137), .B1(new_n818), .B2(new_n784), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n299), .B1(new_n791), .B2(new_n515), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(G294), .B2(new_n812), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n796), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n780), .B1(G68), .B2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1140), .B(new_n1142), .C1(new_n804), .C2(new_n467), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n1134), .A2(new_n1136), .B1(new_n1138), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT120), .ZN(new_n1145));
  OR2_X1    g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n878), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1126), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1125), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n920), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n850), .B2(new_n846), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1124), .B1(new_n1152), .B2(new_n935), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n732), .A2(new_n701), .A3(new_n845), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1151), .B1(new_n1154), .B2(new_n846), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n947), .A2(new_n934), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1153), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n941), .A2(G330), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n942), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1157), .A2(new_n1161), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n763), .A2(G330), .A3(new_n849), .A4(new_n920), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1153), .B(new_n1163), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1150), .B1(new_n1165), .B2(new_n774), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT118), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n464), .A2(new_n1159), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n894), .A2(new_n690), .A3(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n763), .A2(G330), .A3(new_n849), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(new_n1151), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n1160), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n896), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n941), .A2(KEYINPUT117), .A3(G330), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(new_n849), .ZN(new_n1176));
  AOI21_X1  g0976(.A(KEYINPUT117), .B1(new_n941), .B2(G330), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1151), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1178), .A2(new_n846), .A3(new_n1154), .A4(new_n1163), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1174), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1168), .B1(new_n1170), .B2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n717), .B1(new_n1167), .B2(new_n1181), .ZN(new_n1182));
  AND2_X1   g0982(.A1(new_n1167), .A2(new_n1181), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1166), .B1(new_n1182), .B2(new_n1183), .ZN(G378));
  NAND3_X1  g0984(.A1(new_n1162), .A2(new_n1164), .A3(new_n1180), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1185), .A2(new_n1170), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n950), .A2(new_n951), .ZN(new_n1187));
  NOR3_X1   g0987(.A1(new_n940), .A2(new_n939), .A3(new_n943), .ZN(new_n1188));
  AOI21_X1  g0988(.A(KEYINPUT107), .B1(new_n945), .B2(new_n947), .ZN(new_n1189));
  OAI211_X1 g0989(.A(G330), .B(new_n1187), .C1(new_n1188), .C2(new_n1189), .ZN(new_n1190));
  AND2_X1   g0990(.A1(new_n936), .A2(new_n923), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1190), .A2(new_n921), .A3(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n271), .A2(new_n900), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n321), .B(new_n1193), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1194), .B(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n937), .A2(new_n952), .A3(G330), .ZN(new_n1197));
  AND3_X1   g0997(.A1(new_n1192), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1196), .B1(new_n1192), .B2(new_n1197), .ZN(new_n1199));
  OAI21_X1  g0999(.A(KEYINPUT57), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n717), .B1(new_n1186), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1192), .A2(new_n1197), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1196), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1192), .A2(new_n1197), .A3(new_n1196), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1185), .A2(new_n1170), .ZN(new_n1207));
  AOI21_X1  g1007(.A(KEYINPUT57), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n1201), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1196), .A2(new_n833), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n775), .B1(G50), .B2(new_n856), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n302), .A2(G41), .ZN(new_n1212));
  AOI211_X1 g1012(.A(G50), .B(new_n1212), .C1(new_n297), .C2(new_n282), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n796), .A2(new_n792), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n784), .A2(new_n515), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1214), .B(new_n1215), .C1(G97), .C2(new_n798), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1212), .B1(new_n818), .B2(new_n787), .C1(new_n439), .C2(new_n800), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1051), .B(new_n1217), .C1(G77), .C2(new_n1048), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n859), .A2(G107), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1219), .B(KEYINPUT121), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1216), .A2(new_n1218), .A3(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT58), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1213), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(KEYINPUT122), .B(G124), .ZN(new_n1224));
  AOI211_X1 g1024(.A(G33), .B(G41), .C1(new_n812), .C2(new_n1224), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n1127), .A2(new_n784), .B1(new_n870), .B2(new_n865), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n859), .A2(G128), .B1(new_n801), .B2(G137), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n779), .B2(new_n1133), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1226), .B(new_n1228), .C1(G150), .C2(new_n861), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT59), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1225), .B1(new_n326), .B2(new_n796), .C1(new_n1229), .C2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1229), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1232), .A2(KEYINPUT59), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1223), .B1(new_n1222), .B2(new_n1221), .C1(new_n1231), .C2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1211), .B1(new_n1234), .B2(new_n824), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n1206), .A2(new_n774), .B1(new_n1210), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1209), .A2(new_n1236), .ZN(G375));
  INV_X1    g1037(.A(KEYINPUT123), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n1170), .B2(new_n1180), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n850), .A2(new_n846), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(new_n1172), .B2(new_n1160), .ZN(new_n1241));
  AND2_X1   g1041(.A1(new_n1178), .A2(new_n1163), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1154), .A2(new_n846), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1241), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n894), .A2(new_n690), .A3(new_n1169), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1244), .A2(KEYINPUT123), .A3(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1170), .A2(new_n1180), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1239), .A2(new_n1246), .A3(new_n1035), .A4(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n859), .A2(G137), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n1249), .B1(new_n870), .B2(new_n1133), .C1(new_n865), .C2(new_n784), .ZN(new_n1250));
  OR2_X1    g1050(.A1(new_n1250), .A2(KEYINPUT124), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(KEYINPUT124), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n800), .A2(new_n869), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n299), .B(new_n1253), .C1(G128), .C2(new_n812), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n779), .A2(new_n326), .ZN(new_n1255));
  AOI211_X1 g1055(.A(new_n1214), .B(new_n1255), .C1(G50), .C2(new_n861), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1251), .A2(new_n1252), .A3(new_n1254), .A4(new_n1256), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n870), .A2(new_n546), .B1(new_n467), .B2(new_n779), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(G294), .B2(new_n783), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n872), .A2(G107), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n299), .B1(new_n787), .B2(new_n565), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1261), .B1(G283), .B2(new_n859), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n861), .A2(new_n616), .B1(new_n1141), .B2(G77), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1259), .A2(new_n1260), .A3(new_n1262), .A4(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1257), .A2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n824), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n776), .B1(new_n213), .B2(new_n855), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1266), .B(new_n1267), .C1(new_n920), .C2(new_n834), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1268), .B1(new_n1244), .B2(new_n773), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1248), .A2(new_n1270), .ZN(G381));
  INV_X1    g1071(.A(G390), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n841), .B(new_n1095), .C1(new_n1096), .C2(new_n1097), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1272), .A2(new_n882), .A3(new_n1274), .ZN(new_n1275));
  NOR3_X1   g1075(.A1(G387), .A2(new_n1275), .A3(G381), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1149), .B1(new_n1167), .B2(new_n773), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1247), .A2(KEYINPUT118), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n718), .B1(new_n1165), .B2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1167), .A2(new_n1181), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1277), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1276), .A2(new_n1281), .A3(new_n1209), .A4(new_n1236), .ZN(G407));
  INV_X1    g1082(.A(G213), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1283), .A2(G343), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1281), .A2(new_n1284), .ZN(new_n1285));
  OAI211_X1 g1085(.A(G407), .B(G213), .C1(G375), .C2(new_n1285), .ZN(G409));
  OAI211_X1 g1086(.A(G378), .B(new_n1236), .C1(new_n1201), .C2(new_n1208), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1206), .A2(new_n1207), .A3(new_n1035), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1236), .A2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1281), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1287), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1284), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(KEYINPUT60), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1239), .A2(new_n1294), .A3(new_n1246), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1245), .A2(KEYINPUT60), .A3(new_n1174), .A4(new_n1179), .ZN(new_n1296));
  AND2_X1   g1096(.A1(new_n1296), .A2(new_n717), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1270), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n882), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1298), .A2(G384), .A3(new_n1270), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1284), .A2(KEYINPUT125), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1300), .A2(new_n1301), .A3(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1303), .A2(G2897), .A3(new_n1284), .ZN(new_n1304));
  AOI21_X1  g1104(.A(G384), .B1(new_n1298), .B2(new_n1270), .ZN(new_n1305));
  AOI211_X1 g1105(.A(new_n882), .B(new_n1269), .C1(new_n1295), .C2(new_n1297), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1284), .A2(G2897), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1307), .A2(new_n1308), .A3(new_n1302), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1293), .A2(new_n1304), .A3(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1291), .A2(new_n1292), .A3(new_n1307), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT63), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT61), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(G393), .A2(G396), .ZN(new_n1315));
  AND3_X1   g1115(.A1(G390), .A2(new_n1315), .A3(new_n1273), .ZN(new_n1316));
  AOI21_X1  g1116(.A(G390), .B1(new_n1273), .B2(new_n1315), .ZN(new_n1317));
  OAI21_X1  g1117(.A(G387), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1315), .A2(new_n1273), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(new_n1272), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(G390), .A2(new_n1315), .A3(new_n1273), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1320), .A2(new_n1063), .A3(new_n1038), .A4(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1318), .A2(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1284), .B1(new_n1287), .B2(new_n1290), .ZN(new_n1324));
  NOR3_X1   g1124(.A1(new_n1305), .A2(new_n1306), .A3(new_n1312), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1323), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1310), .A2(new_n1313), .A3(new_n1314), .A4(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(KEYINPUT126), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1308), .B1(new_n1307), .B2(new_n1302), .ZN(new_n1329));
  AND4_X1   g1129(.A1(new_n1300), .A2(new_n1301), .A3(new_n1308), .A4(new_n1302), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(KEYINPUT61), .B1(new_n1331), .B2(new_n1293), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT126), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1332), .A2(new_n1333), .A3(new_n1313), .A4(new_n1326), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1328), .A2(new_n1334), .ZN(new_n1335));
  OR2_X1    g1135(.A1(new_n1311), .A2(KEYINPUT62), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1311), .A2(KEYINPUT62), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1332), .A2(new_n1336), .A3(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1338), .A2(new_n1323), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1335), .A2(new_n1339), .ZN(G405));
  NAND2_X1  g1140(.A1(G375), .A2(new_n1281), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1341), .A2(new_n1287), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1342), .A2(KEYINPUT127), .A3(new_n1307), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1307), .A2(KEYINPUT127), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1341), .A2(new_n1287), .A3(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1343), .A2(new_n1345), .ZN(new_n1346));
  XNOR2_X1  g1146(.A(new_n1346), .B(new_n1323), .ZN(G402));
endmodule


