//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 1 0 1 0 0 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1 1 1 0 1 0 1 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n771,
    new_n773, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n989, new_n990, new_n991;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT14), .ZN(new_n203));
  OR3_X1    g002(.A1(new_n203), .A2(G29gat), .A3(G36gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(G29gat), .B2(G36gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT88), .B(G36gat), .ZN(new_n206));
  INV_X1    g005(.A(G29gat), .ZN(new_n207));
  OAI211_X1 g006(.A(new_n204), .B(new_n205), .C1(new_n206), .C2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G43gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n209), .A2(G50gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(G50gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT15), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n208), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n212), .A2(new_n210), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT90), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n210), .B1(new_n215), .B2(new_n211), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n216), .B1(new_n215), .B2(new_n211), .ZN(new_n217));
  XOR2_X1   g016(.A(KEYINPUT89), .B(KEYINPUT15), .Z(new_n218));
  AOI21_X1  g017(.A(new_n214), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n213), .B1(new_n219), .B2(new_n208), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT91), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI211_X1 g021(.A(KEYINPUT91), .B(new_n213), .C1(new_n219), .C2(new_n208), .ZN(new_n223));
  AND2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT16), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n225), .A2(G1gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(G15gat), .B(G22gat), .ZN(new_n227));
  MUX2_X1   g026(.A(G1gat), .B(new_n226), .S(new_n227), .Z(new_n228));
  XOR2_X1   g027(.A(new_n228), .B(G8gat), .Z(new_n229));
  NAND2_X1  g028(.A1(new_n224), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT17), .ZN(new_n231));
  OR2_X1    g030(.A1(new_n220), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT17), .B1(new_n222), .B2(new_n223), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n202), .B(new_n230), .C1(new_n235), .C2(new_n229), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT92), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT18), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT18), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n236), .A2(KEYINPUT92), .A3(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n224), .B(new_n229), .ZN(new_n241));
  XOR2_X1   g040(.A(new_n202), .B(KEYINPUT13), .Z(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n238), .A2(new_n240), .A3(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(G113gat), .B(G141gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(KEYINPUT11), .ZN(new_n246));
  INV_X1    g045(.A(G169gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G197gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n250), .B(KEYINPUT12), .Z(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n244), .A2(new_n252), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n238), .A2(new_n240), .A3(new_n243), .A4(new_n251), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  XOR2_X1   g055(.A(KEYINPUT31), .B(G50gat), .Z(new_n257));
  NAND2_X1  g056(.A1(G228gat), .A2(G233gat), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G197gat), .B(G204gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT22), .ZN(new_n261));
  XNOR2_X1  g060(.A(G211gat), .B(G218gat), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT74), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n261), .A2(KEYINPUT74), .A3(new_n263), .ZN(new_n267));
  AND2_X1   g066(.A1(G211gat), .A2(G218gat), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n262), .B(new_n260), .C1(KEYINPUT22), .C2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n266), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT29), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT3), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(G155gat), .A2(G162gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(G155gat), .A2(G162gat), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G148gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(G141gat), .ZN(new_n277));
  INV_X1    g076(.A(G141gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(G148gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT2), .ZN(new_n281));
  AOI211_X1 g080(.A(new_n273), .B(new_n275), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT77), .ZN(new_n283));
  AND3_X1   g082(.A1(new_n276), .A2(KEYINPUT76), .A3(G141gat), .ZN(new_n284));
  OAI21_X1  g083(.A(KEYINPUT76), .B1(new_n276), .B2(G141gat), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n284), .B1(new_n277), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n275), .B1(new_n281), .B2(new_n273), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n283), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n276), .A2(KEYINPUT76), .A3(G141gat), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT76), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n290), .B1(new_n278), .B2(G148gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n278), .A2(G148gat), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n289), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n273), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n274), .B1(new_n294), .B2(KEYINPUT2), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(KEYINPUT77), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n282), .B1(new_n288), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT3), .ZN(new_n298));
  AOI21_X1  g097(.A(KEYINPUT29), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  OAI221_X1 g098(.A(new_n259), .B1(new_n272), .B2(new_n297), .C1(new_n270), .C2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT81), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n264), .A2(new_n269), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT3), .B1(new_n302), .B2(new_n271), .ZN(new_n303));
  OAI22_X1  g102(.A1(new_n299), .A2(new_n270), .B1(new_n297), .B2(new_n303), .ZN(new_n304));
  XOR2_X1   g103(.A(new_n258), .B(KEYINPUT80), .Z(new_n305));
  AOI21_X1  g104(.A(new_n301), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n282), .ZN(new_n307));
  AND3_X1   g106(.A1(new_n293), .A2(KEYINPUT77), .A3(new_n295), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT77), .B1(new_n293), .B2(new_n295), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n307), .B(new_n298), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n270), .B1(new_n310), .B2(new_n271), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n297), .A2(new_n303), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n301), .B(new_n305), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n300), .B1(new_n306), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G22gat), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n305), .B1(new_n311), .B2(new_n312), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT81), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(new_n313), .ZN(new_n319));
  INV_X1    g118(.A(G22gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n319), .A2(new_n320), .A3(new_n300), .ZN(new_n321));
  XNOR2_X1  g120(.A(G78gat), .B(G106gat), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n316), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n322), .B1(new_n316), .B2(new_n321), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n257), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n322), .ZN(new_n326));
  INV_X1    g125(.A(new_n321), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n320), .B1(new_n319), .B2(new_n300), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n316), .A2(new_n321), .A3(new_n322), .ZN(new_n330));
  INV_X1    g129(.A(new_n257), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  AND2_X1   g131(.A1(new_n325), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT78), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n334), .B1(new_n297), .B2(new_n298), .ZN(new_n335));
  XNOR2_X1  g134(.A(G113gat), .B(G120gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n336), .A2(KEYINPUT1), .ZN(new_n337));
  XNOR2_X1  g136(.A(G127gat), .B(G134gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n338), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n340), .B1(KEYINPUT1), .B2(new_n336), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n343), .B1(new_n297), .B2(new_n298), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n345), .A2(KEYINPUT78), .A3(KEYINPUT3), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n335), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(G225gat), .A2(G233gat), .ZN(new_n348));
  OAI21_X1  g147(.A(KEYINPUT4), .B1(new_n345), .B2(new_n342), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT4), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n297), .A2(new_n350), .A3(new_n343), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n347), .A2(new_n348), .A3(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n297), .B(new_n343), .ZN(new_n354));
  INV_X1    g153(.A(new_n348), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT5), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT5), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n353), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(G1gat), .B(G29gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n362), .B(KEYINPUT0), .ZN(new_n363));
  XOR2_X1   g162(.A(G57gat), .B(G85gat), .Z(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  OR2_X1    g164(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT6), .B1(new_n361), .B2(new_n365), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT79), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n366), .A2(new_n367), .A3(KEYINPUT79), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n361), .A2(new_n365), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(KEYINPUT6), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n370), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  AND3_X1   g173(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT67), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT67), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(G183gat), .A2(G190gat), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n376), .B1(new_n380), .B2(new_n375), .ZN(new_n381));
  INV_X1    g180(.A(G176gat), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n247), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(G169gat), .A2(G176gat), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT65), .B1(new_n384), .B2(KEYINPUT23), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT65), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT23), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n386), .B(new_n387), .C1(G169gat), .C2(G176gat), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n383), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT25), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n390), .B1(new_n384), .B2(KEYINPUT23), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n381), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  AND2_X1   g191(.A1(new_n378), .A2(new_n379), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n393), .A2(new_n375), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n247), .A2(KEYINPUT64), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT64), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(G169gat), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n395), .A2(new_n397), .A3(KEYINPUT23), .A4(new_n382), .ZN(new_n398));
  INV_X1    g197(.A(new_n383), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n247), .A2(new_n382), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n386), .B1(new_n400), .B2(new_n387), .ZN(new_n401));
  NOR3_X1   g200(.A1(new_n384), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n398), .B(new_n399), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT66), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT66), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n405), .A3(new_n398), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n394), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n392), .B1(new_n407), .B2(KEYINPUT25), .ZN(new_n408));
  XNOR2_X1  g207(.A(KEYINPUT27), .B(G183gat), .ZN(new_n409));
  INV_X1    g208(.A(G190gat), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(KEYINPUT28), .A3(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT69), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT68), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT27), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n413), .B1(new_n414), .B2(G183gat), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n410), .B(new_n415), .C1(new_n409), .C2(new_n413), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT28), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n412), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(G183gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT27), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n414), .A2(G183gat), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n413), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n415), .A2(new_n410), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n412), .B(new_n417), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n411), .B1(new_n418), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n400), .B1(new_n383), .B2(KEYINPUT26), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n427), .B1(KEYINPUT26), .B2(new_n400), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n379), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT29), .B1(new_n408), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(G226gat), .A2(G233gat), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(KEYINPUT75), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n392), .ZN(new_n436));
  INV_X1    g235(.A(new_n394), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n385), .A2(new_n388), .ZN(new_n438));
  AND4_X1   g237(.A1(new_n405), .A2(new_n438), .A3(new_n399), .A4(new_n398), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n405), .B1(new_n389), .B2(new_n398), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n437), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n436), .B1(new_n441), .B2(new_n390), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n417), .B1(new_n422), .B2(new_n423), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT69), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n424), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n429), .B1(new_n445), .B2(new_n411), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n271), .B1(new_n442), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT75), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(new_n448), .A3(new_n433), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n433), .B1(new_n408), .B2(new_n431), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n435), .A2(new_n449), .A3(new_n451), .A4(new_n270), .ZN(new_n452));
  INV_X1    g251(.A(new_n270), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n432), .A2(new_n434), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n453), .B1(new_n454), .B2(new_n450), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT30), .ZN(new_n456));
  XNOR2_X1  g255(.A(G8gat), .B(G36gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(G64gat), .B(G92gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n457), .B(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n452), .A2(new_n455), .A3(new_n456), .A4(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n452), .A2(new_n455), .A3(new_n460), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT30), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n460), .B1(new_n452), .B2(new_n455), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n333), .B1(new_n374), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT36), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n343), .B1(new_n442), .B2(new_n446), .ZN(new_n469));
  NAND2_X1  g268(.A1(G227gat), .A2(G233gat), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n408), .A2(new_n342), .A3(new_n431), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n469), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT32), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT33), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  XOR2_X1   g275(.A(G15gat), .B(G43gat), .Z(new_n477));
  XNOR2_X1  g276(.A(new_n477), .B(KEYINPUT70), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n478), .B(KEYINPUT71), .ZN(new_n479));
  XNOR2_X1  g278(.A(G71gat), .B(G99gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n479), .B(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n474), .A2(new_n476), .A3(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n481), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n473), .B(KEYINPUT32), .C1(new_n483), .C2(new_n475), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT73), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n469), .A2(new_n472), .ZN(new_n487));
  OAI211_X1 g286(.A(KEYINPUT72), .B(KEYINPUT34), .C1(new_n487), .C2(new_n471), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT72), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n471), .B1(new_n469), .B2(new_n472), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT34), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n490), .A2(new_n491), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n488), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n486), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n488), .A2(new_n492), .A3(new_n493), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n485), .A2(new_n496), .A3(KEYINPUT73), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n468), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n494), .A2(new_n485), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n496), .A2(new_n484), .A3(new_n482), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT36), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  XOR2_X1   g301(.A(KEYINPUT86), .B(KEYINPUT37), .Z(new_n503));
  NAND3_X1  g302(.A1(new_n452), .A2(new_n455), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n459), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT37), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n506), .B1(new_n452), .B2(new_n455), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT38), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n435), .A2(new_n449), .A3(new_n451), .A4(new_n453), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n270), .B1(new_n454), .B2(new_n450), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT37), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT38), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n511), .A2(new_n504), .A3(new_n512), .A4(new_n459), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n508), .A2(new_n462), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n358), .A2(KEYINPUT84), .A3(new_n360), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT84), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n353), .A2(new_n359), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n359), .B1(new_n353), .B2(new_n356), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n365), .B(KEYINPUT82), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n515), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT85), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(new_n367), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(new_n373), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n522), .B1(new_n521), .B2(new_n367), .ZN(new_n525));
  NOR3_X1   g324(.A1(new_n514), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT87), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n347), .A2(new_n352), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(new_n355), .ZN(new_n529));
  OR2_X1    g328(.A1(new_n529), .A2(KEYINPUT39), .ZN(new_n530));
  INV_X1    g329(.A(new_n520), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT39), .B1(new_n354), .B2(new_n355), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT83), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI211_X1 g333(.A(KEYINPUT83), .B(KEYINPUT39), .C1(new_n354), .C2(new_n355), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n534), .A2(new_n529), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n530), .A2(new_n531), .A3(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT40), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n530), .A2(KEYINPUT40), .A3(new_n536), .A4(new_n531), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n539), .A2(new_n521), .A3(new_n540), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n325), .B(new_n332), .C1(new_n541), .C2(new_n465), .ZN(new_n542));
  NOR3_X1   g341(.A1(new_n526), .A2(new_n527), .A3(new_n542), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n508), .A2(new_n462), .A3(new_n513), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n523), .A2(new_n373), .ZN(new_n545));
  INV_X1    g344(.A(new_n525), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n542), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT87), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n467), .B(new_n502), .C1(new_n543), .C2(new_n549), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n485), .A2(new_n496), .A3(KEYINPUT73), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n496), .B1(new_n485), .B2(KEYINPUT73), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n374), .A2(new_n333), .A3(new_n465), .A4(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n499), .A2(new_n500), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n555), .A2(new_n325), .A3(new_n332), .ZN(new_n556));
  INV_X1    g355(.A(new_n465), .ZN(new_n557));
  NOR3_X1   g356(.A1(new_n556), .A2(KEYINPUT35), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n545), .A2(new_n546), .ZN(new_n559));
  AOI22_X1  g358(.A1(KEYINPUT35), .A2(new_n554), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n256), .B1(new_n550), .B2(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(G183gat), .B(G211gat), .Z(new_n563));
  OR2_X1    g362(.A1(G57gat), .A2(G64gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(G57gat), .A2(G64gat), .ZN(new_n565));
  INV_X1    g364(.A(G71gat), .ZN(new_n566));
  INV_X1    g365(.A(G78gat), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n564), .B(new_n565), .C1(new_n568), .C2(KEYINPUT9), .ZN(new_n569));
  XNOR2_X1  g368(.A(G71gat), .B(G78gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n571), .A2(KEYINPUT21), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT93), .ZN(new_n573));
  NAND2_X1  g372(.A1(G231gat), .A2(G233gat), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n573), .B(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G127gat), .B(G155gat), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n576), .B(new_n577), .Z(new_n578));
  XNOR2_X1  g377(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT94), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n229), .B1(KEYINPUT21), .B2(new_n571), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n576), .B(new_n577), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(new_n580), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n582), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n584), .B1(new_n582), .B2(new_n586), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n563), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n582), .A2(new_n586), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(new_n583), .ZN(new_n592));
  INV_X1    g391(.A(new_n563), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n592), .A2(new_n587), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G134gat), .B(G162gat), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT41), .ZN(new_n598));
  INV_X1    g397(.A(G232gat), .ZN(new_n599));
  INV_X1    g398(.A(G233gat), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n597), .B(new_n601), .ZN(new_n602));
  NOR3_X1   g401(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n603));
  OAI21_X1  g402(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(G85gat), .A2(G92gat), .ZN(new_n605));
  MUX2_X1   g404(.A(KEYINPUT7), .B(new_n604), .S(new_n605), .Z(new_n606));
  INV_X1    g405(.A(KEYINPUT8), .ZN(new_n607));
  INV_X1    g406(.A(G99gat), .ZN(new_n608));
  INV_X1    g407(.A(G106gat), .ZN(new_n609));
  OAI21_X1  g408(.A(KEYINPUT95), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT95), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n611), .A2(G99gat), .A3(G106gat), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n607), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n606), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G99gat), .B(G106gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT96), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n614), .A2(KEYINPUT96), .A3(new_n615), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n614), .A2(new_n615), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n603), .B1(new_n224), .B2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G190gat), .B(G218gat), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n232), .B1(new_n224), .B2(KEYINPUT17), .ZN(new_n626));
  AOI21_X1  g425(.A(KEYINPUT97), .B1(new_n626), .B2(new_n621), .ZN(new_n627));
  OAI211_X1 g426(.A(KEYINPUT97), .B(new_n621), .C1(new_n233), .C2(new_n234), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n623), .B(new_n625), .C1(new_n627), .C2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT98), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n602), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n630), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT97), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n634), .B1(new_n235), .B2(new_n622), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n628), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n625), .B1(new_n636), .B2(new_n623), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n632), .B1(new_n633), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n636), .A2(new_n623), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n624), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n640), .B(new_n630), .C1(new_n631), .C2(new_n602), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n571), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n621), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT10), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n620), .A2(new_n571), .A3(new_n616), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT99), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n645), .A2(KEYINPUT99), .A3(new_n646), .A4(new_n647), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n621), .A2(new_n646), .A3(new_n644), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(G230gat), .A2(G233gat), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(G120gat), .B(G148gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(G176gat), .B(G204gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n647), .ZN(new_n661));
  INV_X1    g460(.A(new_n656), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n657), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n661), .A2(new_n662), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n653), .B1(new_n650), .B2(new_n651), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n656), .B(KEYINPUT100), .Z(new_n667));
  OAI21_X1  g466(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(new_n660), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n664), .A2(new_n669), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n596), .A2(new_n643), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n562), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n374), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g475(.A1(new_n673), .A2(new_n557), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(G8gat), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(KEYINPUT42), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT16), .B(G8gat), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  MUX2_X1   g480(.A(new_n679), .B(KEYINPUT42), .S(new_n681), .Z(G1325gat));
  INV_X1    g481(.A(G15gat), .ZN(new_n683));
  INV_X1    g482(.A(new_n555), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n683), .B1(new_n672), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT101), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n685), .A2(new_n686), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT102), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n689), .B1(new_n498), .B2(new_n501), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n555), .A2(new_n468), .ZN(new_n691));
  OAI21_X1  g490(.A(KEYINPUT36), .B1(new_n551), .B2(new_n552), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n691), .A2(new_n692), .A3(KEYINPUT102), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n673), .A2(G15gat), .A3(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n687), .A2(new_n688), .A3(new_n695), .ZN(new_n696));
  XOR2_X1   g495(.A(new_n696), .B(KEYINPUT103), .Z(G1326gat));
  NOR2_X1   g496(.A1(new_n672), .A2(new_n333), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT43), .B(G22gat), .Z(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1327gat));
  INV_X1    g499(.A(new_n670), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n596), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n702), .A2(new_n642), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n562), .A2(new_n703), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n704), .A2(G29gat), .A3(new_n374), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n705), .B(KEYINPUT45), .Z(new_n706));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n642), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n709), .B1(new_n550), .B2(new_n561), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n527), .B1(new_n526), .B2(new_n542), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n547), .A2(KEYINPUT87), .A3(new_n548), .ZN(new_n712));
  AOI211_X1 g511(.A(new_n466), .B(new_n694), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n643), .B1(new_n713), .B2(new_n560), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n710), .B1(new_n714), .B2(new_n707), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n702), .A2(new_n256), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n717), .A2(new_n674), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n706), .B1(new_n207), .B2(new_n718), .ZN(G1328gat));
  INV_X1    g518(.A(new_n206), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n704), .A2(new_n465), .A3(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT46), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT104), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n717), .A2(new_n557), .ZN(new_n725));
  OAI221_X1 g524(.A(new_n724), .B1(new_n722), .B2(new_n721), .C1(new_n206), .C2(new_n725), .ZN(G1329gat));
  NAND2_X1  g525(.A1(new_n717), .A2(new_n694), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(G43gat), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT105), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT47), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n562), .A2(new_n209), .A3(new_n555), .A4(new_n703), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n730), .B(new_n732), .ZN(G1330gat));
  INV_X1    g532(.A(G50gat), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n466), .B1(new_n711), .B2(new_n712), .ZN(new_n735));
  INV_X1    g534(.A(new_n694), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n560), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n707), .B1(new_n737), .B2(new_n642), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n325), .A2(new_n332), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n550), .A2(new_n561), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n708), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n738), .A2(new_n739), .A3(new_n741), .A4(new_n716), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(KEYINPUT106), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT106), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n715), .A2(new_n744), .A3(new_n739), .A4(new_n716), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n734), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n704), .A2(G50gat), .A3(new_n333), .ZN(new_n747));
  OAI21_X1  g546(.A(KEYINPUT48), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT107), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n742), .A2(G50gat), .ZN(new_n750));
  OR3_X1    g549(.A1(new_n750), .A2(KEYINPUT48), .A3(new_n747), .ZN(new_n751));
  AND3_X1   g550(.A1(new_n748), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n749), .B1(new_n748), .B2(new_n751), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n752), .A2(new_n753), .ZN(G1331gat));
  NAND2_X1  g553(.A1(new_n735), .A2(new_n736), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n561), .ZN(new_n756));
  NOR4_X1   g555(.A1(new_n596), .A2(new_n255), .A3(new_n643), .A4(new_n701), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n674), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g560(.A1(new_n758), .A2(new_n465), .ZN(new_n762));
  OR2_X1    g561(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n763));
  NAND2_X1  g562(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(new_n763), .B2(new_n762), .ZN(new_n766));
  XOR2_X1   g565(.A(new_n766), .B(KEYINPUT108), .Z(G1333gat));
  OAI21_X1  g566(.A(G71gat), .B1(new_n758), .B2(new_n736), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n555), .A2(new_n566), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n758), .B2(new_n769), .ZN(new_n770));
  XNOR2_X1  g569(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n770), .B(new_n771), .ZN(G1334gat));
  NOR2_X1   g571(.A1(new_n758), .A2(new_n333), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(new_n567), .ZN(G1335gat));
  NOR3_X1   g573(.A1(new_n595), .A2(new_n255), .A3(new_n701), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n715), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(G85gat), .B1(new_n776), .B2(new_n374), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n595), .A2(new_n255), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n756), .A2(new_n643), .A3(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT51), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT110), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n779), .A2(KEYINPUT110), .A3(new_n780), .ZN(new_n784));
  OR2_X1    g583(.A1(new_n779), .A2(new_n780), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n374), .A2(G85gat), .A3(new_n701), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(KEYINPUT111), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n777), .B1(new_n787), .B2(new_n789), .ZN(G1336gat));
  NAND3_X1  g589(.A1(new_n715), .A2(new_n557), .A3(new_n775), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(KEYINPUT113), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT52), .B1(new_n792), .B2(G92gat), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT112), .ZN(new_n794));
  OR3_X1    g593(.A1(new_n701), .A2(G92gat), .A3(new_n465), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n794), .B1(new_n786), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n786), .A2(new_n794), .A3(new_n796), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n793), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n791), .A2(G92gat), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n795), .B1(new_n785), .B2(new_n781), .ZN(new_n802));
  OAI21_X1  g601(.A(KEYINPUT52), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n800), .A2(new_n803), .ZN(G1337gat));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n805), .B1(new_n776), .B2(new_n736), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(G99gat), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n776), .A2(new_n805), .A3(new_n736), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n555), .A2(new_n670), .A3(new_n608), .ZN(new_n809));
  OAI22_X1  g608(.A1(new_n807), .A2(new_n808), .B1(new_n787), .B2(new_n809), .ZN(G1338gat));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n715), .A2(new_n739), .A3(new_n775), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(G106gat), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n333), .A2(G106gat), .A3(new_n701), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n786), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n814), .B1(new_n786), .B2(new_n815), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n811), .B(new_n813), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n785), .A2(new_n781), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n815), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n813), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n822), .A2(new_n823), .A3(KEYINPUT53), .ZN(new_n824));
  AOI22_X1  g623(.A1(new_n820), .A2(new_n815), .B1(G106gat), .B2(new_n812), .ZN(new_n825));
  OAI21_X1  g624(.A(KEYINPUT115), .B1(new_n825), .B2(new_n811), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n819), .A2(new_n827), .ZN(G1339gat));
  AND4_X1   g627(.A1(new_n256), .A2(new_n595), .A3(new_n642), .A4(new_n701), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n666), .A2(new_n667), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n657), .A2(KEYINPUT54), .A3(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n832));
  INV_X1    g631(.A(new_n667), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n655), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n831), .A2(KEYINPUT55), .A3(new_n660), .A4(new_n834), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n835), .A2(new_n664), .ZN(new_n836));
  INV_X1    g635(.A(new_n830), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT54), .B1(new_n666), .B2(new_n662), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n660), .B(new_n834), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT55), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n836), .A2(new_n255), .A3(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n250), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n235), .A2(new_n229), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n202), .B1(new_n844), .B2(new_n230), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n241), .A2(new_n242), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n843), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n254), .A2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n670), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n842), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n642), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n638), .A2(new_n641), .A3(new_n841), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT117), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n853), .A2(new_n854), .A3(new_n849), .A4(new_n836), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n853), .A2(new_n849), .A3(new_n836), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(KEYINPUT117), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n852), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n829), .B1(new_n858), .B2(new_n596), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n859), .A2(new_n374), .A3(new_n557), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(new_n333), .A3(new_n553), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(G113gat), .B1(new_n862), .B2(new_n255), .ZN(new_n863));
  INV_X1    g662(.A(new_n860), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n864), .A2(new_n556), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n255), .A2(G113gat), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n863), .B1(new_n865), .B2(new_n866), .ZN(G1340gat));
  OR3_X1    g666(.A1(new_n861), .A2(G120gat), .A3(new_n701), .ZN(new_n868));
  INV_X1    g667(.A(new_n865), .ZN(new_n869));
  OAI21_X1  g668(.A(G120gat), .B1(new_n869), .B2(new_n701), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n870), .A2(KEYINPUT118), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n870), .A2(KEYINPUT118), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n868), .B1(new_n871), .B2(new_n872), .ZN(G1341gat));
  OAI21_X1  g672(.A(G127gat), .B1(new_n869), .B2(new_n596), .ZN(new_n874));
  OR3_X1    g673(.A1(new_n861), .A2(G127gat), .A3(new_n596), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(G1342gat));
  NAND2_X1  g675(.A1(new_n333), .A2(new_n553), .ZN(new_n877));
  NOR4_X1   g676(.A1(new_n864), .A2(G134gat), .A3(new_n877), .A4(new_n642), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n878), .B(KEYINPUT56), .ZN(new_n879));
  OAI21_X1  g678(.A(G134gat), .B1(new_n869), .B2(new_n642), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(G1343gat));
  NOR2_X1   g680(.A1(new_n694), .A2(new_n333), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n860), .A2(new_n278), .A3(new_n255), .A4(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT58), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n374), .A2(new_n557), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n736), .A2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT57), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n887), .B1(new_n859), .B2(new_n333), .ZN(new_n888));
  AOI22_X1  g687(.A1(new_n851), .A2(new_n642), .B1(new_n856), .B2(KEYINPUT117), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n595), .B1(new_n889), .B2(new_n855), .ZN(new_n890));
  OAI211_X1 g689(.A(KEYINPUT57), .B(new_n739), .C1(new_n890), .C2(new_n829), .ZN(new_n891));
  AOI211_X1 g690(.A(new_n256), .B(new_n886), .C1(new_n888), .C2(new_n891), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n883), .B(new_n884), .C1(new_n892), .C2(new_n278), .ZN(new_n893));
  INV_X1    g692(.A(new_n883), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n888), .A2(new_n891), .ZN(new_n895));
  INV_X1    g694(.A(new_n886), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT119), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT119), .ZN(new_n898));
  AOI211_X1 g697(.A(new_n898), .B(new_n886), .C1(new_n888), .C2(new_n891), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n255), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n894), .B1(new_n901), .B2(G141gat), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n893), .B1(new_n902), .B2(new_n884), .ZN(G1344gat));
  NAND2_X1  g702(.A1(new_n860), .A2(new_n882), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n904), .A2(G148gat), .A3(new_n701), .ZN(new_n905));
  XOR2_X1   g704(.A(new_n905), .B(KEYINPUT120), .Z(new_n906));
  INV_X1    g705(.A(KEYINPUT59), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n853), .A2(KEYINPUT121), .A3(new_n836), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n638), .A2(new_n641), .A3(new_n841), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n835), .A2(new_n664), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n849), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(KEYINPUT122), .A3(new_n852), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT122), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n848), .B1(new_n908), .B2(new_n912), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n643), .B1(new_n842), .B2(new_n850), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n915), .A2(new_n596), .A3(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(new_n829), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n333), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n891), .B1(new_n922), .B2(KEYINPUT57), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n923), .A2(KEYINPUT123), .A3(new_n670), .A4(new_n896), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n924), .A2(G148gat), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n923), .A2(new_n670), .A3(new_n896), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT123), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n907), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  AOI211_X1 g728(.A(KEYINPUT59), .B(new_n276), .C1(new_n900), .C2(new_n670), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n906), .B1(new_n929), .B2(new_n930), .ZN(G1345gat));
  NOR3_X1   g730(.A1(new_n897), .A2(new_n899), .A3(new_n596), .ZN(new_n932));
  INV_X1    g731(.A(G155gat), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n595), .A2(new_n933), .ZN(new_n934));
  OAI22_X1  g733(.A1(new_n932), .A2(new_n933), .B1(new_n904), .B2(new_n934), .ZN(G1346gat));
  INV_X1    g734(.A(G162gat), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n936), .B1(new_n900), .B2(new_n643), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n643), .A2(new_n936), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n904), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g738(.A(KEYINPUT124), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT124), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n897), .A2(new_n899), .A3(new_n642), .ZN(new_n942));
  OAI221_X1 g741(.A(new_n941), .B1(new_n904), .B2(new_n938), .C1(new_n942), .C2(new_n936), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n940), .A2(new_n943), .ZN(G1347gat));
  INV_X1    g743(.A(new_n877), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n674), .A2(new_n465), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n945), .B(new_n946), .C1(new_n890), .C2(new_n829), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n948), .A2(new_n395), .A3(new_n397), .A4(new_n255), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n946), .A2(new_n555), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n333), .B1(new_n950), .B2(KEYINPUT125), .ZN(new_n951));
  AOI211_X1 g750(.A(new_n951), .B(new_n859), .C1(KEYINPUT125), .C2(new_n950), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n952), .A2(new_n255), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n949), .B1(new_n953), .B2(new_n247), .ZN(G1348gat));
  NAND3_X1  g753(.A1(new_n948), .A2(new_n382), .A3(new_n670), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n952), .A2(new_n670), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n955), .B1(new_n956), .B2(new_n382), .ZN(G1349gat));
  AOI21_X1  g756(.A(new_n419), .B1(new_n952), .B2(new_n595), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n948), .A2(new_n409), .A3(new_n595), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT126), .ZN(new_n960));
  OAI22_X1  g759(.A1(new_n958), .A2(new_n959), .B1(new_n960), .B2(KEYINPUT60), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(KEYINPUT60), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n961), .B(new_n962), .ZN(G1350gat));
  AOI21_X1  g762(.A(new_n410), .B1(new_n952), .B2(new_n643), .ZN(new_n964));
  XOR2_X1   g763(.A(new_n964), .B(KEYINPUT61), .Z(new_n965));
  NAND3_X1  g764(.A1(new_n948), .A2(new_n410), .A3(new_n643), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(G1351gat));
  NAND2_X1  g766(.A1(new_n736), .A2(new_n946), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n859), .A2(new_n333), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g768(.A(G197gat), .B1(new_n969), .B2(new_n255), .ZN(new_n970));
  INV_X1    g769(.A(new_n923), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n971), .A2(new_n968), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n256), .A2(new_n249), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n970), .B1(new_n972), .B2(new_n973), .ZN(G1352gat));
  NOR2_X1   g773(.A1(new_n701), .A2(G204gat), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n969), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n976), .B(KEYINPUT127), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT62), .ZN(new_n978));
  XNOR2_X1  g777(.A(new_n977), .B(new_n978), .ZN(new_n979));
  INV_X1    g778(.A(G204gat), .ZN(new_n980));
  NOR3_X1   g779(.A1(new_n971), .A2(new_n701), .A3(new_n968), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n979), .B1(new_n980), .B2(new_n981), .ZN(G1353gat));
  INV_X1    g781(.A(new_n969), .ZN(new_n983));
  OR3_X1    g782(.A1(new_n983), .A2(G211gat), .A3(new_n596), .ZN(new_n984));
  NAND4_X1  g783(.A1(new_n923), .A2(new_n595), .A3(new_n736), .A4(new_n946), .ZN(new_n985));
  AND3_X1   g784(.A1(new_n985), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n986));
  AOI21_X1  g785(.A(KEYINPUT63), .B1(new_n985), .B2(G211gat), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n984), .B1(new_n986), .B2(new_n987), .ZN(G1354gat));
  INV_X1    g787(.A(G218gat), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n969), .A2(new_n989), .A3(new_n643), .ZN(new_n990));
  NOR3_X1   g789(.A1(new_n971), .A2(new_n642), .A3(new_n968), .ZN(new_n991));
  OAI21_X1  g790(.A(new_n990), .B1(new_n991), .B2(new_n989), .ZN(G1355gat));
endmodule


