

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583;

  NOR2_X2 U323 ( .A1(n557), .A2(n556), .ZN(n568) );
  INV_X1 U324 ( .A(KEYINPUT54), .ZN(n394) );
  AND2_X1 U325 ( .A1(G230GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U326 ( .A(n366), .B(n291), .ZN(n330) );
  XNOR2_X1 U327 ( .A(n424), .B(n330), .ZN(n334) );
  XNOR2_X1 U328 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U329 ( .A(n342), .B(n341), .ZN(n572) );
  XOR2_X1 U330 ( .A(G64GAT), .B(G204GAT), .Z(n293) );
  XNOR2_X1 U331 ( .A(G176GAT), .B(G92GAT), .ZN(n292) );
  XNOR2_X1 U332 ( .A(n293), .B(n292), .ZN(n336) );
  XOR2_X1 U333 ( .A(KEYINPUT89), .B(KEYINPUT21), .Z(n295) );
  XNOR2_X1 U334 ( .A(G197GAT), .B(G218GAT), .ZN(n294) );
  XNOR2_X1 U335 ( .A(n295), .B(n294), .ZN(n423) );
  XNOR2_X1 U336 ( .A(n336), .B(n423), .ZN(n306) );
  XOR2_X1 U337 ( .A(G36GAT), .B(G190GAT), .Z(n370) );
  XOR2_X1 U338 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n301) );
  XOR2_X1 U339 ( .A(KEYINPUT86), .B(KEYINPUT17), .Z(n297) );
  XNOR2_X1 U340 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n296) );
  XNOR2_X1 U341 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U342 ( .A(G169GAT), .B(n298), .Z(n449) );
  XNOR2_X1 U343 ( .A(G8GAT), .B(G183GAT), .ZN(n299) );
  XNOR2_X1 U344 ( .A(n299), .B(G211GAT), .ZN(n346) );
  XNOR2_X1 U345 ( .A(n449), .B(n346), .ZN(n300) );
  XNOR2_X1 U346 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U347 ( .A(n370), .B(n302), .Z(n304) );
  NAND2_X1 U348 ( .A1(G226GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U349 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U350 ( .A(n306), .B(n305), .ZN(n490) );
  XNOR2_X1 U351 ( .A(KEYINPUT121), .B(n490), .ZN(n392) );
  XOR2_X1 U352 ( .A(G22GAT), .B(G197GAT), .Z(n308) );
  XNOR2_X1 U353 ( .A(G169GAT), .B(G8GAT), .ZN(n307) );
  XNOR2_X1 U354 ( .A(n308), .B(n307), .ZN(n312) );
  XOR2_X1 U355 ( .A(KEYINPUT72), .B(KEYINPUT67), .Z(n310) );
  XNOR2_X1 U356 ( .A(G15GAT), .B(KEYINPUT68), .ZN(n309) );
  XNOR2_X1 U357 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U358 ( .A(n312), .B(n311), .Z(n317) );
  XOR2_X1 U359 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n314) );
  NAND2_X1 U360 ( .A1(G229GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U361 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U362 ( .A(KEYINPUT66), .B(n315), .ZN(n316) );
  XNOR2_X1 U363 ( .A(n317), .B(n316), .ZN(n322) );
  XOR2_X1 U364 ( .A(G50GAT), .B(G36GAT), .Z(n320) );
  XNOR2_X1 U365 ( .A(G1GAT), .B(KEYINPUT71), .ZN(n318) );
  XNOR2_X1 U366 ( .A(n318), .B(KEYINPUT70), .ZN(n358) );
  XNOR2_X1 U367 ( .A(G113GAT), .B(n358), .ZN(n319) );
  XNOR2_X1 U368 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U369 ( .A(n322), .B(n321), .Z(n327) );
  XOR2_X1 U370 ( .A(KEYINPUT7), .B(KEYINPUT69), .Z(n324) );
  XNOR2_X1 U371 ( .A(G43GAT), .B(G29GAT), .ZN(n323) );
  XNOR2_X1 U372 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U373 ( .A(KEYINPUT8), .B(n325), .Z(n378) );
  XNOR2_X1 U374 ( .A(n378), .B(G141GAT), .ZN(n326) );
  XNOR2_X1 U375 ( .A(n327), .B(n326), .ZN(n558) );
  XOR2_X1 U376 ( .A(KEYINPUT74), .B(KEYINPUT75), .Z(n329) );
  XNOR2_X1 U377 ( .A(G148GAT), .B(G106GAT), .ZN(n328) );
  XNOR2_X1 U378 ( .A(n329), .B(n328), .ZN(n424) );
  XOR2_X1 U379 ( .A(G99GAT), .B(G85GAT), .Z(n366) );
  XOR2_X1 U380 ( .A(KEYINPUT33), .B(KEYINPUT73), .Z(n332) );
  XNOR2_X1 U381 ( .A(KEYINPUT77), .B(KEYINPUT31), .ZN(n331) );
  XNOR2_X1 U382 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U383 ( .A(n334), .B(n333), .Z(n342) );
  XNOR2_X1 U384 ( .A(G71GAT), .B(G57GAT), .ZN(n335) );
  XNOR2_X1 U385 ( .A(n335), .B(KEYINPUT13), .ZN(n347) );
  XNOR2_X1 U386 ( .A(n336), .B(n347), .ZN(n340) );
  XOR2_X1 U387 ( .A(KEYINPUT76), .B(KEYINPUT32), .Z(n338) );
  XNOR2_X1 U388 ( .A(G120GAT), .B(G78GAT), .ZN(n337) );
  XOR2_X1 U389 ( .A(n338), .B(n337), .Z(n339) );
  XNOR2_X1 U390 ( .A(n572), .B(KEYINPUT41), .ZN(n560) );
  NAND2_X1 U391 ( .A1(n558), .A2(n560), .ZN(n345) );
  XOR2_X1 U392 ( .A(KEYINPUT46), .B(KEYINPUT109), .Z(n343) );
  XNOR2_X1 U393 ( .A(KEYINPUT108), .B(n343), .ZN(n344) );
  XNOR2_X1 U394 ( .A(n345), .B(n344), .ZN(n383) );
  XNOR2_X1 U395 ( .A(n347), .B(n346), .ZN(n362) );
  XOR2_X1 U396 ( .A(G15GAT), .B(G127GAT), .Z(n443) );
  XOR2_X1 U397 ( .A(KEYINPUT82), .B(KEYINPUT15), .Z(n349) );
  XNOR2_X1 U398 ( .A(G64GAT), .B(KEYINPUT81), .ZN(n348) );
  XNOR2_X1 U399 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U400 ( .A(n443), .B(n350), .Z(n352) );
  NAND2_X1 U401 ( .A1(G231GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U402 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U403 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n354) );
  XNOR2_X1 U404 ( .A(KEYINPUT84), .B(KEYINPUT83), .ZN(n353) );
  XNOR2_X1 U405 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U406 ( .A(n356), .B(n355), .Z(n360) );
  XNOR2_X1 U407 ( .A(G22GAT), .B(G155GAT), .ZN(n357) );
  XNOR2_X1 U408 ( .A(n357), .B(G78GAT), .ZN(n422) );
  XNOR2_X1 U409 ( .A(n358), .B(n422), .ZN(n359) );
  XNOR2_X1 U410 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U411 ( .A(n362), .B(n361), .ZN(n482) );
  INV_X1 U412 ( .A(n482), .ZN(n576) );
  XNOR2_X1 U413 ( .A(KEYINPUT107), .B(n576), .ZN(n565) );
  XOR2_X1 U414 ( .A(KEYINPUT10), .B(KEYINPUT65), .Z(n364) );
  XNOR2_X1 U415 ( .A(G106GAT), .B(G218GAT), .ZN(n363) );
  XNOR2_X1 U416 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U417 ( .A(n365), .B(KEYINPUT79), .Z(n368) );
  XNOR2_X1 U418 ( .A(G92GAT), .B(n366), .ZN(n367) );
  XNOR2_X1 U419 ( .A(n368), .B(n367), .ZN(n374) );
  XNOR2_X1 U420 ( .A(G50GAT), .B(G162GAT), .ZN(n369) );
  XNOR2_X1 U421 ( .A(n369), .B(KEYINPUT78), .ZN(n433) );
  XOR2_X1 U422 ( .A(n370), .B(n433), .Z(n372) );
  NAND2_X1 U423 ( .A1(G232GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U424 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U425 ( .A(n374), .B(n373), .Z(n380) );
  XOR2_X1 U426 ( .A(KEYINPUT11), .B(KEYINPUT80), .Z(n376) );
  XNOR2_X1 U427 ( .A(G134GAT), .B(KEYINPUT9), .ZN(n375) );
  XNOR2_X1 U428 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U429 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U430 ( .A(n380), .B(n379), .ZN(n567) );
  INV_X1 U431 ( .A(n567), .ZN(n381) );
  AND2_X1 U432 ( .A1(n565), .A2(n381), .ZN(n382) );
  AND2_X1 U433 ( .A1(n383), .A2(n382), .ZN(n385) );
  XNOR2_X1 U434 ( .A(KEYINPUT47), .B(KEYINPUT110), .ZN(n384) );
  XNOR2_X1 U435 ( .A(n385), .B(n384), .ZN(n390) );
  XOR2_X1 U436 ( .A(KEYINPUT36), .B(n567), .Z(n581) );
  NOR2_X1 U437 ( .A1(n581), .A2(n482), .ZN(n386) );
  XOR2_X1 U438 ( .A(KEYINPUT45), .B(n386), .Z(n387) );
  NOR2_X1 U439 ( .A1(n558), .A2(n387), .ZN(n388) );
  NAND2_X1 U440 ( .A1(n572), .A2(n388), .ZN(n389) );
  NAND2_X1 U441 ( .A1(n390), .A2(n389), .ZN(n391) );
  XNOR2_X1 U442 ( .A(n391), .B(KEYINPUT48), .ZN(n520) );
  NAND2_X1 U443 ( .A1(n392), .A2(n520), .ZN(n393) );
  XNOR2_X1 U444 ( .A(n393), .B(KEYINPUT122), .ZN(n395) );
  XNOR2_X1 U445 ( .A(n395), .B(n394), .ZN(n416) );
  XOR2_X1 U446 ( .A(G162GAT), .B(G85GAT), .Z(n397) );
  XNOR2_X1 U447 ( .A(G29GAT), .B(G1GAT), .ZN(n396) );
  XNOR2_X1 U448 ( .A(n397), .B(n396), .ZN(n401) );
  XOR2_X1 U449 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n399) );
  XNOR2_X1 U450 ( .A(G127GAT), .B(G148GAT), .ZN(n398) );
  XNOR2_X1 U451 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U452 ( .A(n401), .B(n400), .Z(n406) );
  XOR2_X1 U453 ( .A(KEYINPUT91), .B(G57GAT), .Z(n403) );
  NAND2_X1 U454 ( .A1(G225GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U455 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U456 ( .A(KEYINPUT1), .B(n404), .ZN(n405) );
  XNOR2_X1 U457 ( .A(n406), .B(n405), .ZN(n410) );
  XOR2_X1 U458 ( .A(KEYINPUT6), .B(G155GAT), .Z(n408) );
  XNOR2_X1 U459 ( .A(KEYINPUT4), .B(KEYINPUT5), .ZN(n407) );
  XNOR2_X1 U460 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U461 ( .A(n410), .B(n409), .Z(n415) );
  XOR2_X1 U462 ( .A(G120GAT), .B(KEYINPUT0), .Z(n412) );
  XNOR2_X1 U463 ( .A(G113GAT), .B(G134GAT), .ZN(n411) );
  XNOR2_X1 U464 ( .A(n412), .B(n411), .ZN(n442) );
  XNOR2_X1 U465 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n413) );
  XNOR2_X1 U466 ( .A(n413), .B(KEYINPUT2), .ZN(n425) );
  XNOR2_X1 U467 ( .A(n442), .B(n425), .ZN(n414) );
  XNOR2_X1 U468 ( .A(n415), .B(n414), .ZN(n487) );
  NAND2_X1 U469 ( .A1(n416), .A2(n487), .ZN(n417) );
  XOR2_X1 U470 ( .A(n417), .B(KEYINPUT64), .Z(n553) );
  XOR2_X1 U471 ( .A(KEYINPUT87), .B(KEYINPUT24), .Z(n419) );
  XNOR2_X1 U472 ( .A(KEYINPUT22), .B(KEYINPUT88), .ZN(n418) );
  XNOR2_X1 U473 ( .A(n419), .B(n418), .ZN(n421) );
  XOR2_X1 U474 ( .A(G204GAT), .B(G211GAT), .Z(n420) );
  XNOR2_X1 U475 ( .A(n421), .B(n420), .ZN(n429) );
  XOR2_X1 U476 ( .A(n423), .B(n422), .Z(n427) );
  XNOR2_X1 U477 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U478 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U479 ( .A(n429), .B(n428), .ZN(n431) );
  NAND2_X1 U480 ( .A1(G228GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U481 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U482 ( .A(n432), .B(KEYINPUT90), .Z(n435) );
  XNOR2_X1 U483 ( .A(n433), .B(KEYINPUT23), .ZN(n434) );
  XNOR2_X1 U484 ( .A(n435), .B(n434), .ZN(n554) );
  XOR2_X1 U485 ( .A(G183GAT), .B(G99GAT), .Z(n437) );
  XNOR2_X1 U486 ( .A(G43GAT), .B(G190GAT), .ZN(n436) );
  XNOR2_X1 U487 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U488 ( .A(KEYINPUT20), .B(KEYINPUT85), .Z(n439) );
  XNOR2_X1 U489 ( .A(G176GAT), .B(G71GAT), .ZN(n438) );
  XNOR2_X1 U490 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U491 ( .A(n441), .B(n440), .ZN(n447) );
  XOR2_X1 U492 ( .A(n443), .B(n442), .Z(n445) );
  NAND2_X1 U493 ( .A1(G227GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U494 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U495 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U496 ( .A(n449), .B(n448), .ZN(n557) );
  INV_X1 U497 ( .A(n557), .ZN(n523) );
  NOR2_X1 U498 ( .A1(n554), .A2(n523), .ZN(n450) );
  XNOR2_X1 U499 ( .A(n450), .B(KEYINPUT26), .ZN(n462) );
  NAND2_X1 U500 ( .A1(n553), .A2(n462), .ZN(n580) );
  INV_X1 U501 ( .A(n580), .ZN(n577) );
  NAND2_X1 U502 ( .A1(n577), .A2(n558), .ZN(n452) );
  XOR2_X1 U503 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n451) );
  XNOR2_X1 U504 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U505 ( .A(n453), .B(KEYINPUT59), .ZN(n455) );
  XOR2_X1 U506 ( .A(G197GAT), .B(KEYINPUT124), .Z(n454) );
  XNOR2_X1 U507 ( .A(n455), .B(n454), .ZN(G1352GAT) );
  XOR2_X1 U508 ( .A(KEYINPUT99), .B(KEYINPUT34), .Z(n471) );
  NAND2_X1 U509 ( .A1(n558), .A2(n572), .ZN(n485) );
  NOR2_X1 U510 ( .A1(n567), .A2(n482), .ZN(n456) );
  XNOR2_X1 U511 ( .A(KEYINPUT16), .B(n456), .ZN(n469) );
  NOR2_X1 U512 ( .A1(n490), .A2(n557), .ZN(n457) );
  XOR2_X1 U513 ( .A(KEYINPUT98), .B(n457), .Z(n458) );
  NAND2_X1 U514 ( .A1(n458), .A2(n554), .ZN(n459) );
  XOR2_X1 U515 ( .A(KEYINPUT25), .B(n459), .Z(n460) );
  NAND2_X1 U516 ( .A1(n487), .A2(n460), .ZN(n464) );
  XOR2_X1 U517 ( .A(n490), .B(KEYINPUT96), .Z(n461) );
  XNOR2_X1 U518 ( .A(KEYINPUT27), .B(n461), .ZN(n465) );
  NAND2_X1 U519 ( .A1(n462), .A2(n465), .ZN(n542) );
  XNOR2_X1 U520 ( .A(KEYINPUT97), .B(n542), .ZN(n463) );
  NOR2_X1 U521 ( .A1(n464), .A2(n463), .ZN(n468) );
  XNOR2_X1 U522 ( .A(n554), .B(KEYINPUT28), .ZN(n495) );
  NAND2_X1 U523 ( .A1(n465), .A2(n495), .ZN(n522) );
  NOR2_X1 U524 ( .A1(n522), .A2(n523), .ZN(n466) );
  NOR2_X1 U525 ( .A1(n487), .A2(n466), .ZN(n467) );
  NOR2_X1 U526 ( .A1(n468), .A2(n467), .ZN(n481) );
  NAND2_X1 U527 ( .A1(n469), .A2(n481), .ZN(n500) );
  NOR2_X1 U528 ( .A1(n485), .A2(n500), .ZN(n478) );
  INV_X1 U529 ( .A(n487), .ZN(n521) );
  NAND2_X1 U530 ( .A1(n478), .A2(n521), .ZN(n470) );
  XNOR2_X1 U531 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U532 ( .A(G1GAT), .B(n472), .ZN(G1324GAT) );
  INV_X1 U533 ( .A(n490), .ZN(n512) );
  NAND2_X1 U534 ( .A1(n512), .A2(n478), .ZN(n473) );
  XNOR2_X1 U535 ( .A(n473), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U536 ( .A(KEYINPUT35), .B(KEYINPUT101), .Z(n475) );
  NAND2_X1 U537 ( .A1(n478), .A2(n523), .ZN(n474) );
  XNOR2_X1 U538 ( .A(n475), .B(n474), .ZN(n477) );
  XOR2_X1 U539 ( .A(G15GAT), .B(KEYINPUT100), .Z(n476) );
  XNOR2_X1 U540 ( .A(n477), .B(n476), .ZN(G1326GAT) );
  INV_X1 U541 ( .A(n495), .ZN(n515) );
  NAND2_X1 U542 ( .A1(n478), .A2(n515), .ZN(n479) );
  XNOR2_X1 U543 ( .A(n479), .B(KEYINPUT102), .ZN(n480) );
  XNOR2_X1 U544 ( .A(G22GAT), .B(n480), .ZN(G1327GAT) );
  NAND2_X1 U545 ( .A1(n482), .A2(n481), .ZN(n483) );
  NOR2_X1 U546 ( .A1(n483), .A2(n581), .ZN(n484) );
  XNOR2_X1 U547 ( .A(n484), .B(KEYINPUT37), .ZN(n510) );
  NOR2_X1 U548 ( .A1(n510), .A2(n485), .ZN(n486) );
  XOR2_X1 U549 ( .A(KEYINPUT38), .B(n486), .Z(n496) );
  NOR2_X1 U550 ( .A1(n487), .A2(n496), .ZN(n488) );
  XNOR2_X1 U551 ( .A(n488), .B(KEYINPUT39), .ZN(n489) );
  XNOR2_X1 U552 ( .A(G29GAT), .B(n489), .ZN(G1328GAT) );
  NOR2_X1 U553 ( .A1(n490), .A2(n496), .ZN(n491) );
  XOR2_X1 U554 ( .A(G36GAT), .B(n491), .Z(G1329GAT) );
  NOR2_X1 U555 ( .A1(n496), .A2(n557), .ZN(n493) );
  XNOR2_X1 U556 ( .A(KEYINPUT103), .B(KEYINPUT40), .ZN(n492) );
  XNOR2_X1 U557 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U558 ( .A(G43GAT), .B(n494), .ZN(G1330GAT) );
  NOR2_X1 U559 ( .A1(n496), .A2(n495), .ZN(n497) );
  XOR2_X1 U560 ( .A(KEYINPUT104), .B(n497), .Z(n498) );
  XNOR2_X1 U561 ( .A(G50GAT), .B(n498), .ZN(G1331GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT42), .B(KEYINPUT105), .Z(n502) );
  INV_X1 U563 ( .A(n558), .ZN(n499) );
  NAND2_X1 U564 ( .A1(n499), .A2(n560), .ZN(n509) );
  NOR2_X1 U565 ( .A1(n509), .A2(n500), .ZN(n506) );
  NAND2_X1 U566 ( .A1(n506), .A2(n521), .ZN(n501) );
  XNOR2_X1 U567 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(n503), .ZN(G1332GAT) );
  NAND2_X1 U569 ( .A1(n512), .A2(n506), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n504), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U571 ( .A1(n506), .A2(n523), .ZN(n505) );
  XNOR2_X1 U572 ( .A(n505), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U573 ( .A(G78GAT), .B(KEYINPUT43), .Z(n508) );
  NAND2_X1 U574 ( .A1(n506), .A2(n515), .ZN(n507) );
  XNOR2_X1 U575 ( .A(n508), .B(n507), .ZN(G1335GAT) );
  NOR2_X1 U576 ( .A1(n510), .A2(n509), .ZN(n516) );
  NAND2_X1 U577 ( .A1(n516), .A2(n521), .ZN(n511) );
  XNOR2_X1 U578 ( .A(G85GAT), .B(n511), .ZN(G1336GAT) );
  NAND2_X1 U579 ( .A1(n512), .A2(n516), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n513), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U581 ( .A1(n516), .A2(n523), .ZN(n514) );
  XNOR2_X1 U582 ( .A(n514), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT106), .B(KEYINPUT44), .Z(n518) );
  NAND2_X1 U584 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U586 ( .A(G106GAT), .B(n519), .Z(G1339GAT) );
  XNOR2_X1 U587 ( .A(G113GAT), .B(KEYINPUT112), .ZN(n527) );
  NAND2_X1 U588 ( .A1(n520), .A2(n521), .ZN(n541) );
  NOR2_X1 U589 ( .A1(n522), .A2(n541), .ZN(n524) );
  NAND2_X1 U590 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n525), .B(KEYINPUT111), .ZN(n537) );
  NAND2_X1 U592 ( .A1(n558), .A2(n537), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n527), .B(n526), .ZN(G1340GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT49), .B(KEYINPUT114), .Z(n529) );
  NAND2_X1 U595 ( .A1(n537), .A2(n560), .ZN(n528) );
  XNOR2_X1 U596 ( .A(n529), .B(n528), .ZN(n531) );
  XOR2_X1 U597 ( .A(G120GAT), .B(KEYINPUT113), .Z(n530) );
  XNOR2_X1 U598 ( .A(n531), .B(n530), .ZN(G1341GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n533) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n532) );
  XNOR2_X1 U601 ( .A(n533), .B(n532), .ZN(n536) );
  INV_X1 U602 ( .A(n537), .ZN(n534) );
  NOR2_X1 U603 ( .A1(n565), .A2(n534), .ZN(n535) );
  XOR2_X1 U604 ( .A(n536), .B(n535), .Z(G1342GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n539) );
  NAND2_X1 U606 ( .A1(n537), .A2(n567), .ZN(n538) );
  XNOR2_X1 U607 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U608 ( .A(G134GAT), .B(n540), .Z(G1343GAT) );
  XNOR2_X1 U609 ( .A(G141GAT), .B(KEYINPUT118), .ZN(n544) );
  NOR2_X1 U610 ( .A1(n542), .A2(n541), .ZN(n550) );
  NAND2_X1 U611 ( .A1(n558), .A2(n550), .ZN(n543) );
  XNOR2_X1 U612 ( .A(n544), .B(n543), .ZN(G1344GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT52), .B(KEYINPUT119), .Z(n546) );
  NAND2_X1 U614 ( .A1(n550), .A2(n560), .ZN(n545) );
  XNOR2_X1 U615 ( .A(n546), .B(n545), .ZN(n548) );
  XOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT53), .Z(n547) );
  XNOR2_X1 U617 ( .A(n548), .B(n547), .ZN(G1345GAT) );
  NAND2_X1 U618 ( .A1(n576), .A2(n550), .ZN(n549) );
  XNOR2_X1 U619 ( .A(n549), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U620 ( .A1(n550), .A2(n567), .ZN(n551) );
  XNOR2_X1 U621 ( .A(n551), .B(KEYINPUT120), .ZN(n552) );
  XNOR2_X1 U622 ( .A(G162GAT), .B(n552), .ZN(G1347GAT) );
  AND2_X1 U623 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n555), .B(KEYINPUT55), .ZN(n556) );
  INV_X1 U625 ( .A(n568), .ZN(n564) );
  NAND2_X1 U626 ( .A1(n568), .A2(n558), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n559), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U628 ( .A1(n568), .A2(n560), .ZN(n562) );
  XOR2_X1 U629 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n561) );
  XNOR2_X1 U630 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n563), .B(G176GAT), .ZN(G1349GAT) );
  NOR2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U633 ( .A(G183GAT), .B(n566), .Z(G1350GAT) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n570) );
  XOR2_X1 U635 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(G190GAT), .B(n571), .ZN(G1351GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n574) );
  OR2_X1 U639 ( .A1(n580), .A2(n572), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(G204GAT), .B(n575), .ZN(G1353GAT) );
  XOR2_X1 U642 ( .A(G211GAT), .B(KEYINPUT127), .Z(n579) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1354GAT) );
  NOR2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U646 ( .A(KEYINPUT62), .B(n582), .Z(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

