//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 1 1 1 0 0 1 1 0 1 0 0 1 1 0 1 1 1 0 0 0 0 1 1 0 1 0 0 1 1 1 0 0 0 1 1 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n562, new_n564, new_n565, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n627, new_n630, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1208,
    new_n1209, new_n1210;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT66), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  OR4_X1    g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n454), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND4_X1  g041(.A1(new_n463), .A2(new_n465), .A3(G137), .A4(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT69), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT3), .B(G2104), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n470), .A2(KEYINPUT69), .A3(G137), .A4(new_n466), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n462), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n463), .A2(new_n465), .ZN(new_n477));
  INV_X1    g052(.A(G125), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n475), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  AND3_X1   g057(.A1(new_n463), .A2(new_n465), .A3(G2105), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT70), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g060(.A(KEYINPUT70), .B1(new_n477), .B2(new_n466), .ZN(new_n486));
  AND2_X1   g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n477), .A2(G2105), .ZN(new_n489));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G112), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n462), .B1(new_n491), .B2(G2105), .ZN(new_n492));
  AOI22_X1  g067(.A1(new_n489), .A2(G136), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G162));
  INV_X1    g070(.A(KEYINPUT71), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(new_n466), .B2(G114), .ZN(new_n497));
  NOR2_X1   g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OR2_X1    g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(G114), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G2105), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n500), .A2(new_n502), .A3(KEYINPUT71), .A4(G2104), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n470), .A2(G126), .A3(G2105), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n463), .A2(new_n465), .A3(G138), .A4(new_n466), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n470), .A2(KEYINPUT4), .A3(G138), .A4(new_n466), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n504), .A2(new_n505), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(G164));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  OAI21_X1  g087(.A(KEYINPUT72), .B1(new_n512), .B2(KEYINPUT6), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n514), .A2(new_n515), .A3(G651), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n513), .A2(new_n516), .B1(KEYINPUT6), .B2(new_n512), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(G50), .B1(G75), .B2(G651), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT5), .B(G543), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n521), .A2(G62), .A3(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n513), .A2(new_n516), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n512), .A2(KEYINPUT6), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n523), .A2(new_n524), .A3(new_n521), .ZN(new_n525));
  XOR2_X1   g100(.A(KEYINPUT73), .B(G88), .Z(new_n526));
  OAI21_X1  g101(.A(new_n522), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n520), .A2(new_n527), .ZN(G166));
  NAND3_X1  g103(.A1(new_n517), .A2(G89), .A3(new_n521), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n517), .A2(G51), .A3(G543), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n529), .A2(new_n530), .A3(new_n532), .A4(new_n533), .ZN(G286));
  INV_X1    g109(.A(G286), .ZN(G168));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n519), .A2(KEYINPUT5), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT5), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G543), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(G64), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n536), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G651), .ZN(new_n543));
  XOR2_X1   g118(.A(KEYINPUT74), .B(G52), .Z(new_n544));
  NAND3_X1  g119(.A1(new_n517), .A2(G543), .A3(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(G90), .ZN(new_n546));
  OAI211_X1 g121(.A(new_n543), .B(new_n545), .C1(new_n546), .C2(new_n525), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  AND2_X1   g123(.A1(new_n517), .A2(G543), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G43), .ZN(new_n550));
  INV_X1    g125(.A(new_n525), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G81), .ZN(new_n552));
  NAND2_X1  g127(.A1(G68), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G56), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n540), .B2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT75), .ZN(new_n556));
  AND3_X1   g131(.A1(new_n555), .A2(new_n556), .A3(G651), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n556), .B1(new_n555), .B2(G651), .ZN(new_n558));
  OAI211_X1 g133(.A(new_n550), .B(new_n552), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  AND3_X1   g136(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G36), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n562), .A2(new_n565), .ZN(G188));
  NOR2_X1   g141(.A1(KEYINPUT78), .A2(G65), .ZN(new_n567));
  AND2_X1   g142(.A1(KEYINPUT78), .A2(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n521), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT77), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n512), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(G91), .ZN(new_n573));
  OAI21_X1  g148(.A(KEYINPUT76), .B1(new_n525), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT76), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n517), .A2(new_n575), .A3(G91), .A4(new_n521), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n572), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n523), .A2(G53), .A3(G543), .A4(new_n524), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT9), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(KEYINPUT79), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT79), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n577), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(G299));
  INV_X1    g159(.A(G166), .ZN(G303));
  NAND4_X1  g160(.A1(new_n523), .A2(G49), .A3(G543), .A4(new_n524), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n523), .A2(G87), .A3(new_n524), .A4(new_n521), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G288));
  AND4_X1   g164(.A1(G86), .A2(new_n523), .A3(new_n524), .A4(new_n521), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n523), .A2(G48), .A3(G543), .A4(new_n524), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(KEYINPUT81), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT81), .ZN(new_n593));
  NAND4_X1  g168(.A1(new_n517), .A2(new_n593), .A3(G48), .A4(G543), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n590), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n521), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n596));
  OAI21_X1  g171(.A(KEYINPUT80), .B1(new_n596), .B2(new_n512), .ZN(new_n597));
  NAND2_X1  g172(.A1(G73), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G61), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n540), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT80), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n600), .A2(new_n601), .A3(G651), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n595), .A2(new_n603), .ZN(G305));
  NAND2_X1  g179(.A1(G72), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G60), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n540), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n549), .A2(G47), .B1(G651), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n551), .A2(G85), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(G290));
  NAND2_X1  g185(.A1(G301), .A2(G868), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n517), .A2(G92), .A3(new_n521), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT10), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n612), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n549), .A2(KEYINPUT82), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n517), .A2(G543), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT82), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n615), .A2(G54), .A3(new_n618), .ZN(new_n619));
  AOI22_X1  g194(.A1(new_n521), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n620));
  OR2_X1    g195(.A1(new_n620), .A2(new_n512), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n614), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n611), .B1(new_n623), .B2(G868), .ZN(G284));
  OAI21_X1  g199(.A(new_n611), .B1(new_n623), .B2(G868), .ZN(G321));
  INV_X1    g200(.A(G868), .ZN(new_n626));
  NAND2_X1  g201(.A1(G299), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(new_n626), .B2(G168), .ZN(G297));
  OAI21_X1  g203(.A(new_n627), .B1(new_n626), .B2(G168), .ZN(G280));
  INV_X1    g204(.A(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n623), .B1(new_n630), .B2(G860), .ZN(G148));
  NAND2_X1  g206(.A1(new_n559), .A2(new_n626), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n622), .A2(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(new_n633), .B2(new_n626), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g210(.A1(new_n489), .A2(G135), .ZN(new_n636));
  NOR2_X1   g211(.A1(G99), .A2(G2105), .ZN(new_n637));
  OAI21_X1  g212(.A(G2104), .B1(new_n466), .B2(G111), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n485), .A2(new_n486), .ZN(new_n639));
  INV_X1    g214(.A(G123), .ZN(new_n640));
  OAI221_X1 g215(.A(new_n636), .B1(new_n637), .B2(new_n638), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(G2096), .Z(new_n642));
  NAND2_X1  g217(.A1(new_n470), .A2(new_n473), .ZN(new_n643));
  XOR2_X1   g218(.A(KEYINPUT83), .B(KEYINPUT12), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT13), .B(G2100), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n642), .A2(new_n647), .ZN(G156));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XOR2_X1   g225(.A(G2443), .B(G2446), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2427), .B(G2438), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2430), .ZN(new_n656));
  XOR2_X1   g231(.A(KEYINPUT15), .B(G2435), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(KEYINPUT14), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n654), .B(new_n659), .ZN(new_n660));
  AND2_X1   g235(.A1(new_n660), .A2(G14), .ZN(G401));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2067), .B(G2678), .Z(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n664), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n666), .A2(new_n667), .A3(KEYINPUT17), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT18), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2072), .B(G2078), .ZN(new_n671));
  OAI211_X1 g246(.A(new_n670), .B(new_n671), .C1(new_n669), .C2(new_n665), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n672), .B1(new_n671), .B2(new_n670), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2096), .B(G2100), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(G227));
  XNOR2_X1  g250(.A(G1971), .B(G1976), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT19), .ZN(new_n677));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n677), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n678), .A2(new_n679), .ZN(new_n683));
  AOI22_X1  g258(.A1(new_n681), .A2(KEYINPUT20), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n683), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n685), .A2(new_n677), .A3(new_n680), .ZN(new_n686));
  OAI211_X1 g261(.A(new_n684), .B(new_n686), .C1(KEYINPUT20), .C2(new_n681), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1986), .B(G1996), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G1981), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(G1991), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n689), .B(new_n692), .ZN(G229));
  INV_X1    g268(.A(G29), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G25), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT84), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n487), .A2(new_n696), .A3(G119), .ZN(new_n697));
  INV_X1    g272(.A(G119), .ZN(new_n698));
  OAI21_X1  g273(.A(KEYINPUT84), .B1(new_n639), .B2(new_n698), .ZN(new_n699));
  AOI22_X1  g274(.A1(new_n697), .A2(new_n699), .B1(G131), .B2(new_n489), .ZN(new_n700));
  OR2_X1    g275(.A1(G95), .A2(G2105), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n701), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n695), .B1(new_n703), .B2(new_n694), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT35), .B(G1991), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n704), .B(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT36), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(KEYINPUT87), .B2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G305), .ZN(new_n710));
  INV_X1    g285(.A(G16), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(G6), .B2(new_n711), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT32), .B(G1981), .Z(new_n714));
  OR2_X1    g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n711), .A2(G22), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G166), .B2(new_n711), .ZN(new_n717));
  AOI22_X1  g292(.A1(new_n713), .A2(new_n714), .B1(G1971), .B2(new_n717), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n717), .A2(G1971), .ZN(new_n719));
  NOR2_X1   g294(.A1(G16), .A2(G23), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT86), .ZN(new_n721));
  NAND2_X1  g296(.A1(G288), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g297(.A1(new_n586), .A2(new_n587), .A3(KEYINPUT86), .A4(new_n588), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n720), .B1(new_n724), .B2(G16), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT33), .B(G1976), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n715), .A2(new_n718), .A3(new_n719), .A4(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n709), .B1(KEYINPUT34), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n711), .A2(G24), .ZN(new_n730));
  INV_X1    g305(.A(G290), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(new_n711), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT85), .B(G1986), .Z(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n728), .A2(KEYINPUT34), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n729), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n708), .A2(KEYINPUT87), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n487), .A2(G129), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT93), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND3_X1  g316(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT26), .Z(new_n743));
  INV_X1    g318(.A(new_n489), .ZN(new_n744));
  INV_X1    g319(.A(G141), .ZN(new_n745));
  OR3_X1    g320(.A1(new_n744), .A2(KEYINPUT92), .A3(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(KEYINPUT92), .B1(new_n744), .B2(new_n745), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n746), .A2(new_n747), .B1(G105), .B2(new_n473), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n741), .A2(new_n743), .A3(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(G29), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G29), .B2(G32), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT27), .B(G1996), .Z(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n510), .A2(G29), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n694), .A2(G27), .ZN(new_n757));
  AND2_X1   g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G2078), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n751), .B(new_n753), .C1(G29), .C2(G32), .ZN(new_n761));
  OR2_X1    g336(.A1(G29), .A2(G33), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n470), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n763), .A2(new_n466), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n473), .A2(G103), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT25), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT90), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n489), .A2(G139), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n768), .B1(new_n767), .B2(new_n769), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n764), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n762), .B1(new_n773), .B2(new_n694), .ZN(new_n774));
  INV_X1    g349(.A(G2072), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n758), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n776), .B1(G2078), .B2(new_n777), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n755), .A2(new_n760), .A3(new_n761), .A4(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  AND2_X1   g355(.A1(KEYINPUT24), .A2(G34), .ZN(new_n781));
  NOR2_X1   g356(.A1(KEYINPUT24), .A2(G34), .ZN(new_n782));
  NOR3_X1   g357(.A1(new_n781), .A2(new_n782), .A3(G29), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n481), .B2(G29), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G2084), .ZN(new_n785));
  NOR2_X1   g360(.A1(G5), .A2(G16), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G171), .B2(G16), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(G1961), .ZN(new_n788));
  INV_X1    g363(.A(G28), .ZN(new_n789));
  AOI21_X1  g364(.A(G29), .B1(new_n789), .B2(KEYINPUT30), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(KEYINPUT30), .B2(new_n789), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n788), .B(new_n791), .C1(new_n694), .C2(new_n641), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n711), .A2(G21), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G168), .B2(new_n711), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1966), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT31), .B(G11), .Z(new_n796));
  NOR3_X1   g371(.A1(new_n792), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT94), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n774), .A2(new_n775), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT91), .Z(new_n800));
  NOR2_X1   g375(.A1(new_n787), .A2(G1961), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n780), .A2(new_n785), .A3(new_n798), .A4(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT95), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR3_X1   g380(.A1(new_n779), .A2(new_n800), .A3(new_n801), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n806), .A2(KEYINPUT95), .A3(new_n785), .A4(new_n798), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n711), .A2(G4), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(new_n623), .B2(new_n711), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT88), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT89), .B(G1348), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n694), .A2(G35), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G162), .B2(new_n694), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT29), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n711), .A2(G19), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n560), .B2(new_n711), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n815), .A2(G2090), .B1(G1341), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(G1341), .B2(new_n817), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT96), .B(KEYINPUT23), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n711), .A2(G20), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(G299), .B2(G16), .ZN(new_n823));
  INV_X1    g398(.A(G1956), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT28), .ZN(new_n826));
  INV_X1    g401(.A(G26), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n827), .B2(G29), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n827), .A2(G29), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n489), .A2(G140), .ZN(new_n830));
  NOR2_X1   g405(.A1(G104), .A2(G2105), .ZN(new_n831));
  OAI21_X1  g406(.A(G2104), .B1(new_n466), .B2(G116), .ZN(new_n832));
  INV_X1    g407(.A(G128), .ZN(new_n833));
  OAI221_X1 g408(.A(new_n830), .B1(new_n831), .B2(new_n832), .C1(new_n639), .C2(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n829), .B1(new_n834), .B2(G29), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n828), .B1(new_n835), .B2(new_n826), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(G2067), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n815), .B2(G2090), .ZN(new_n838));
  NOR4_X1   g413(.A1(new_n812), .A2(new_n819), .A3(new_n825), .A4(new_n838), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n738), .A2(new_n805), .A3(new_n807), .A4(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n836), .A2(G2067), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n736), .A2(new_n737), .ZN(new_n842));
  NOR3_X1   g417(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(G311));
  AND3_X1   g418(.A1(new_n805), .A2(new_n807), .A3(new_n839), .ZN(new_n844));
  INV_X1    g419(.A(new_n841), .ZN(new_n845));
  INV_X1    g420(.A(new_n842), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n844), .A2(new_n845), .A3(new_n846), .A4(new_n738), .ZN(G150));
  AOI22_X1  g422(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n848), .A2(new_n512), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n517), .A2(G55), .A3(G543), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n517), .A2(G93), .A3(new_n521), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT97), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(KEYINPUT97), .B1(new_n850), .B2(new_n851), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n849), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(G860), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(KEYINPUT37), .Z(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n560), .ZN(new_n859));
  OAI211_X1 g434(.A(new_n559), .B(new_n849), .C1(new_n855), .C2(new_n854), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT39), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n623), .A2(G559), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT38), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n862), .B(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n858), .B1(new_n865), .B2(G860), .ZN(G145));
  XNOR2_X1  g441(.A(new_n494), .B(new_n481), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n773), .A2(G164), .ZN(new_n868));
  INV_X1    g443(.A(new_n772), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(new_n770), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n510), .B1(new_n870), .B2(new_n764), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n703), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n489), .A2(G142), .ZN(new_n873));
  NOR2_X1   g448(.A1(G106), .A2(G2105), .ZN(new_n874));
  OAI21_X1  g449(.A(G2104), .B1(new_n466), .B2(G118), .ZN(new_n875));
  INV_X1    g450(.A(G130), .ZN(new_n876));
  OAI221_X1 g451(.A(new_n873), .B1(new_n874), .B2(new_n875), .C1(new_n639), .C2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n834), .B(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n700), .A2(new_n702), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n773), .A2(G164), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n870), .A2(new_n510), .A3(new_n764), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n872), .A2(new_n878), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n878), .B1(new_n872), .B2(new_n882), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n750), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n872), .A2(new_n882), .ZN(new_n886));
  INV_X1    g461(.A(new_n878), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n872), .A2(new_n878), .A3(new_n882), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n888), .A2(new_n749), .A3(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n641), .B(new_n645), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n885), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n891), .B1(new_n885), .B2(new_n890), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n867), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n891), .ZN(new_n895));
  NOR3_X1   g470(.A1(new_n883), .A2(new_n884), .A3(new_n750), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n749), .B1(new_n888), .B2(new_n889), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n867), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n885), .A2(new_n890), .A3(new_n891), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  XOR2_X1   g476(.A(KEYINPUT98), .B(G37), .Z(new_n902));
  NAND3_X1  g477(.A1(new_n894), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g479(.A1(new_n856), .A2(new_n626), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n731), .A2(G303), .ZN(new_n906));
  NAND2_X1  g481(.A1(G290), .A2(G166), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n724), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n906), .A2(new_n724), .A3(new_n907), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n910), .A2(new_n710), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n710), .B1(new_n910), .B2(new_n911), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(KEYINPUT42), .ZN(new_n915));
  XOR2_X1   g490(.A(new_n861), .B(new_n633), .Z(new_n916));
  INV_X1    g491(.A(new_n583), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n582), .B1(new_n577), .B2(new_n579), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n623), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT99), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n581), .A2(new_n583), .A3(new_n622), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n622), .B1(new_n581), .B2(new_n583), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(KEYINPUT99), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n916), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n922), .A2(new_n924), .A3(KEYINPUT41), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT41), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n919), .A2(new_n928), .A3(new_n921), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n926), .B1(new_n916), .B2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n915), .B(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n905), .B1(new_n932), .B2(new_n626), .ZN(G295));
  OAI21_X1  g508(.A(new_n905), .B1(new_n932), .B2(new_n626), .ZN(G331));
  INV_X1    g509(.A(new_n914), .ZN(new_n935));
  XNOR2_X1  g510(.A(G301), .B(G286), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n861), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n859), .A2(new_n860), .A3(new_n936), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n922), .A2(new_n924), .A3(new_n938), .A4(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT101), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n940), .B(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n938), .A2(KEYINPUT100), .A3(new_n939), .ZN(new_n943));
  INV_X1    g518(.A(new_n921), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT41), .B1(new_n944), .B2(new_n923), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT100), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n861), .A2(new_n946), .A3(new_n937), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n943), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT41), .B1(new_n922), .B2(new_n924), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n935), .B1(new_n942), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT43), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n943), .A2(new_n947), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(new_n925), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n938), .A2(new_n939), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n927), .A2(new_n929), .A3(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n954), .A2(new_n914), .A3(new_n956), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n951), .A2(new_n952), .A3(new_n902), .A4(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n954), .A2(new_n956), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n935), .ZN(new_n960));
  INV_X1    g535(.A(G37), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n960), .A2(new_n961), .A3(new_n957), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n958), .B1(new_n962), .B2(new_n952), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT44), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n940), .B(KEYINPUT101), .ZN(new_n966));
  OR2_X1    g541(.A1(new_n948), .A2(new_n949), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n914), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n957), .A2(new_n902), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT43), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT103), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT103), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n972), .B(KEYINPUT43), .C1(new_n968), .C2(new_n969), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n971), .A2(KEYINPUT44), .A3(new_n973), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n960), .A2(new_n952), .A3(new_n961), .A4(new_n957), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT102), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n975), .B(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n965), .B1(new_n974), .B2(new_n977), .ZN(G397));
  INV_X1    g553(.A(G1996), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n750), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n834), .B(G2067), .ZN(new_n981));
  OR2_X1    g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G1384), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n462), .B1(new_n501), .B2(G2105), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT71), .B1(new_n984), .B2(new_n500), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n497), .A2(new_n496), .A3(new_n498), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n505), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n508), .A2(new_n509), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n983), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n472), .A2(new_n480), .A3(G40), .A4(new_n474), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n979), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n994), .B(KEYINPUT104), .ZN(new_n995));
  AOI22_X1  g570(.A1(new_n982), .A2(new_n993), .B1(new_n750), .B2(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n703), .A2(new_n706), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n879), .A2(new_n705), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n993), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g575(.A(G290), .B(G1986), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1000), .B1(new_n993), .B2(new_n1001), .ZN(new_n1002));
  AND4_X1   g577(.A1(G40), .A2(new_n472), .A3(new_n480), .A4(new_n474), .ZN(new_n1003));
  XNOR2_X1  g578(.A(KEYINPUT106), .B(KEYINPUT50), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n510), .A2(new_n983), .A3(new_n1004), .ZN(new_n1005));
  AND2_X1   g580(.A1(new_n508), .A2(new_n509), .ZN(new_n1006));
  AOI22_X1  g581(.A1(new_n499), .A2(new_n503), .B1(new_n483), .B2(G126), .ZN(new_n1007));
  AOI21_X1  g582(.A(G1384), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n1003), .B(new_n1005), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT115), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1961), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n989), .A2(KEYINPUT50), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1014), .A2(KEYINPUT115), .A3(new_n1003), .A4(new_n1005), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1012), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g591(.A(KEYINPUT121), .B(KEYINPUT53), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n510), .A2(KEYINPUT45), .A3(new_n983), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n991), .A2(new_n1003), .A3(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1017), .B1(new_n1019), .B2(G2078), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n510), .A2(KEYINPUT45), .A3(new_n983), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT45), .B1(new_n510), .B2(new_n983), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n1021), .A2(new_n1022), .A3(new_n992), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1023), .A2(KEYINPUT53), .A3(new_n759), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1016), .A2(new_n1020), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(G171), .ZN(new_n1026));
  INV_X1    g601(.A(G2084), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1014), .A2(new_n1027), .A3(new_n1003), .A4(new_n1005), .ZN(new_n1028));
  OAI211_X1 g603(.A(G168), .B(new_n1028), .C1(new_n1023), .C2(G1966), .ZN(new_n1029));
  INV_X1    g604(.A(G1966), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1019), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(G168), .B1(new_n1031), .B2(new_n1028), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT51), .ZN(new_n1033));
  OAI211_X1 g608(.A(G8), .B(new_n1029), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1029), .A2(G8), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(KEYINPUT51), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT120), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1034), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1037), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT62), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1026), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT62), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT127), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G1976), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1046), .B1(new_n722), .B2(new_n723), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G8), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1049), .B1(new_n1003), .B2(new_n1008), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n1051));
  NAND2_X1  g626(.A1(G288), .A2(new_n1046), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1048), .A2(new_n1050), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT110), .ZN(new_n1054));
  OAI21_X1  g629(.A(G8), .B1(new_n989), .B2(new_n992), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1055), .A2(new_n1047), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT110), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1056), .A2(new_n1057), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1054), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT111), .ZN(new_n1060));
  INV_X1    g635(.A(G1981), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n595), .A2(new_n1061), .A3(new_n603), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1061), .B1(new_n595), .B2(new_n603), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1060), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT49), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT49), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1060), .B(new_n1066), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1065), .A2(new_n1050), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT109), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1069), .B1(new_n1056), .B2(new_n1051), .ZN(new_n1070));
  OAI211_X1 g645(.A(KEYINPUT109), .B(KEYINPUT52), .C1(new_n1055), .C2(new_n1047), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n1059), .A2(new_n1068), .A3(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(G8), .B1(new_n520), .B2(new_n527), .ZN(new_n1074));
  XNOR2_X1  g649(.A(KEYINPUT108), .B(KEYINPUT55), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n1074), .B(new_n1076), .ZN(new_n1077));
  XNOR2_X1  g652(.A(KEYINPUT105), .B(G1971), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1019), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n510), .A2(new_n1009), .A3(new_n983), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1003), .B(new_n1080), .C1(new_n1008), .C2(new_n1004), .ZN(new_n1081));
  XNOR2_X1  g656(.A(KEYINPUT107), .B(G2090), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1079), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1077), .B1(new_n1083), .B2(G8), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1082), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1014), .A2(new_n1003), .A3(new_n1005), .A4(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1079), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1088), .A2(G8), .A3(new_n1077), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1073), .A2(KEYINPUT125), .A3(new_n1085), .A4(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT125), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1059), .A2(new_n1068), .A3(new_n1089), .A4(new_n1072), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1091), .B1(new_n1092), .B2(new_n1084), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1094));
  OAI211_X1 g669(.A(KEYINPUT127), .B(KEYINPUT62), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1042), .A2(new_n1045), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1096));
  OR2_X1    g671(.A1(new_n1073), .A2(KEYINPUT112), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1089), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1073), .A2(KEYINPUT112), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G288), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1068), .A2(new_n1046), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1062), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1055), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1049), .B1(new_n1079), .B2(new_n1087), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT63), .B1(new_n1105), .B2(new_n1077), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1029), .A2(G8), .A3(G168), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n1098), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1097), .A2(new_n1099), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT63), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1073), .A2(new_n1085), .A3(new_n1089), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1110), .B1(new_n1111), .B2(new_n1107), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1104), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1096), .A2(new_n1100), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(KEYINPUT120), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1034), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT122), .ZN(new_n1118));
  OR2_X1    g693(.A1(new_n479), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n479), .A2(new_n1118), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1119), .A2(new_n1120), .A3(G2105), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1121), .A2(G40), .A3(new_n475), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT123), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT123), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1121), .A2(new_n1125), .A3(G40), .A4(new_n475), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n759), .A2(KEYINPUT53), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1123), .A2(new_n1124), .A3(new_n1126), .A4(new_n1127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1016), .A2(G301), .A3(new_n1020), .A4(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT54), .B1(new_n1026), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1116), .A2(new_n1117), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1016), .A2(new_n1020), .A3(new_n1128), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(G171), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1016), .A2(G301), .A3(new_n1020), .A4(new_n1024), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1134), .A2(KEYINPUT54), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(KEYINPUT126), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT126), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1134), .A2(new_n1138), .A3(KEYINPUT54), .A4(new_n1135), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  OR2_X1    g715(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1132), .A2(new_n1094), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT114), .ZN(new_n1143));
  XNOR2_X1  g718(.A(KEYINPUT56), .B(G2072), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1023), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT113), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1081), .A2(new_n1146), .A3(new_n824), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1146), .B1(new_n1081), .B2(new_n824), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1145), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  XOR2_X1   g725(.A(new_n580), .B(KEYINPUT57), .Z(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1143), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1081), .A2(new_n824), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(KEYINPUT113), .ZN(new_n1155));
  AOI22_X1  g730(.A1(new_n1155), .A2(new_n1147), .B1(new_n1023), .B2(new_n1144), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1156), .A2(KEYINPUT114), .A3(new_n1151), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT116), .ZN(new_n1158));
  INV_X1    g733(.A(new_n811), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1012), .A2(new_n1159), .A3(new_n1015), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n989), .A2(new_n992), .ZN(new_n1161));
  INV_X1    g736(.A(G2067), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1158), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1160), .A2(new_n1158), .A3(new_n1163), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1167), .A2(new_n622), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1156), .A2(new_n1151), .ZN(new_n1169));
  OAI211_X1 g744(.A(new_n1153), .B(new_n1157), .C1(new_n1168), .C2(new_n1169), .ZN(new_n1170));
  OR2_X1    g745(.A1(new_n622), .A2(KEYINPUT119), .ZN(new_n1171));
  AND3_X1   g746(.A1(new_n1160), .A2(new_n1158), .A3(new_n1163), .ZN(new_n1172));
  OAI211_X1 g747(.A(KEYINPUT60), .B(new_n1171), .C1(new_n1172), .C2(new_n1164), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1173), .A2(KEYINPUT119), .A3(new_n622), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n622), .A2(KEYINPUT119), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1167), .A2(KEYINPUT60), .A3(new_n1171), .A4(new_n1175), .ZN(new_n1176));
  OR3_X1    g751(.A1(new_n1172), .A2(new_n1164), .A3(KEYINPUT60), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1174), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g753(.A(KEYINPUT58), .B(G1341), .ZN(new_n1179));
  OAI22_X1  g754(.A1(new_n1019), .A2(G1996), .B1(new_n1161), .B2(new_n1179), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n1180), .A2(new_n560), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n1181), .A2(KEYINPUT117), .A3(KEYINPUT59), .ZN(new_n1182));
  OAI22_X1  g757(.A1(new_n1156), .A2(new_n1151), .B1(KEYINPUT118), .B2(KEYINPUT61), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT118), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1150), .A2(new_n1184), .A3(new_n1152), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1183), .A2(new_n1153), .A3(new_n1157), .A4(new_n1185), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1187));
  OAI21_X1  g762(.A(KEYINPUT61), .B1(new_n1169), .B2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1182), .B1(new_n1186), .B2(new_n1188), .ZN(new_n1189));
  XOR2_X1   g764(.A(KEYINPUT117), .B(KEYINPUT59), .Z(new_n1190));
  NAND2_X1  g765(.A1(new_n1181), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1178), .A2(new_n1189), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1142), .B1(new_n1170), .B2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1002), .B1(new_n1114), .B2(new_n1193), .ZN(new_n1194));
  XOR2_X1   g769(.A(new_n995), .B(KEYINPUT46), .Z(new_n1195));
  OAI21_X1  g770(.A(new_n993), .B1(new_n749), .B2(new_n981), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  XOR2_X1   g772(.A(new_n1197), .B(KEYINPUT47), .Z(new_n1198));
  NOR2_X1   g773(.A1(new_n834), .A2(G2067), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1199), .B1(new_n996), .B2(new_n998), .ZN(new_n1200));
  INV_X1    g775(.A(new_n993), .ZN(new_n1201));
  NOR3_X1   g776(.A1(new_n1201), .A2(G1986), .A3(G290), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1202), .B(KEYINPUT48), .ZN(new_n1203));
  OAI22_X1  g778(.A1(new_n1200), .A2(new_n1201), .B1(new_n1000), .B2(new_n1203), .ZN(new_n1204));
  NOR2_X1   g779(.A1(new_n1198), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1194), .A2(new_n1205), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g781(.A1(G401), .A2(G227), .ZN(new_n1208));
  AND2_X1   g782(.A1(new_n903), .A2(new_n1208), .ZN(new_n1209));
  NOR2_X1   g783(.A1(G229), .A2(new_n460), .ZN(new_n1210));
  AND3_X1   g784(.A1(new_n1209), .A2(new_n963), .A3(new_n1210), .ZN(G308));
  NAND3_X1  g785(.A1(new_n1209), .A2(new_n963), .A3(new_n1210), .ZN(G225));
endmodule


