//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 1 1 0 1 0 0 0 1 0 0 1 1 1 0 1 1 0 1 1 1 0 0 0 0 0 1 0 0 1 0 0 1 0 1 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1296, new_n1297,
    new_n1298, new_n1299, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  AND2_X1   g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G20), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n202), .A2(G50), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT64), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n217), .A2(new_n218), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n208), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n211), .B1(new_n213), .B2(new_n214), .C1(new_n224), .C2(KEYINPUT1), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G250), .B(G257), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT65), .ZN(new_n228));
  XOR2_X1   g0028(.A(G264), .B(G270), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n230), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  INV_X1    g0038(.A(G50), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n239), .A2(G68), .ZN(new_n240));
  INV_X1    g0040(.A(G68), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(G50), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n238), .B(new_n245), .ZN(G351));
  AND2_X1   g0046(.A1(G33), .A2(G41), .ZN(new_n247));
  NAND2_X1  g0047(.A1(G1), .A2(G13), .ZN(new_n248));
  OAI21_X1  g0048(.A(KEYINPUT66), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT66), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n212), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND4_X1  g0054(.A1(new_n249), .A2(new_n252), .A3(new_n254), .A4(G274), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n249), .A2(new_n252), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(new_n254), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n256), .B1(G226), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  OR2_X1    g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  AND2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n263), .A2(G223), .B1(new_n266), .B2(G77), .ZN(new_n267));
  AOI21_X1  g0067(.A(G1698), .B1(new_n261), .B2(new_n262), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G222), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n247), .A2(new_n248), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AND3_X1   g0072(.A1(new_n259), .A2(new_n272), .A3(KEYINPUT67), .ZN(new_n273));
  AOI21_X1  g0073(.A(KEYINPUT67), .B1(new_n259), .B2(new_n272), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G179), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n248), .ZN(new_n280));
  NOR2_X1   g0080(.A1(KEYINPUT8), .A2(G58), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT68), .B(G58), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT8), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n206), .A2(G33), .ZN(new_n286));
  INV_X1    g0086(.A(G150), .ZN(new_n287));
  NOR2_X1   g0087(.A1(G20), .A2(G33), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  OAI22_X1  g0089(.A1(new_n285), .A2(new_n286), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n290), .A2(KEYINPUT69), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n206), .B1(new_n201), .B2(new_n239), .ZN(new_n292));
  XOR2_X1   g0092(.A(new_n292), .B(KEYINPUT70), .Z(new_n293));
  OAI21_X1  g0093(.A(new_n293), .B1(new_n290), .B2(KEYINPUT69), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n280), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(G50), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n280), .B1(new_n205), .B2(G20), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n297), .B1(new_n298), .B2(G50), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n275), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n278), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n300), .B(KEYINPUT9), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n275), .A2(G200), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n276), .A2(G190), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT10), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT10), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n305), .A2(new_n310), .A3(new_n306), .A4(new_n307), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n304), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  OAI22_X1  g0112(.A1(new_n289), .A2(new_n239), .B1(new_n206), .B2(G68), .ZN(new_n313));
  INV_X1    g0113(.A(G77), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n286), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n280), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT11), .ZN(new_n317));
  OR2_X1    g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n317), .ZN(new_n319));
  OR3_X1    g0119(.A1(new_n296), .A2(KEYINPUT12), .A3(G68), .ZN(new_n320));
  OAI21_X1  g0120(.A(KEYINPUT12), .B1(new_n296), .B2(G68), .ZN(new_n321));
  AOI22_X1  g0121(.A1(G68), .A2(new_n298), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n318), .A2(new_n319), .A3(new_n322), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n323), .B(KEYINPUT73), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT14), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n256), .B1(G238), .B2(new_n258), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n268), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT3), .B(G33), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n328), .A2(G232), .A3(G1698), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n271), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT13), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n326), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n332), .B1(new_n326), .B2(new_n331), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n325), .B(G169), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n335), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n333), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n336), .B1(new_n277), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n325), .B1(new_n338), .B2(G169), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n324), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n324), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n338), .A2(G200), .ZN(new_n343));
  INV_X1    g0143(.A(G190), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n342), .B(new_n343), .C1(new_n344), .C2(new_n338), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n202), .B1(new_n283), .B2(new_n241), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n348), .A2(G20), .B1(G159), .B2(new_n288), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n261), .A2(new_n206), .A3(new_n262), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT7), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n261), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n262), .ZN(new_n353));
  AND3_X1   g0153(.A1(new_n352), .A2(KEYINPUT74), .A3(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(G68), .B1(new_n352), .B2(KEYINPUT74), .ZN(new_n355));
  OAI211_X1 g0155(.A(KEYINPUT16), .B(new_n349), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT16), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n288), .A2(G159), .ZN(new_n358));
  INV_X1    g0158(.A(G58), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(KEYINPUT68), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT68), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(G58), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n201), .B1(new_n363), .B2(G68), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n358), .B1(new_n364), .B2(new_n206), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n241), .B1(new_n352), .B2(new_n353), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n357), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n356), .A2(new_n280), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n285), .A2(new_n296), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n285), .B2(new_n298), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  AND3_X1   g0171(.A1(new_n249), .A2(G274), .A3(new_n252), .ZN(new_n372));
  INV_X1    g0172(.A(G226), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(G1698), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(G223), .B2(G1698), .ZN(new_n375));
  INV_X1    g0175(.A(G33), .ZN(new_n376));
  INV_X1    g0176(.A(G87), .ZN(new_n377));
  OAI22_X1  g0177(.A1(new_n375), .A2(new_n266), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n254), .A2(new_n372), .B1(new_n378), .B2(new_n271), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n249), .A2(new_n252), .A3(G232), .A4(new_n253), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n379), .A2(G179), .A3(new_n380), .ZN(new_n381));
  NOR2_X1   g0181(.A1(G223), .A2(G1698), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n382), .B1(new_n373), .B2(G1698), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n383), .A2(new_n328), .B1(G33), .B2(G87), .ZN(new_n384));
  INV_X1    g0184(.A(new_n271), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n255), .B(new_n380), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(G169), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n381), .A2(new_n387), .ZN(new_n388));
  AND3_X1   g0188(.A1(new_n371), .A2(new_n388), .A3(KEYINPUT18), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT18), .B1(new_n371), .B2(new_n388), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT75), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n379), .A2(new_n392), .A3(new_n344), .A4(new_n380), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT75), .B1(new_n386), .B2(G190), .ZN(new_n394));
  INV_X1    g0194(.A(G200), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n386), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n393), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n397), .A2(new_n368), .A3(new_n370), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT17), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n397), .A2(KEYINPUT17), .A3(new_n368), .A4(new_n370), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n391), .A2(new_n402), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n263), .A2(G238), .B1(new_n266), .B2(G107), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n328), .A2(G232), .A3(new_n260), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n271), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n258), .A2(G244), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n407), .A2(new_n255), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(G190), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n409), .A2(G200), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n298), .A2(G77), .ZN(new_n413));
  XOR2_X1   g0213(.A(new_n413), .B(KEYINPUT72), .Z(new_n414));
  XOR2_X1   g0214(.A(KEYINPUT8), .B(G58), .Z(new_n415));
  OR2_X1    g0215(.A1(new_n288), .A2(KEYINPUT71), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n288), .A2(KEYINPUT71), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  XNOR2_X1  g0218(.A(KEYINPUT15), .B(G87), .ZN(new_n419));
  OAI221_X1 g0219(.A(new_n418), .B1(new_n206), .B2(new_n314), .C1(new_n286), .C2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n296), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n420), .A2(new_n280), .B1(new_n314), .B2(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n411), .A2(new_n412), .A3(new_n414), .A4(new_n422), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n414), .A2(new_n422), .B1(new_n409), .B2(new_n301), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n410), .A2(new_n277), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n312), .A2(new_n347), .A3(new_n403), .A4(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  OAI211_X1 g0229(.A(G264), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT78), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n328), .A2(KEYINPUT78), .A3(G264), .A4(G1698), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n266), .A2(G303), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n328), .A2(G257), .A3(new_n260), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n432), .A2(new_n433), .A3(new_n434), .A4(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n271), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n205), .A2(G45), .ZN(new_n438));
  OR2_X1    g0238(.A1(KEYINPUT5), .A2(G41), .ZN(new_n439));
  NAND2_X1  g0239(.A1(KEYINPUT5), .A2(G41), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n441), .A2(G274), .A3(new_n249), .A4(new_n252), .ZN(new_n442));
  INV_X1    g0242(.A(G45), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(G1), .ZN(new_n444));
  INV_X1    g0244(.A(new_n440), .ZN(new_n445));
  NOR2_X1   g0245(.A1(KEYINPUT5), .A2(G41), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n447), .A2(new_n249), .A3(G270), .A4(new_n252), .ZN(new_n448));
  AND2_X1   g0248(.A1(new_n442), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n437), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT79), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n205), .A2(G33), .ZN(new_n453));
  AND2_X1   g0253(.A1(new_n296), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT80), .ZN(new_n455));
  INV_X1    g0255(.A(new_n280), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n454), .A2(new_n455), .A3(new_n456), .A4(G116), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n455), .B1(new_n296), .B2(G116), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n296), .A2(new_n453), .A3(new_n248), .A4(new_n279), .ZN(new_n459));
  INV_X1    g0259(.A(G116), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n279), .A2(new_n248), .B1(G20), .B2(new_n460), .ZN(new_n462));
  NAND2_X1  g0262(.A1(G33), .A2(G283), .ZN(new_n463));
  INV_X1    g0263(.A(G97), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n463), .B(new_n206), .C1(G33), .C2(new_n464), .ZN(new_n465));
  AND3_X1   g0265(.A1(new_n462), .A2(KEYINPUT20), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(KEYINPUT20), .B1(new_n462), .B2(new_n465), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n457), .B(new_n461), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT81), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n462), .A2(new_n465), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT20), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n462), .A2(KEYINPUT20), .A3(new_n465), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n475), .A2(KEYINPUT81), .A3(new_n461), .A4(new_n457), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n470), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n437), .A2(KEYINPUT79), .A3(new_n449), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n452), .A2(new_n477), .A3(G169), .A4(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT21), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n450), .A2(new_n277), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n477), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n301), .B1(new_n470), .B2(new_n476), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n484), .A2(new_n452), .A3(KEYINPUT21), .A4(new_n478), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n481), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n452), .A2(G200), .A3(new_n478), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT82), .ZN(new_n488));
  INV_X1    g0288(.A(new_n477), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n452), .A2(new_n478), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(G190), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n488), .B1(new_n487), .B2(new_n489), .ZN(new_n494));
  OAI21_X1  g0294(.A(KEYINPUT83), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n487), .A2(new_n489), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT82), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT83), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n497), .A2(new_n498), .A3(new_n492), .A4(new_n490), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n486), .B1(new_n495), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n296), .A2(G97), .ZN(new_n501));
  INV_X1    g0301(.A(new_n459), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n501), .B1(new_n502), .B2(G97), .ZN(new_n503));
  AOI21_X1  g0303(.A(KEYINPUT7), .B1(new_n266), .B2(new_n206), .ZN(new_n504));
  NOR4_X1   g0304(.A1(new_n264), .A2(new_n265), .A3(new_n351), .A4(G20), .ZN(new_n505));
  OAI21_X1  g0305(.A(G107), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n289), .A2(new_n314), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT6), .ZN(new_n508));
  AND2_X1   g0308(.A1(G97), .A2(G107), .ZN(new_n509));
  NOR2_X1   g0309(.A1(G97), .A2(G107), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(G107), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n512), .A2(KEYINPUT6), .A3(G97), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n507), .B1(new_n514), .B2(G20), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n456), .B1(new_n506), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT76), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI211_X1 g0318(.A(KEYINPUT76), .B(new_n456), .C1(new_n506), .C2(new_n515), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n503), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(G250), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n521));
  OAI211_X1 g0321(.A(G244), .B(new_n260), .C1(new_n264), .C2(new_n265), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT4), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n463), .B(new_n521), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(KEYINPUT4), .B1(new_n268), .B2(G244), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n271), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n447), .A2(new_n249), .A3(G257), .A4(new_n252), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n442), .A2(new_n527), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n526), .A2(new_n528), .A3(new_n277), .ZN(new_n529));
  AOI21_X1  g0329(.A(G169), .B1(new_n526), .B2(new_n528), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n520), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n514), .A2(G20), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n288), .A2(G77), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n512), .B1(new_n352), .B2(new_n353), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n280), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT76), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n516), .A2(new_n517), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n526), .A2(new_n528), .A3(new_n344), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n442), .A2(new_n527), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n268), .A2(KEYINPUT4), .A3(G244), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n522), .A2(new_n523), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n543), .A2(new_n544), .A3(new_n463), .A4(new_n521), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n542), .B1(new_n545), .B2(new_n271), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n541), .B1(new_n546), .B2(G200), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n540), .A2(new_n503), .A3(new_n547), .ZN(new_n548));
  NOR3_X1   g0348(.A1(new_n247), .A2(KEYINPUT66), .A3(new_n248), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n250), .B1(new_n212), .B2(new_n251), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n551), .A2(G264), .A3(new_n447), .ZN(new_n552));
  OAI211_X1 g0352(.A(G250), .B(new_n260), .C1(new_n264), .C2(new_n265), .ZN(new_n553));
  INV_X1    g0353(.A(G294), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n553), .B1(new_n376), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT85), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n263), .A2(new_n556), .A3(G257), .ZN(new_n557));
  OAI211_X1 g0357(.A(G257), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT85), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n555), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n442), .B(new_n552), .C1(new_n560), .C2(new_n385), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(G200), .ZN(new_n562));
  XNOR2_X1  g0362(.A(new_n558), .B(new_n556), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n271), .B1(new_n563), .B2(new_n555), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n564), .A2(G190), .A3(new_n442), .A4(new_n552), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n206), .B(G87), .C1(new_n264), .C2(new_n265), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT22), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT22), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n328), .A2(new_n568), .A3(new_n206), .A4(G87), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n206), .A2(KEYINPUT23), .A3(G107), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT23), .ZN(new_n572));
  OAI22_X1  g0372(.A1(new_n571), .A2(KEYINPUT84), .B1(new_n572), .B2(new_n512), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n572), .A2(new_n512), .A3(G20), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT84), .ZN(new_n575));
  AOI21_X1  g0375(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n576));
  OAI22_X1  g0376(.A1(new_n574), .A2(new_n575), .B1(new_n576), .B2(G20), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT24), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n570), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n579), .B1(new_n570), .B2(new_n578), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n280), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT25), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n296), .B2(G107), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NOR3_X1   g0386(.A1(new_n296), .A2(new_n584), .A3(G107), .ZN(new_n587));
  OAI22_X1  g0387(.A1(new_n586), .A2(new_n587), .B1(new_n512), .B2(new_n459), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n562), .A2(new_n565), .A3(new_n583), .A4(new_n589), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n532), .A2(new_n548), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n561), .A2(new_n301), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n564), .A2(new_n277), .A3(new_n442), .A4(new_n552), .ZN(new_n593));
  INV_X1    g0393(.A(new_n582), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n456), .B1(new_n594), .B2(new_n580), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n592), .B(new_n593), .C1(new_n595), .C2(new_n588), .ZN(new_n596));
  NAND3_X1  g0396(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n206), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n510), .A2(new_n377), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n206), .B(G68), .C1(new_n264), .C2(new_n265), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT19), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(new_n286), .B2(new_n464), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n280), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n419), .A2(new_n421), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n502), .A2(G87), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(G250), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(new_n443), .B2(G1), .ZN(new_n610));
  INV_X1    g0410(.A(G274), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n205), .A2(new_n611), .A3(G45), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n249), .A2(new_n252), .A3(new_n610), .A4(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT77), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n610), .A2(new_n612), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT77), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n615), .A2(new_n616), .A3(new_n249), .A4(new_n252), .ZN(new_n617));
  OAI211_X1 g0417(.A(G238), .B(new_n260), .C1(new_n264), .C2(new_n265), .ZN(new_n618));
  OAI211_X1 g0418(.A(G244), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n619));
  NAND2_X1  g0419(.A1(G33), .A2(G116), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n614), .A2(new_n617), .B1(new_n271), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n608), .B1(new_n622), .B2(G190), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n621), .A2(new_n271), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n616), .B1(new_n551), .B2(new_n615), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n610), .A2(new_n612), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n257), .A2(KEYINPUT77), .A3(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n624), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(G200), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n623), .A2(new_n629), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n277), .B(new_n624), .C1(new_n625), .C2(new_n627), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n605), .B(new_n606), .C1(new_n419), .C2(new_n459), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n631), .B(new_n632), .C1(G169), .C2(new_n622), .ZN(new_n633));
  AND4_X1   g0433(.A1(new_n591), .A2(new_n596), .A3(new_n630), .A4(new_n633), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n429), .A2(new_n500), .A3(new_n634), .ZN(G372));
  NAND3_X1  g0435(.A1(new_n345), .A2(new_n425), .A3(new_n424), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n402), .B1(new_n636), .B2(new_n341), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT87), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n638), .B1(new_n389), .B2(new_n390), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n371), .A2(new_n388), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT18), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n368), .A2(new_n370), .B1(new_n387), .B2(new_n381), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(KEYINPUT18), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n642), .A2(KEYINPUT87), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n639), .A2(new_n645), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n637), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n309), .A2(new_n311), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n304), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  AND4_X1   g0449(.A1(new_n481), .A2(new_n483), .A3(new_n485), .A4(new_n596), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n628), .A2(KEYINPUT86), .A3(G200), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT86), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n622), .B2(new_n395), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n623), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n654), .A2(new_n633), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n655), .A2(new_n532), .A3(new_n548), .A4(new_n590), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n650), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n526), .A2(new_n528), .A3(new_n277), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(new_n546), .B2(G169), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n659), .B1(new_n540), .B2(new_n503), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT26), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n660), .A2(new_n661), .A3(new_n633), .A4(new_n654), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n520), .A2(new_n630), .A3(new_n531), .A4(new_n633), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(KEYINPUT26), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n662), .A2(new_n664), .A3(new_n633), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n657), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n649), .B1(new_n428), .B2(new_n666), .ZN(G369));
  NAND3_X1  g0467(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT27), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n670), .A2(new_n205), .A3(new_n206), .A4(G13), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n669), .A2(G213), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g0472(.A(new_n672), .B(KEYINPUT88), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(G343), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n674), .B(KEYINPUT89), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(new_n489), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n500), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n486), .A2(new_n676), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n596), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT89), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n674), .B(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n583), .A2(new_n589), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n682), .B1(new_n590), .B2(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n596), .A2(new_n684), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n681), .A2(G330), .A3(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n688), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n689), .A2(new_n486), .A3(new_n675), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(G399));
  INV_X1    g0493(.A(new_n209), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(G41), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n599), .A2(G116), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(G1), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n214), .B2(new_n696), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n699), .B(KEYINPUT28), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n661), .B1(new_n655), .B2(new_n660), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n633), .B1(new_n663), .B2(KEYINPUT26), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n481), .A2(new_n483), .A3(new_n485), .A4(new_n596), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n591), .B(new_n655), .C1(new_n704), .C2(KEYINPUT90), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n704), .A2(KEYINPUT90), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n703), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n707), .A2(KEYINPUT91), .A3(KEYINPUT29), .A4(new_n675), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n707), .A2(KEYINPUT29), .A3(new_n675), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT91), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n662), .A2(new_n664), .A3(new_n633), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n704), .A2(new_n591), .A3(new_n655), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n684), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n710), .B1(new_n713), .B2(KEYINPUT29), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n708), .B1(new_n709), .B2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(G330), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n500), .A2(new_n634), .A3(new_n675), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n564), .A2(new_n552), .A3(new_n622), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n718), .A2(new_n482), .A3(new_n546), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n718), .A2(new_n482), .A3(KEYINPUT30), .A4(new_n546), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n546), .A2(G179), .A3(new_n622), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n723), .A2(new_n452), .A3(new_n478), .A4(new_n561), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n721), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n684), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n726), .B(KEYINPUT31), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n716), .B1(new_n717), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n715), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n700), .B1(new_n729), .B2(G1), .ZN(G364));
  AOI21_X1  g0530(.A(new_n248), .B1(G20), .B2(new_n301), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n344), .A2(G179), .A3(G200), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n206), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n206), .A2(G179), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n734), .A2(new_n344), .A3(G200), .ZN(new_n735));
  OAI22_X1  g0535(.A1(new_n733), .A2(new_n464), .B1(new_n735), .B2(new_n512), .ZN(new_n736));
  NOR2_X1   g0536(.A1(G190), .A2(G200), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G159), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XOR2_X1   g0540(.A(new_n740), .B(KEYINPUT32), .Z(new_n741));
  NOR2_X1   g0541(.A1(new_n206), .A2(new_n277), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n743), .A2(G190), .A3(new_n395), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n734), .A2(G190), .A3(G200), .ZN(new_n746));
  OAI22_X1  g0546(.A1(new_n745), .A2(new_n241), .B1(new_n746), .B2(new_n377), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n742), .A2(new_n737), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n742), .A2(G190), .A3(new_n395), .ZN(new_n749));
  OAI221_X1 g0549(.A(new_n328), .B1(new_n748), .B2(new_n314), .C1(new_n283), .C2(new_n749), .ZN(new_n750));
  OR4_X1    g0550(.A1(new_n736), .A2(new_n741), .A3(new_n747), .A4(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n742), .A2(G190), .A3(G200), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT93), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n752), .A2(new_n753), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n751), .B1(G50), .B2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n733), .ZN(new_n760));
  INV_X1    g0560(.A(new_n735), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n760), .A2(G294), .B1(new_n761), .B2(G283), .ZN(new_n762));
  INV_X1    g0562(.A(G317), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(KEYINPUT33), .ZN(new_n764));
  OR2_X1    g0564(.A1(new_n763), .A2(KEYINPUT33), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n744), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G303), .ZN(new_n767));
  OAI211_X1 g0567(.A(new_n762), .B(new_n766), .C1(new_n767), .C2(new_n746), .ZN(new_n768));
  INV_X1    g0568(.A(new_n749), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n328), .B1(new_n769), .B2(G322), .ZN(new_n770));
  INV_X1    g0570(.A(G311), .ZN(new_n771));
  INV_X1    g0571(.A(new_n738), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n772), .A2(KEYINPUT94), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(KEYINPUT94), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G329), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n770), .B1(new_n771), .B2(new_n748), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n768), .B(new_n777), .C1(G326), .C2(new_n758), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n731), .B1(new_n759), .B2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G13), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G20), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n205), .B1(new_n781), .B2(G45), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n695), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n694), .A2(new_n266), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n786), .A2(G355), .B1(new_n460), .B2(new_n694), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n694), .A2(new_n328), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n788), .B1(G45), .B2(new_n214), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n245), .A2(new_n443), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n787), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(KEYINPUT92), .B1(G13), .B2(G33), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR3_X1   g0593(.A1(KEYINPUT92), .A2(G13), .A3(G33), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(G20), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n731), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n785), .B1(new_n791), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n779), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT95), .ZN(new_n800));
  INV_X1    g0600(.A(new_n796), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n800), .B1(new_n681), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n681), .A2(G330), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(new_n785), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n681), .A2(G330), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(G396));
  INV_X1    g0606(.A(new_n748), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n744), .A2(G283), .B1(G116), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT97), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n758), .A2(G303), .ZN(new_n810));
  INV_X1    g0610(.A(new_n775), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G311), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n266), .B1(new_n749), .B2(new_n554), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n377), .A2(new_n735), .B1(new_n746), .B2(new_n512), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n813), .B(new_n814), .C1(G97), .C2(new_n760), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n809), .A2(new_n810), .A3(new_n812), .A4(new_n815), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n769), .A2(G143), .B1(new_n807), .B2(G159), .ZN(new_n817));
  INV_X1    g0617(.A(G137), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n817), .B1(new_n287), .B2(new_n745), .C1(new_n757), .C2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT34), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n811), .A2(G132), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n733), .A2(new_n283), .B1(new_n746), .B2(new_n239), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n266), .B(new_n823), .C1(G68), .C2(new_n761), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n821), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n819), .A2(new_n820), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n816), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n731), .ZN(new_n828));
  INV_X1    g0628(.A(new_n795), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n829), .A2(new_n731), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT96), .Z(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n785), .B1(new_n832), .B2(new_n314), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n426), .A2(new_n684), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n422), .A2(new_n414), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n423), .B1(new_n835), .B2(new_n675), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n834), .B1(new_n836), .B2(new_n426), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n828), .B(new_n833), .C1(new_n837), .C2(new_n795), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n675), .B(new_n837), .C1(new_n657), .C2(new_n665), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(KEYINPUT98), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT98), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(new_n713), .B2(new_n837), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n841), .A2(new_n843), .B1(new_n713), .B2(new_n837), .ZN(new_n844));
  INV_X1    g0644(.A(new_n728), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n784), .B1(new_n844), .B2(new_n845), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n839), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(G384));
  NAND2_X1  g0650(.A1(new_n514), .A2(KEYINPUT35), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n213), .A2(new_n460), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n514), .B2(KEYINPUT35), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT99), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n851), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(new_n854), .B2(new_n853), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT36), .Z(new_n857));
  AOI211_X1 g0657(.A(new_n314), .B(new_n214), .C1(new_n363), .C2(G68), .ZN(new_n858));
  XOR2_X1   g0658(.A(new_n240), .B(KEYINPUT100), .Z(new_n859));
  OAI211_X1 g0659(.A(G1), .B(new_n780), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  XOR2_X1   g0661(.A(new_n861), .B(KEYINPUT101), .Z(new_n862));
  INV_X1    g0662(.A(new_n834), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n841), .B2(new_n843), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT38), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n356), .A2(new_n280), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n349), .B1(new_n354), .B2(new_n355), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT16), .B1(new_n867), .B2(KEYINPUT102), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT102), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n869), .B(new_n349), .C1(new_n354), .C2(new_n355), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n866), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n370), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n673), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n400), .A2(new_n401), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n642), .A2(new_n644), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n388), .B1(new_n871), .B2(new_n872), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n873), .A2(new_n877), .A3(KEYINPUT37), .A4(new_n398), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n371), .A2(new_n673), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n640), .A2(new_n879), .A3(new_n398), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT37), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n865), .B1(new_n876), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n673), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n352), .A2(KEYINPUT74), .A3(new_n353), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT74), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n241), .B1(new_n504), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n365), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n456), .B1(new_n889), .B2(KEYINPUT16), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n357), .B1(new_n889), .B2(new_n869), .ZN(new_n891));
  INV_X1    g0691(.A(new_n870), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n885), .B1(new_n893), .B2(new_n370), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n391), .B2(new_n402), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n895), .A2(KEYINPUT38), .A3(new_n882), .A4(new_n878), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n884), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n342), .A2(new_n675), .ZN(new_n898));
  OR2_X1    g0698(.A1(new_n346), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n346), .A2(new_n898), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n864), .A2(new_n897), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n646), .A2(new_n885), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT104), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n874), .A2(new_n639), .A3(new_n645), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n885), .B1(new_n368), .B2(new_n370), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n879), .A2(new_n398), .A3(new_n638), .ZN(new_n910));
  INV_X1    g0710(.A(new_n371), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n908), .B1(new_n911), .B2(new_n397), .ZN(new_n912));
  AOI22_X1  g0712(.A1(KEYINPUT37), .A2(new_n910), .B1(new_n912), .B2(new_n640), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n879), .A2(new_n398), .ZN(new_n914));
  NOR4_X1   g0714(.A1(new_n914), .A2(new_n638), .A3(new_n881), .A4(new_n643), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n909), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n865), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT39), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n896), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n906), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT38), .B1(new_n909), .B2(new_n916), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n896), .A2(new_n919), .ZN(new_n923));
  NOR3_X1   g0723(.A1(new_n922), .A2(new_n923), .A3(KEYINPUT104), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT103), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(new_n897), .B2(KEYINPUT39), .ZN(new_n926));
  AOI211_X1 g0726(.A(KEYINPUT103), .B(new_n919), .C1(new_n884), .C2(new_n896), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n921), .A2(new_n924), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n339), .A2(new_n340), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n929), .A2(new_n324), .A3(new_n675), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n905), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n715), .A2(new_n429), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n649), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n933), .B(new_n935), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n901), .A2(new_n837), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n717), .A2(new_n727), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n918), .A2(new_n896), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n937), .A2(KEYINPUT40), .A3(new_n938), .A4(new_n939), .ZN(new_n940));
  XOR2_X1   g0740(.A(KEYINPUT105), .B(KEYINPUT40), .Z(new_n941));
  NAND3_X1  g0741(.A1(new_n938), .A2(new_n901), .A3(new_n837), .ZN(new_n942));
  INV_X1    g0742(.A(new_n897), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AND2_X1   g0744(.A1(new_n940), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n428), .B1(new_n717), .B2(new_n727), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n716), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n946), .B2(new_n945), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n936), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n205), .B2(new_n781), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n936), .A2(new_n948), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n862), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n952), .B(KEYINPUT106), .Z(G367));
  AND2_X1   g0753(.A1(new_n230), .A2(new_n788), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n797), .B1(new_n209), .B2(new_n419), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n784), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n744), .A2(G159), .B1(G50), .B2(new_n807), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n758), .A2(G143), .B1(KEYINPUT112), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n328), .B1(new_n738), .B2(new_n818), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(G150), .B2(new_n769), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n314), .A2(new_n735), .B1(new_n746), .B2(new_n283), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(G68), .B2(new_n760), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n957), .A2(KEYINPUT112), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n958), .A2(new_n960), .A3(new_n962), .A4(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n735), .A2(new_n464), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n965), .B1(G107), .B2(new_n760), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n966), .B1(new_n554), .B2(new_n745), .C1(new_n757), .C2(new_n771), .ZN(new_n967));
  AOI22_X1  g0767(.A1(G283), .A2(new_n807), .B1(new_n772), .B2(G317), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n328), .B1(new_n769), .B2(G303), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT46), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n746), .B2(new_n460), .ZN(new_n971));
  INV_X1    g0771(.A(new_n746), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n972), .A2(KEYINPUT46), .A3(G116), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n968), .A2(new_n969), .A3(new_n971), .A4(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n964), .B1(new_n967), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT47), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n956), .B1(new_n976), .B2(new_n731), .ZN(new_n977));
  AND2_X1   g0777(.A1(new_n684), .A2(new_n608), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n633), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n655), .B2(new_n978), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n796), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n977), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT108), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n684), .A2(new_n520), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n984), .A2(new_n532), .A3(new_n548), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n985), .A2(new_n596), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n684), .B1(new_n986), .B2(new_n532), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n660), .A2(new_n684), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n692), .A2(new_n989), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n990), .A2(KEYINPUT42), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(KEYINPUT42), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n987), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n980), .A2(KEYINPUT107), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT43), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n980), .A2(KEYINPUT107), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n995), .B2(new_n980), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n993), .A2(new_n998), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n987), .B(new_n997), .C1(new_n991), .C2(new_n992), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n983), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n997), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n993), .A2(new_n1002), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1003), .B(KEYINPUT108), .C1(new_n993), .C2(new_n998), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n690), .A2(new_n989), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1001), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n486), .A2(new_n675), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n691), .B1(new_n1011), .B2(new_n687), .ZN(new_n1012));
  OR3_X1    g0812(.A1(new_n1012), .A2(KEYINPUT110), .A3(new_n989), .ZN(new_n1013));
  OAI21_X1  g0813(.A(KEYINPUT110), .B1(new_n1012), .B2(new_n989), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT45), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1012), .A2(new_n989), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT44), .Z(new_n1019));
  NAND3_X1  g0819(.A1(new_n1013), .A2(KEYINPUT45), .A3(new_n1014), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1017), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n690), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1017), .A2(new_n1019), .A3(new_n690), .A4(new_n1020), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n689), .B(new_n1011), .Z(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n803), .B2(KEYINPUT111), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n803), .A2(KEYINPUT111), .A3(new_n1026), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n729), .B1(new_n1025), .B2(new_n1030), .ZN(new_n1031));
  XOR2_X1   g0831(.A(KEYINPUT109), .B(KEYINPUT41), .Z(new_n1032));
  XNOR2_X1  g0832(.A(new_n695), .B(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n783), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n982), .B1(new_n1010), .B2(new_n1034), .ZN(G387));
  INV_X1    g0835(.A(new_n1029), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1036), .A2(new_n1027), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n783), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n731), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n769), .A2(G317), .B1(new_n807), .B2(G303), .ZN(new_n1040));
  INV_X1    g0840(.A(G322), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1040), .B1(new_n771), .B2(new_n745), .C1(new_n757), .C2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT48), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n760), .A2(G283), .B1(new_n972), .B2(G294), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT49), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n735), .A2(new_n460), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n328), .B(new_n1051), .C1(G326), .C2(new_n772), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1049), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n758), .A2(G159), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n749), .A2(new_n239), .B1(new_n748), .B2(new_n241), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n266), .B(new_n1055), .C1(G150), .C2(new_n772), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n733), .A2(new_n419), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n965), .B(new_n1057), .C1(G77), .C2(new_n972), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n285), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n744), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1054), .A2(new_n1056), .A3(new_n1058), .A4(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1039), .B1(new_n1053), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n697), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n786), .A2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(G107), .B2(new_n209), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n788), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n415), .A2(new_n239), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT50), .Z(new_n1068));
  AOI211_X1 g0868(.A(G45), .B(new_n1063), .C1(G68), .C2(G77), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1066), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n234), .A2(G45), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1065), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n797), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n784), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT113), .Z(new_n1075));
  OR3_X1    g0875(.A1(new_n1062), .A2(KEYINPUT114), .A3(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(KEYINPUT114), .B1(new_n1062), .B2(new_n1075), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1076), .B(new_n1077), .C1(new_n689), .C2(new_n801), .ZN(new_n1078));
  AND2_X1   g0878(.A1(new_n1038), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1037), .A2(new_n729), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n1036), .A2(new_n1027), .B1(new_n728), .B2(new_n715), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1080), .A2(new_n695), .A3(new_n1081), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n1079), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(G393));
  INV_X1    g0884(.A(new_n1025), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1080), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1025), .A2(new_n1080), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1087), .A2(new_n1088), .A3(new_n695), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n989), .A2(new_n796), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1066), .A2(new_n238), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n797), .B1(new_n464), .B2(new_n209), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n784), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n757), .A2(new_n287), .B1(new_n739), .B2(new_n749), .ZN(new_n1094));
  XOR2_X1   g0894(.A(new_n1094), .B(KEYINPUT51), .Z(new_n1095));
  OAI22_X1  g0895(.A1(new_n745), .A2(new_n239), .B1(new_n735), .B2(new_n377), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n733), .A2(new_n314), .B1(new_n746), .B2(new_n241), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n807), .A2(new_n415), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n266), .B1(new_n772), .B2(G143), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n757), .A2(new_n763), .B1(new_n771), .B2(new_n749), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT52), .Z(new_n1103));
  OAI22_X1  g0903(.A1(new_n745), .A2(new_n767), .B1(new_n735), .B2(new_n512), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n266), .B1(new_n738), .B2(new_n1041), .C1(new_n554), .C2(new_n748), .ZN(new_n1105));
  INV_X1    g0905(.A(G283), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n733), .A2(new_n460), .B1(new_n746), .B2(new_n1106), .ZN(new_n1107));
  OR3_X1    g0907(.A1(new_n1104), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n1095), .A2(new_n1101), .B1(new_n1103), .B2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1093), .B1(new_n1109), .B2(new_n731), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1085), .A2(new_n783), .B1(new_n1090), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1089), .A2(new_n1111), .ZN(G390));
  NAND2_X1  g0912(.A1(new_n429), .A2(new_n728), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n934), .A2(new_n649), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT116), .ZN(new_n1116));
  AND4_X1   g0916(.A1(G330), .A2(new_n938), .A3(new_n901), .A4(new_n837), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n901), .B1(new_n728), .B2(new_n837), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1116), .B(new_n864), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n938), .A2(G330), .A3(new_n837), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n901), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n728), .A2(new_n837), .A3(new_n901), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n707), .A2(new_n675), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n836), .A2(new_n426), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n834), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1122), .A2(new_n1123), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1119), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n840), .A2(KEYINPUT98), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n713), .A2(new_n842), .A3(new_n837), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n834), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1132), .A2(new_n1116), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1115), .B1(new_n1128), .B2(new_n1133), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n930), .B(new_n939), .C1(new_n1126), .C2(new_n1121), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n931), .B1(new_n864), .B2(new_n901), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1135), .B1(new_n928), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT115), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n930), .B1(new_n1131), .B2(new_n1121), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n896), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n398), .A2(KEYINPUT37), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n894), .A2(new_n1142), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1143), .A2(new_n877), .B1(new_n881), .B2(new_n880), .ZN(new_n1144));
  AOI21_X1  g0944(.A(KEYINPUT38), .B1(new_n1144), .B2(new_n895), .ZN(new_n1145));
  OAI21_X1  g0945(.A(KEYINPUT39), .B1(new_n1141), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(KEYINPUT103), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n897), .A2(new_n925), .A3(KEYINPUT39), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n918), .A2(new_n920), .A3(new_n906), .ZN(new_n1150));
  OAI21_X1  g0950(.A(KEYINPUT104), .B1(new_n922), .B2(new_n923), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1140), .A2(new_n1149), .A3(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1153), .A2(KEYINPUT115), .A3(new_n1135), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1123), .B1(new_n1139), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1117), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1134), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n930), .B1(new_n922), .B2(new_n1141), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n707), .A2(new_n675), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1125), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n863), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1158), .B1(new_n1161), .B2(new_n901), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n1147), .A2(new_n1148), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n1138), .B(new_n1162), .C1(new_n1163), .C2(new_n1140), .ZN(new_n1164));
  AOI21_X1  g0964(.A(KEYINPUT115), .B1(new_n1153), .B2(new_n1135), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1117), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1156), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n1132), .A2(new_n1116), .B1(new_n1168), .B2(new_n1126), .ZN(new_n1169));
  OAI21_X1  g0969(.A(KEYINPUT116), .B1(new_n1168), .B2(new_n1131), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1114), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1166), .A2(new_n1167), .A3(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1157), .A2(new_n695), .A3(new_n1172), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n758), .A2(G128), .B1(G132), .B2(new_n769), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT117), .ZN(new_n1175));
  INV_X1    g0975(.A(G125), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n775), .A2(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(KEYINPUT54), .B(G143), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n328), .B1(new_n748), .B2(new_n1178), .C1(new_n745), .C2(new_n818), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n972), .A2(G150), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1180), .B(KEYINPUT53), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n733), .A2(new_n739), .B1(new_n735), .B2(new_n239), .ZN(new_n1182));
  NOR4_X1   g0982(.A1(new_n1177), .A2(new_n1179), .A3(new_n1181), .A4(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n758), .A2(G283), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n775), .A2(new_n554), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n745), .A2(new_n512), .B1(new_n314), .B2(new_n733), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n241), .A2(new_n735), .B1(new_n746), .B2(new_n377), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n266), .B1(new_n748), .B2(new_n464), .C1(new_n460), .C2(new_n749), .ZN(new_n1188));
  NOR4_X1   g0988(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n1175), .A2(new_n1183), .B1(new_n1184), .B2(new_n1189), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n784), .B1(new_n1059), .B2(new_n831), .C1(new_n1190), .C2(new_n1039), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(new_n1163), .B2(new_n829), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1139), .A2(new_n1154), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1156), .B1(new_n1193), .B2(new_n1117), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1192), .B1(new_n1194), .B2(new_n783), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1173), .A2(new_n1195), .ZN(G378));
  NAND2_X1  g0996(.A1(new_n300), .A2(new_n673), .ZN(new_n1197));
  OR2_X1    g0997(.A1(new_n312), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n312), .A2(new_n1197), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1198), .A2(new_n1199), .A3(new_n1201), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1203), .A2(new_n829), .A3(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n784), .B1(new_n831), .B2(G50), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n757), .A2(new_n460), .B1(new_n241), .B2(new_n733), .ZN(new_n1207));
  XOR2_X1   g1007(.A(new_n1207), .B(KEYINPUT118), .Z(new_n1208));
  AOI22_X1  g1008(.A1(new_n972), .A2(G77), .B1(new_n761), .B2(new_n363), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n464), .B2(new_n745), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n775), .A2(new_n1106), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n328), .A2(G41), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1212), .B1(new_n748), .B2(new_n419), .C1(new_n512), .C2(new_n749), .ZN(new_n1213));
  NOR4_X1   g1013(.A1(new_n1208), .A2(new_n1210), .A3(new_n1211), .A4(new_n1213), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n1214), .A2(KEYINPUT58), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(KEYINPUT58), .ZN(new_n1216));
  INV_X1    g1016(.A(G128), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n749), .A2(new_n1217), .B1(new_n748), .B2(new_n818), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(G132), .B2(new_n744), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1178), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n760), .A2(G150), .B1(new_n972), .B2(new_n1220), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1219), .B(new_n1221), .C1(new_n757), .C2(new_n1176), .ZN(new_n1222));
  OR2_X1    g1022(.A1(new_n1222), .A2(KEYINPUT59), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(KEYINPUT59), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n761), .A2(G159), .ZN(new_n1225));
  AOI211_X1 g1025(.A(G33), .B(G41), .C1(new_n772), .C2(G124), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1223), .A2(new_n1224), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1212), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1228), .B(new_n239), .C1(G33), .C2(G41), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1215), .A2(new_n1216), .A3(new_n1227), .A4(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1206), .B1(new_n1230), .B2(new_n731), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1205), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n932), .ZN(new_n1234));
  OAI21_X1  g1034(.A(KEYINPUT119), .B1(new_n1234), .B2(new_n904), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n940), .A2(new_n944), .A3(G330), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1236), .A2(new_n1204), .A3(new_n1203), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1238), .A2(G330), .A3(new_n944), .A4(new_n940), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1235), .A2(new_n1240), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1235), .A2(new_n1240), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1233), .B1(new_n1243), .B2(new_n783), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1114), .B1(new_n1194), .B2(new_n1245), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1240), .A2(new_n933), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n1237), .A2(new_n1239), .B1(new_n905), .B2(new_n932), .ZN(new_n1248));
  OAI21_X1  g1048(.A(KEYINPUT57), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n695), .B1(new_n1246), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1172), .A2(new_n1115), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT57), .B1(new_n1251), .B2(new_n1243), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1244), .B1(new_n1250), .B2(new_n1252), .ZN(G375));
  NAND2_X1  g1053(.A1(new_n1121), .A2(new_n829), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n784), .B1(new_n831), .B2(G68), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n745), .A2(new_n460), .B1(new_n746), .B2(new_n464), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1057), .B(new_n1256), .C1(G77), .C2(new_n761), .ZN(new_n1257));
  OAI221_X1 g1057(.A(new_n266), .B1(new_n748), .B2(new_n512), .C1(new_n1106), .C2(new_n749), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(new_n811), .B2(G303), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1257), .B(new_n1259), .C1(new_n554), .C2(new_n757), .ZN(new_n1260));
  XOR2_X1   g1060(.A(new_n1260), .B(KEYINPUT120), .Z(new_n1261));
  OAI221_X1 g1061(.A(new_n328), .B1(new_n748), .B2(new_n287), .C1(new_n283), .C2(new_n735), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n760), .A2(G50), .B1(new_n972), .B2(G159), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1263), .B(new_n1264), .C1(new_n775), .C2(new_n1217), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1266), .A2(KEYINPUT121), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n745), .A2(new_n1178), .B1(new_n818), .B2(new_n749), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1268), .B1(new_n758), .B2(G132), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT121), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1269), .B1(new_n1265), .B2(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1261), .B1(new_n1267), .B2(new_n1271), .ZN(new_n1272));
  OR2_X1    g1072(.A1(new_n1272), .A2(KEYINPUT122), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1039), .B1(new_n1272), .B2(KEYINPUT122), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1255), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n1245), .A2(new_n783), .B1(new_n1254), .B2(new_n1275), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1170), .A2(new_n1114), .A3(new_n1127), .A4(new_n1119), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1134), .A2(new_n1277), .A3(new_n1033), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1276), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(G381));
  INV_X1    g1080(.A(new_n1244), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1249), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n696), .B1(new_n1282), .B2(new_n1251), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1251), .A2(new_n1243), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT57), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1281), .B1(new_n1283), .B2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(G396), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n1079), .A2(new_n1288), .A3(new_n1082), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1289), .A2(new_n1089), .A3(new_n849), .A4(new_n1111), .ZN(new_n1290));
  NOR4_X1   g1090(.A1(G378), .A2(G381), .A3(new_n1290), .A4(G387), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT123), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1287), .A2(new_n1291), .A3(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1292), .B1(new_n1287), .B2(new_n1291), .ZN(new_n1294));
  OR2_X1    g1094(.A1(new_n1293), .A2(new_n1294), .ZN(G407));
  INV_X1    g1095(.A(G213), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(G378), .A2(G343), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1296), .B1(new_n1287), .B2(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1298), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(new_n1299), .B(KEYINPUT124), .ZN(G409));
  NOR2_X1   g1100(.A1(new_n1296), .A2(G343), .ZN(new_n1301));
  OAI211_X1 g1101(.A(G378), .B(new_n1244), .C1(new_n1250), .C2(new_n1252), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1251), .A2(new_n1243), .A3(new_n1033), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(new_n1240), .B(new_n933), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1233), .B1(new_n1304), .B2(new_n783), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1303), .A2(new_n1305), .ZN(new_n1306));
  AND2_X1   g1106(.A1(new_n1173), .A2(new_n1195), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1301), .B1(new_n1302), .B2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT60), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1277), .A2(new_n1310), .ZN(new_n1311));
  AND3_X1   g1111(.A1(new_n1311), .A2(new_n695), .A3(new_n1134), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT125), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1313), .B1(new_n1277), .B2(new_n1310), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1128), .A2(new_n1133), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1315), .A2(KEYINPUT125), .A3(KEYINPUT60), .A4(new_n1114), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1314), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1312), .A2(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(G384), .B1(new_n1318), .B2(new_n1276), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1275), .A2(new_n1254), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1320), .B1(new_n1315), .B2(new_n782), .ZN(new_n1321));
  AOI211_X1 g1121(.A(new_n849), .B(new_n1321), .C1(new_n1312), .C2(new_n1317), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1319), .A2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1309), .A2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT63), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1083), .A2(new_n1288), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1327), .A2(new_n1289), .ZN(new_n1328));
  OAI211_X1 g1128(.A(G390), .B(new_n982), .C1(new_n1034), .C2(new_n1010), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1329), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1328), .B1(new_n1330), .B2(KEYINPUT126), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(G387), .A2(new_n1089), .A3(new_n1111), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(new_n1329), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1331), .A2(new_n1333), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1332), .A2(new_n1328), .A3(new_n1329), .A4(KEYINPUT126), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1336), .A2(KEYINPUT61), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1301), .A2(G2897), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1338), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1339), .B1(new_n1319), .B2(new_n1322), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1311), .A2(new_n695), .A3(new_n1134), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1341), .B1(new_n1314), .B2(new_n1316), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n849), .B1(new_n1342), .B2(new_n1321), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1318), .A2(G384), .A3(new_n1276), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1343), .A2(new_n1344), .A3(new_n1338), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1340), .A2(new_n1345), .ZN(new_n1346));
  OR2_X1    g1146(.A1(new_n1309), .A2(new_n1346), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1309), .A2(KEYINPUT63), .A3(new_n1323), .ZN(new_n1348));
  NAND4_X1  g1148(.A1(new_n1326), .A2(new_n1337), .A3(new_n1347), .A4(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT62), .ZN(new_n1350));
  AND3_X1   g1150(.A1(new_n1309), .A2(new_n1350), .A3(new_n1323), .ZN(new_n1351));
  XNOR2_X1  g1151(.A(KEYINPUT127), .B(KEYINPUT61), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1352), .B1(new_n1309), .B2(new_n1346), .ZN(new_n1353));
  AOI21_X1  g1153(.A(new_n1350), .B1(new_n1309), .B2(new_n1323), .ZN(new_n1354));
  NOR3_X1   g1154(.A1(new_n1351), .A2(new_n1353), .A3(new_n1354), .ZN(new_n1355));
  AND2_X1   g1155(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1349), .B1(new_n1355), .B2(new_n1356), .ZN(G405));
  NAND2_X1  g1157(.A1(G375), .A2(new_n1307), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1358), .A2(new_n1302), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1356), .A2(new_n1359), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(new_n1336), .A2(new_n1302), .A3(new_n1358), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1360), .A2(new_n1361), .ZN(new_n1362));
  INV_X1    g1162(.A(new_n1323), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1362), .A2(new_n1363), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1360), .A2(new_n1323), .A3(new_n1361), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1364), .A2(new_n1365), .ZN(G402));
endmodule


