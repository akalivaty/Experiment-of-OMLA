//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 1 0 0 0 1 1 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 1 1 0 1 0 0 1 0 1 1 0 0 0 0 0 0 0 1 1 0 1 1 0 1 0 1 1 0 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n529, new_n530, new_n531, new_n532, new_n533, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n545,
    new_n546, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n556, new_n557, new_n558, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n592, new_n593, new_n596, new_n598,
    new_n599, new_n600, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G567), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  OR2_X1    g031(.A1(new_n456), .A2(KEYINPUT66), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(KEYINPUT66), .ZN(new_n458));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  OAI211_X1 g034(.A(new_n457), .B(new_n458), .C1(new_n459), .C2(new_n451), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G137), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT3), .B(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n470), .A2(new_n475), .ZN(G160));
  NAND2_X1  g051(.A1(new_n472), .A2(new_n471), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(KEYINPUT67), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n465), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT68), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT69), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n471), .B1(new_n463), .B2(new_n464), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(G124), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  AND2_X1   g066(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n492));
  OAI211_X1 g067(.A(G138), .B(new_n471), .C1(new_n492), .C2(new_n462), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n493), .B(KEYINPUT4), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT70), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n471), .A2(G114), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OR2_X1    g073(.A1(G102), .A2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(G114), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n499), .A2(new_n501), .A3(KEYINPUT70), .A4(G2104), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n472), .A2(G126), .A3(G2105), .ZN(new_n504));
  AND3_X1   g079(.A1(new_n503), .A2(KEYINPUT71), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g080(.A(KEYINPUT71), .B1(new_n503), .B2(new_n504), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n494), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  XNOR2_X1  g083(.A(KEYINPUT5), .B(G543), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n509), .A2(new_n510), .A3(G88), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n510), .A2(G50), .A3(G543), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  OAI211_X1 g089(.A(new_n511), .B(new_n512), .C1(new_n513), .C2(new_n514), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  NAND3_X1  g091(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n510), .A2(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G51), .ZN(new_n519));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n509), .A2(new_n510), .ZN(new_n522));
  INV_X1    g097(.A(G89), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT72), .ZN(new_n525));
  OAI211_X1 g100(.A(new_n517), .B(new_n519), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n524), .A2(new_n525), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(G168));
  INV_X1    g103(.A(new_n522), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n529), .A2(G90), .B1(new_n518), .B2(G52), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT73), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n530), .B(new_n531), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n514), .B2(new_n533), .ZN(G301));
  INV_X1    g109(.A(G301), .ZN(G171));
  INV_X1    g110(.A(G81), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n510), .A2(G543), .ZN(new_n537));
  INV_X1    g112(.A(G43), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n522), .A2(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n514), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  NAND4_X1  g118(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND4_X1  g121(.A1(G319), .A2(G483), .A3(G661), .A4(new_n546), .ZN(G188));
  NAND2_X1  g122(.A1(new_n518), .A2(G53), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT9), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n509), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(new_n514), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n529), .A2(G91), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n549), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  XOR2_X1   g128(.A(new_n553), .B(KEYINPUT74), .Z(G299));
  INV_X1    g129(.A(G168), .ZN(G286));
  NAND2_X1  g130(.A1(new_n529), .A2(G87), .ZN(new_n556));
  OAI21_X1  g131(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n518), .A2(G49), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(G288));
  INV_X1    g134(.A(G86), .ZN(new_n560));
  INV_X1    g135(.A(G48), .ZN(new_n561));
  OAI22_X1  g136(.A1(new_n522), .A2(new_n560), .B1(new_n537), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n509), .A2(G61), .ZN(new_n563));
  NAND2_X1  g138(.A1(G73), .A2(G543), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT75), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n514), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(G305));
  AND2_X1   g143(.A1(new_n509), .A2(G60), .ZN(new_n569));
  AND2_X1   g144(.A1(G72), .A2(G543), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT76), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n529), .A2(G85), .B1(new_n518), .B2(G47), .ZN(new_n574));
  AND2_X1   g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OR2_X1    g150(.A1(new_n571), .A2(new_n572), .ZN(new_n576));
  AND2_X1   g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(G290));
  NAND2_X1  g153(.A1(G301), .A2(G868), .ZN(new_n579));
  AND3_X1   g154(.A1(new_n509), .A2(new_n510), .A3(G92), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT77), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(KEYINPUT10), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n509), .A2(G66), .ZN(new_n583));
  NAND2_X1  g158(.A1(G79), .A2(G543), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n514), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n585), .B1(G54), .B2(new_n518), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n581), .A2(KEYINPUT10), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n579), .B1(new_n589), .B2(G868), .ZN(G284));
  OAI21_X1  g165(.A(new_n579), .B1(new_n589), .B2(G868), .ZN(G321));
  NAND2_X1  g166(.A1(G286), .A2(G868), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n553), .B(KEYINPUT74), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n593), .B2(G868), .ZN(G297));
  OAI21_X1  g169(.A(new_n592), .B1(new_n593), .B2(G868), .ZN(G280));
  INV_X1    g170(.A(G559), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n589), .B1(new_n596), .B2(G860), .ZN(G148));
  NOR2_X1   g172(.A1(new_n542), .A2(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n589), .A2(new_n596), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(G868), .ZN(new_n600));
  XOR2_X1   g175(.A(new_n600), .B(KEYINPUT78), .Z(G323));
  XNOR2_X1  g176(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g177(.A1(new_n472), .A2(new_n468), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT12), .ZN(new_n604));
  XNOR2_X1  g179(.A(KEYINPUT79), .B(KEYINPUT13), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n604), .B(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  OR2_X1    g182(.A1(new_n607), .A2(G2100), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n482), .A2(G135), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n471), .A2(G111), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n610), .A2(KEYINPUT80), .ZN(new_n611));
  OAI21_X1  g186(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n612), .B1(new_n610), .B2(KEYINPUT80), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n611), .A2(new_n613), .B1(new_n488), .B2(G123), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  OR2_X1    g190(.A1(new_n615), .A2(G2096), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n607), .A2(G2100), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n615), .A2(G2096), .ZN(new_n618));
  NAND4_X1  g193(.A1(new_n608), .A2(new_n616), .A3(new_n617), .A4(new_n618), .ZN(G156));
  INV_X1    g194(.A(KEYINPUT83), .ZN(new_n620));
  XNOR2_X1  g195(.A(G2427), .B(G2438), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2430), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT15), .B(G2435), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n624), .A2(KEYINPUT14), .A3(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT82), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G1341), .ZN(new_n629));
  INV_X1    g204(.A(G1348), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G2451), .B(G2454), .Z(new_n632));
  XNOR2_X1  g207(.A(G2443), .B(G2446), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n634), .B(new_n635), .Z(new_n636));
  NAND2_X1  g211(.A1(new_n629), .A2(new_n630), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n631), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(G14), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n636), .B1(new_n631), .B2(new_n637), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n620), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n631), .A2(new_n637), .ZN(new_n642));
  INV_X1    g217(.A(new_n636), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g219(.A1(new_n644), .A2(KEYINPUT83), .A3(G14), .A4(new_n638), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(G401));
  XOR2_X1   g222(.A(G2084), .B(G2090), .Z(new_n648));
  XNOR2_X1  g223(.A(G2067), .B(G2678), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2072), .B(G2078), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT18), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n651), .B(KEYINPUT17), .Z(new_n655));
  INV_X1    g230(.A(new_n648), .ZN(new_n656));
  INV_X1    g231(.A(new_n649), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n655), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n656), .A2(new_n652), .A3(new_n657), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(new_n650), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n654), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2096), .B(G2100), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(G227));
  XOR2_X1   g238(.A(G1971), .B(G1976), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1956), .B(G2474), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1961), .B(G1966), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AND2_X1   g243(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  NOR3_X1   g244(.A1(new_n665), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n665), .A2(new_n668), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT84), .B(KEYINPUT20), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  AOI211_X1 g248(.A(new_n670), .B(new_n673), .C1(new_n665), .C2(new_n669), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G1991), .B(G1996), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1981), .B(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(G229));
  OR2_X1    g255(.A1(G16), .A2(G23), .ZN(new_n681));
  NAND2_X1  g256(.A1(G288), .A2(KEYINPUT88), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT88), .ZN(new_n683));
  NAND4_X1  g258(.A1(new_n556), .A2(new_n558), .A3(new_n683), .A4(new_n557), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(G16), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n681), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT33), .B(G1976), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT89), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n689), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n686), .A2(G22), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT90), .Z(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(G166), .B2(new_n686), .ZN(new_n694));
  INV_X1    g269(.A(G1971), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(G6), .A2(G16), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(new_n567), .B2(G16), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT32), .B(G1981), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND4_X1  g275(.A1(new_n690), .A2(new_n691), .A3(new_n696), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT34), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n482), .A2(G131), .ZN(new_n703));
  NOR2_X1   g278(.A1(G95), .A2(G2105), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT85), .ZN(new_n705));
  INV_X1    g280(.A(G107), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n467), .B1(new_n706), .B2(G2105), .ZN(new_n707));
  AOI22_X1  g282(.A1(new_n705), .A2(new_n707), .B1(new_n488), .B2(G119), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n703), .A2(new_n708), .ZN(new_n709));
  MUX2_X1   g284(.A(G25), .B(new_n709), .S(G29), .Z(new_n710));
  XOR2_X1   g285(.A(KEYINPUT35), .B(G1991), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT86), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n710), .B(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n686), .A2(G24), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(new_n577), .B2(new_n686), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT87), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n713), .B1(new_n717), .B2(G1986), .ZN(new_n718));
  AOI211_X1 g293(.A(new_n702), .B(new_n718), .C1(G1986), .C2(new_n717), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT36), .ZN(new_n720));
  NOR2_X1   g295(.A1(G29), .A2(G35), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G162), .B2(G29), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT29), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(G2090), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n686), .A2(G20), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT23), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(new_n593), .B2(new_n686), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(G1956), .Z(new_n728));
  INV_X1    g303(.A(G29), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G26), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT92), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT28), .ZN(new_n732));
  OAI21_X1  g307(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n733));
  INV_X1    g308(.A(G116), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n733), .B1(new_n734), .B2(G2105), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(new_n488), .B2(G128), .ZN(new_n736));
  INV_X1    g311(.A(G140), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n481), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT91), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n732), .B1(new_n740), .B2(G29), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G2067), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n686), .A2(G5), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G171), .B2(new_n686), .ZN(new_n744));
  INV_X1    g319(.A(G1966), .ZN(new_n745));
  NOR2_X1   g320(.A1(G168), .A2(new_n686), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n686), .B2(G21), .ZN(new_n747));
  OAI22_X1  g322(.A1(new_n744), .A2(G1961), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G1961), .B2(new_n744), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n728), .A2(new_n742), .A3(new_n749), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT25), .Z(new_n752));
  AOI22_X1  g327(.A1(new_n472), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n753), .B2(new_n471), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n482), .B2(G139), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n755), .A2(new_n729), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n729), .B2(G33), .ZN(new_n757));
  INV_X1    g332(.A(G2072), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n488), .A2(G129), .ZN(new_n759));
  NAND3_X1  g334(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT26), .Z(new_n761));
  NAND2_X1  g336(.A1(new_n468), .A2(G105), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n759), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n482), .B2(G141), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n764), .A2(new_n729), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n729), .B2(G32), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT27), .B(G1996), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n757), .A2(new_n758), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n766), .B2(new_n767), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT93), .B(KEYINPUT24), .Z(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(G34), .ZN(new_n772));
  AOI21_X1  g347(.A(G29), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT94), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n773), .A2(KEYINPUT94), .B1(G34), .B2(new_n770), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n776), .A2(new_n777), .B1(G29), .B2(G160), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n778), .A2(G2084), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(G2084), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT30), .B(G28), .ZN(new_n781));
  OR2_X1    g356(.A1(KEYINPUT31), .A2(G11), .ZN(new_n782));
  NAND2_X1  g357(.A1(KEYINPUT31), .A2(G11), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n781), .A2(new_n729), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n780), .B(new_n784), .C1(new_n729), .C2(new_n615), .ZN(new_n785));
  NOR2_X1   g360(.A1(G16), .A2(G19), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n542), .B2(G16), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(G1341), .Z(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n757), .B2(new_n758), .ZN(new_n789));
  NOR4_X1   g364(.A1(new_n769), .A2(new_n779), .A3(new_n785), .A4(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(G27), .ZN(new_n791));
  OR3_X1    g366(.A1(new_n791), .A2(KEYINPUT96), .A3(G29), .ZN(new_n792));
  OAI21_X1  g367(.A(KEYINPUT96), .B1(new_n791), .B2(G29), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n792), .B(new_n793), .C1(G164), .C2(new_n729), .ZN(new_n794));
  INV_X1    g369(.A(G2078), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n686), .A2(G4), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n589), .B2(new_n686), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(new_n630), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n747), .A2(new_n745), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT95), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n790), .A2(new_n796), .A3(new_n799), .A4(new_n801), .ZN(new_n802));
  OR4_X1    g377(.A1(new_n720), .A2(new_n724), .A3(new_n750), .A4(new_n802), .ZN(G150));
  XNOR2_X1  g378(.A(G150), .B(KEYINPUT97), .ZN(G311));
  NAND2_X1  g379(.A1(new_n589), .A2(G559), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT38), .Z(new_n806));
  INV_X1    g381(.A(G93), .ZN(new_n807));
  INV_X1    g382(.A(G55), .ZN(new_n808));
  OAI22_X1  g383(.A1(new_n522), .A2(new_n807), .B1(new_n537), .B2(new_n808), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n810), .A2(new_n514), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n542), .B(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n806), .B(new_n813), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n814), .A2(KEYINPUT39), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n814), .A2(KEYINPUT39), .ZN(new_n816));
  NOR3_X1   g391(.A1(new_n815), .A2(new_n816), .A3(G860), .ZN(new_n817));
  OAI21_X1  g392(.A(G860), .B1(new_n809), .B2(new_n811), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT37), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n817), .A2(new_n819), .ZN(G145));
  XNOR2_X1  g395(.A(new_n615), .B(G160), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n490), .B(new_n821), .Z(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n739), .B(KEYINPUT98), .ZN(new_n824));
  AOI22_X1  g399(.A1(G126), .A2(new_n488), .B1(new_n498), .B2(new_n502), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n494), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n764), .B(new_n826), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n824), .A2(new_n827), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT99), .ZN(new_n830));
  OAI211_X1 g405(.A(new_n828), .B(new_n829), .C1(new_n830), .C2(new_n755), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n755), .A2(new_n830), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n488), .A2(G130), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n471), .A2(G118), .ZN(new_n835));
  OAI21_X1  g410(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(new_n482), .B2(G142), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(new_n604), .Z(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(new_n709), .Z(new_n840));
  NAND2_X1  g415(.A1(new_n833), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n833), .A2(new_n840), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n823), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n843), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n845), .A2(new_n822), .A3(new_n841), .ZN(new_n846));
  INV_X1    g421(.A(G37), .ZN(new_n847));
  AND3_X1   g422(.A1(new_n844), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(KEYINPUT40), .Z(G395));
  NOR2_X1   g424(.A1(new_n812), .A2(G868), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n599), .B(new_n813), .ZN(new_n851));
  NAND2_X1  g426(.A1(G299), .A2(new_n589), .ZN(new_n852));
  INV_X1    g427(.A(new_n589), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n593), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT41), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n852), .A2(new_n854), .A3(KEYINPUT41), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n857), .A2(KEYINPUT100), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n855), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT100), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n860), .A2(new_n861), .A3(KEYINPUT41), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n851), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n863), .B1(new_n851), .B2(new_n860), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n567), .B(G303), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n577), .B(new_n685), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n865), .B1(new_n866), .B2(KEYINPUT101), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(KEYINPUT101), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT42), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n864), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n864), .A2(new_n870), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n871), .A2(G868), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n850), .B1(new_n873), .B2(KEYINPUT102), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n874), .B1(KEYINPUT102), .B2(new_n873), .ZN(G295));
  OAI21_X1  g450(.A(new_n874), .B1(KEYINPUT102), .B2(new_n873), .ZN(G331));
  INV_X1    g451(.A(KEYINPUT44), .ZN(new_n877));
  XNOR2_X1  g452(.A(G301), .B(new_n813), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(G286), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n859), .A2(new_n862), .A3(new_n879), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n879), .A2(new_n860), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n869), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n847), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT103), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n880), .A2(new_n885), .A3(new_n881), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n869), .B1(new_n882), .B2(KEYINPUT103), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n884), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT43), .ZN(new_n889));
  OAI21_X1  g464(.A(KEYINPUT104), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n882), .A2(KEYINPUT103), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n891), .A2(new_n883), .A3(new_n886), .ZN(new_n892));
  INV_X1    g467(.A(new_n884), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT104), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n894), .A2(new_n895), .A3(KEYINPUT43), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n857), .A2(new_n897), .A3(new_n858), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n879), .B1(new_n857), .B2(new_n897), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n881), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n883), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n893), .A2(new_n889), .A3(new_n901), .ZN(new_n902));
  AND4_X1   g477(.A1(new_n877), .A2(new_n890), .A3(new_n896), .A4(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n892), .A2(new_n893), .A3(new_n889), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n893), .A2(new_n901), .ZN(new_n905));
  AOI22_X1  g480(.A1(new_n904), .A2(KEYINPUT106), .B1(new_n905), .B2(KEYINPUT43), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT106), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n888), .A2(new_n907), .A3(new_n889), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n877), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n903), .A2(new_n909), .ZN(G397));
  INV_X1    g485(.A(G1384), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT4), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n493), .B(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n497), .ZN(new_n914));
  AOI21_X1  g489(.A(KEYINPUT70), .B1(new_n914), .B2(new_n501), .ZN(new_n915));
  NOR3_X1   g490(.A1(new_n496), .A2(new_n497), .A3(new_n495), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n504), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n911), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(G40), .ZN(new_n919));
  NOR3_X1   g494(.A1(new_n470), .A2(new_n475), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT45), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n918), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT107), .ZN(new_n923));
  OR2_X1    g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n923), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n739), .B(G2067), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n764), .B(G1996), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n929), .A2(new_n703), .A3(new_n708), .A4(new_n711), .ZN(new_n930));
  INV_X1    g505(.A(G2067), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n739), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n926), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n709), .B(new_n711), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n926), .B1(new_n929), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(G1986), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n577), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT108), .ZN(new_n938));
  INV_X1    g513(.A(new_n926), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT48), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n935), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n938), .A2(KEYINPUT48), .A3(new_n939), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n933), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT47), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n926), .B1(new_n927), .B2(new_n764), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n945), .B(KEYINPUT123), .ZN(new_n946));
  INV_X1    g521(.A(G1996), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n939), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(KEYINPUT46), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n943), .B1(new_n944), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n951), .B1(new_n944), .B2(new_n950), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT54), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT50), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n954), .B1(new_n507), .B2(new_n911), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n920), .B1(new_n918), .B2(KEYINPUT50), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT116), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT116), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n473), .A2(new_n474), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(G2105), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n960), .A2(G40), .A3(new_n469), .A4(new_n466), .ZN(new_n961));
  AOI21_X1  g536(.A(G1384), .B1(new_n494), .B2(new_n825), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n961), .B1(new_n962), .B2(new_n954), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT71), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n917), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n503), .A2(KEYINPUT71), .A3(new_n504), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(G1384), .B1(new_n967), .B2(new_n494), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n958), .B(new_n963), .C1(new_n968), .C2(new_n954), .ZN(new_n969));
  INV_X1    g544(.A(G1961), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n957), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n961), .B1(new_n918), .B2(new_n921), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n962), .A2(KEYINPUT45), .ZN(new_n973));
  OR2_X1    g548(.A1(new_n795), .A2(KEYINPUT120), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT53), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n975), .B1(KEYINPUT120), .B2(new_n795), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n972), .A2(new_n973), .A3(new_n974), .A4(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT110), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT45), .B1(new_n507), .B2(new_n911), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n920), .B1(new_n918), .B2(new_n921), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n978), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n961), .B1(new_n962), .B2(KEYINPUT45), .ZN(new_n982));
  OAI211_X1 g557(.A(KEYINPUT110), .B(new_n982), .C1(new_n968), .C2(KEYINPUT45), .ZN(new_n983));
  AOI21_X1  g558(.A(G2078), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n971), .B(new_n977), .C1(new_n984), .C2(KEYINPUT53), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n953), .B1(new_n985), .B2(G171), .ZN(new_n986));
  OR2_X1    g561(.A1(new_n984), .A2(KEYINPUT53), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT119), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n507), .A2(KEYINPUT45), .A3(new_n911), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n989), .A2(new_n972), .A3(KEYINPUT53), .A4(new_n795), .ZN(new_n990));
  AND3_X1   g565(.A1(new_n971), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n988), .B1(new_n971), .B2(new_n990), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n987), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n986), .B1(new_n993), .B2(G171), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT51), .ZN(new_n995));
  INV_X1    g570(.A(G8), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n955), .A2(new_n956), .A3(G2084), .ZN(new_n999));
  AOI21_X1  g574(.A(G1966), .B1(new_n989), .B2(new_n972), .ZN(new_n1000));
  OAI21_X1  g575(.A(G168), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n989), .A2(new_n972), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n745), .ZN(new_n1003));
  INV_X1    g578(.A(G2084), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n1004), .B(new_n963), .C1(new_n968), .C2(new_n954), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1003), .A2(G286), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n998), .B1(new_n1001), .B2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1003), .A2(G168), .A3(new_n1005), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT51), .B1(new_n1008), .B2(G8), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n509), .A2(G62), .ZN(new_n1011));
  NAND2_X1  g586(.A1(G75), .A2(G543), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n514), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n511), .A2(new_n512), .ZN(new_n1014));
  OAI211_X1 g589(.A(KEYINPUT55), .B(G8), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT111), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g592(.A1(G303), .A2(KEYINPUT111), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n1017), .A2(KEYINPUT112), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT112), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1021));
  NOR3_X1   g596(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n981), .A2(new_n983), .A3(new_n695), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n961), .B1(new_n918), .B2(KEYINPUT50), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n507), .A2(new_n911), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1025), .B1(new_n1026), .B2(KEYINPUT50), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1024), .B1(G2090), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1023), .B1(new_n1028), .B2(G8), .ZN(new_n1029));
  OR3_X1    g604(.A1(new_n955), .A2(new_n956), .A3(G2090), .ZN(new_n1030));
  AOI211_X1 g605(.A(new_n996), .B(new_n1022), .C1(new_n1024), .C2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n682), .A2(G1976), .A3(new_n684), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n996), .B1(new_n962), .B2(new_n920), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT52), .ZN(new_n1035));
  OR3_X1    g610(.A1(new_n562), .A2(new_n566), .A3(G1981), .ZN(new_n1036));
  OAI21_X1  g611(.A(G1981), .B1(new_n562), .B2(new_n566), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT49), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1036), .A2(KEYINPUT49), .A3(new_n1037), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(new_n1033), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(G1976), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT52), .B1(G288), .B2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1032), .A2(new_n1033), .A3(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1035), .A2(new_n1042), .A3(new_n1045), .ZN(new_n1046));
  NOR3_X1   g621(.A1(new_n1029), .A2(new_n1031), .A3(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n994), .A2(new_n1010), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n993), .A2(G171), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n985), .A2(G171), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT54), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(KEYINPUT121), .B1(new_n1048), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n971), .A2(new_n990), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT119), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n971), .A2(new_n988), .A3(new_n990), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(G301), .B1(new_n1057), .B2(new_n987), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n953), .B1(new_n1058), .B2(new_n1050), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT121), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1028), .A2(G8), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(new_n1022), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n996), .B1(new_n1024), .B2(new_n1030), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1046), .B1(new_n1063), .B2(new_n1023), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1062), .A2(new_n1010), .A3(new_n1064), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1059), .A2(new_n1060), .A3(new_n994), .A4(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT57), .ZN(new_n1067));
  XNOR2_X1  g642(.A(new_n553), .B(new_n1067), .ZN(new_n1068));
  XOR2_X1   g643(.A(KEYINPUT115), .B(G1956), .Z(new_n1069));
  NAND2_X1  g644(.A1(new_n1027), .A2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n982), .B1(new_n968), .B2(KEYINPUT45), .ZN(new_n1071));
  XOR2_X1   g646(.A(KEYINPUT56), .B(G2072), .Z(new_n1072));
  OAI211_X1 g647(.A(new_n1068), .B(new_n1070), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n553), .B(KEYINPUT57), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n1027), .A2(new_n1069), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1074), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n957), .A2(new_n969), .A3(new_n630), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n918), .A2(new_n961), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n931), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n853), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1073), .B1(new_n1078), .B2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1079), .A2(KEYINPUT60), .A3(new_n1081), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1084), .A2(new_n589), .ZN(new_n1085));
  XNOR2_X1  g660(.A(KEYINPUT58), .B(G1341), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1080), .A2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n979), .A2(new_n980), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1087), .B1(new_n1088), .B2(new_n947), .ZN(new_n1089));
  INV_X1    g664(.A(new_n542), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1091), .A2(KEYINPUT59), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT59), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n1089), .A2(new_n1093), .A3(new_n1090), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1085), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1077), .A2(new_n1073), .A3(KEYINPUT61), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1096), .A2(KEYINPUT118), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1096), .A2(KEYINPUT118), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1095), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT60), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1102), .A2(new_n589), .A3(new_n1084), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT117), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1077), .A2(new_n1073), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT61), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1104), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  AOI211_X1 g682(.A(KEYINPUT117), .B(KEYINPUT61), .C1(new_n1077), .C2(new_n1073), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1103), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1083), .B1(new_n1099), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1053), .A2(new_n1066), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT113), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1046), .A2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1035), .A2(new_n1042), .A3(KEYINPUT113), .A4(new_n1045), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(G288), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1042), .A2(new_n1043), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n1036), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1031), .A2(new_n1115), .B1(new_n1033), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1001), .A2(new_n1006), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n997), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1008), .A2(G8), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(new_n995), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1121), .A2(new_n1123), .A3(KEYINPUT62), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT62), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1124), .A2(new_n1126), .A3(new_n993), .A4(G171), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1119), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1001), .A2(new_n996), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1115), .A2(KEYINPUT63), .A3(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1063), .A2(new_n1023), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n1131), .A2(new_n1031), .A3(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1062), .A2(new_n1064), .A3(new_n1130), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT63), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1133), .B1(new_n1136), .B2(KEYINPUT114), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT114), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1134), .A2(new_n1138), .A3(new_n1135), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1129), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1111), .A2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n577), .A2(new_n936), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n938), .A2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1143), .A2(new_n926), .ZN(new_n1144));
  OR2_X1    g719(.A1(new_n1144), .A2(new_n935), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1145), .B(KEYINPUT109), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(KEYINPUT122), .B1(new_n1141), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT122), .ZN(new_n1149));
  AOI211_X1 g724(.A(new_n1149), .B(new_n1146), .C1(new_n1111), .C2(new_n1140), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n952), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT124), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g728(.A(KEYINPUT124), .B(new_n952), .C1(new_n1148), .C2(new_n1150), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g730(.A(KEYINPUT127), .ZN(new_n1157));
  NOR2_X1   g731(.A1(G227), .A2(new_n460), .ZN(new_n1158));
  XOR2_X1   g732(.A(new_n1158), .B(KEYINPUT125), .Z(new_n1159));
  AOI21_X1  g733(.A(new_n1159), .B1(new_n641), .B2(new_n645), .ZN(new_n1160));
  INV_X1    g734(.A(KEYINPUT126), .ZN(new_n1161));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g736(.A(G229), .ZN(new_n1163));
  NAND2_X1  g737(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g738(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1165));
  OAI21_X1  g739(.A(new_n1157), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g740(.A(G229), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1167));
  OAI211_X1 g741(.A(new_n1167), .B(KEYINPUT127), .C1(new_n1161), .C2(new_n1160), .ZN(new_n1168));
  AOI21_X1  g742(.A(new_n848), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g743(.A1(new_n890), .A2(new_n896), .A3(new_n902), .ZN(new_n1170));
  AND2_X1   g744(.A1(new_n1169), .A2(new_n1170), .ZN(G308));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(G225));
endmodule


