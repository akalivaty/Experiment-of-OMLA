//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 1 0 0 0 0 1 1 1 0 0 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n574, new_n576, new_n577, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n631, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  XOR2_X1   g007(.A(KEYINPUT66), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XNOR2_X1  g015(.A(KEYINPUT67), .B(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT68), .Z(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  AOI22_X1  g035(.A1(new_n460), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n460), .A2(new_n462), .ZN(new_n464));
  INV_X1    g039(.A(G137), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(KEYINPUT69), .B1(new_n466), .B2(G2105), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT69), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(new_n462), .A3(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G101), .ZN(new_n471));
  OAI22_X1  g046(.A1(new_n464), .A2(new_n465), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n463), .A2(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(new_n460), .A2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(G124), .ZN(new_n475));
  OR3_X1    g050(.A1(new_n474), .A2(KEYINPUT70), .A3(new_n475), .ZN(new_n476));
  OAI21_X1  g051(.A(KEYINPUT70), .B1(new_n474), .B2(new_n475), .ZN(new_n477));
  INV_X1    g052(.A(new_n464), .ZN(new_n478));
  AOI22_X1  g053(.A1(new_n476), .A2(new_n477), .B1(G136), .B2(new_n478), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  NAND2_X1  g058(.A1(G114), .A2(G2104), .ZN(new_n484));
  AND2_X1   g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  NOR2_X1   g060(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(G126), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n484), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n466), .A2(G2105), .ZN(new_n490));
  AOI22_X1  g065(.A1(new_n489), .A2(G2105), .B1(G102), .B2(new_n490), .ZN(new_n491));
  OAI211_X1 g066(.A(G138), .B(new_n462), .C1(new_n485), .C2(new_n486), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n460), .A2(new_n494), .A3(G138), .A4(new_n462), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  INV_X1    g073(.A(G651), .ZN(new_n499));
  OAI21_X1  g074(.A(KEYINPUT72), .B1(new_n499), .B2(KEYINPUT6), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT72), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n501), .A2(new_n502), .A3(G651), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT71), .B(G651), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n500), .B(new_n503), .C1(new_n504), .C2(new_n502), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n505), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(G50), .A2(new_n507), .B1(new_n512), .B2(G88), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT73), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n512), .A2(G88), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n507), .A2(G50), .ZN(new_n517));
  AND3_X1   g092(.A1(new_n516), .A2(new_n517), .A3(new_n514), .ZN(new_n518));
  INV_X1    g093(.A(G62), .ZN(new_n519));
  OR3_X1    g094(.A1(new_n511), .A2(KEYINPUT74), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(G75), .A2(G543), .ZN(new_n521));
  OAI21_X1  g096(.A(KEYINPUT74), .B1(new_n511), .B2(new_n519), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g098(.A(KEYINPUT75), .B1(new_n523), .B2(new_n504), .ZN(new_n524));
  AND3_X1   g099(.A1(new_n523), .A2(KEYINPUT75), .A3(new_n504), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n515), .A2(new_n518), .B1(new_n524), .B2(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT76), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n509), .A2(G543), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n506), .A2(KEYINPUT5), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n508), .A2(new_n510), .A3(KEYINPUT76), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n535), .A2(G63), .A3(G651), .ZN(new_n536));
  NOR3_X1   g111(.A1(new_n499), .A2(KEYINPUT72), .A3(KEYINPUT6), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n499), .A2(KEYINPUT71), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT71), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G651), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n537), .B1(new_n541), .B2(KEYINPUT6), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n531), .A2(new_n532), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n542), .A2(G89), .A3(new_n543), .A4(new_n500), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n542), .A2(G51), .A3(G543), .A4(new_n500), .ZN(new_n545));
  AND4_X1   g120(.A1(new_n529), .A2(new_n536), .A3(new_n544), .A4(new_n545), .ZN(G168));
  INV_X1    g121(.A(KEYINPUT77), .ZN(new_n547));
  NAND4_X1  g122(.A1(new_n542), .A2(G52), .A3(G543), .A4(new_n500), .ZN(new_n548));
  NAND4_X1  g123(.A1(new_n542), .A2(G90), .A3(new_n543), .A4(new_n500), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AND3_X1   g125(.A1(new_n508), .A2(new_n510), .A3(KEYINPUT76), .ZN(new_n551));
  AOI21_X1  g126(.A(KEYINPUT76), .B1(new_n508), .B2(new_n510), .ZN(new_n552));
  OAI21_X1  g127(.A(G64), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(G77), .A2(G543), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n541), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n547), .B1(new_n550), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(G64), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n557), .B1(new_n533), .B2(new_n534), .ZN(new_n558));
  INV_X1    g133(.A(new_n554), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n504), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n560), .A2(KEYINPUT77), .A3(new_n548), .A4(new_n549), .ZN(new_n561));
  AND2_X1   g136(.A1(new_n556), .A2(new_n561), .ZN(G301));
  INV_X1    g137(.A(G301), .ZN(G171));
  NAND2_X1  g138(.A1(new_n507), .A2(G43), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n512), .A2(G81), .ZN(new_n565));
  INV_X1    g140(.A(G56), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n566), .B1(new_n533), .B2(new_n534), .ZN(new_n567));
  INV_X1    g142(.A(G68), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n568), .A2(new_n506), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n504), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n564), .A2(new_n565), .A3(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G860), .ZN(G153));
  AND3_X1   g148(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G36), .ZN(G176));
  NAND2_X1  g150(.A1(G1), .A2(G3), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT8), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n574), .A2(new_n577), .ZN(G188));
  INV_X1    g153(.A(KEYINPUT9), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n541), .A2(KEYINPUT6), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n580), .A2(G543), .A3(new_n500), .A4(new_n503), .ZN(new_n581));
  INV_X1    g156(.A(G53), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n579), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n512), .A2(G91), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n502), .B1(new_n538), .B2(new_n540), .ZN(new_n585));
  INV_X1    g160(.A(new_n500), .ZN(new_n586));
  NOR3_X1   g161(.A1(new_n585), .A2(new_n586), .A3(new_n537), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n587), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n588));
  NAND2_X1  g163(.A1(G78), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G65), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n511), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(G651), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n583), .A2(new_n584), .A3(new_n588), .A4(new_n592), .ZN(G299));
  INV_X1    g168(.A(G168), .ZN(G286));
  NAND2_X1  g169(.A1(new_n507), .A2(G49), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n512), .A2(G87), .ZN(new_n596));
  OAI21_X1  g171(.A(G651), .B1(new_n535), .B2(G74), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(G288));
  NAND3_X1  g173(.A1(new_n543), .A2(KEYINPUT78), .A3(G61), .ZN(new_n599));
  NAND2_X1  g174(.A1(G73), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT78), .ZN(new_n601));
  INV_X1    g176(.A(G61), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n511), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n599), .A2(new_n600), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(new_n504), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n512), .A2(G86), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n507), .A2(G48), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(G305));
  AOI22_X1  g183(.A1(new_n535), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n609), .A2(new_n541), .ZN(new_n610));
  INV_X1    g185(.A(G47), .ZN(new_n611));
  NAND4_X1  g186(.A1(new_n580), .A2(new_n543), .A3(new_n500), .A4(new_n503), .ZN(new_n612));
  XNOR2_X1  g187(.A(KEYINPUT79), .B(G85), .ZN(new_n613));
  OAI22_X1  g188(.A1(new_n611), .A2(new_n581), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(G290));
  NAND2_X1  g191(.A1(new_n507), .A2(G54), .ZN(new_n617));
  NAND2_X1  g192(.A1(G79), .A2(G543), .ZN(new_n618));
  INV_X1    g193(.A(G66), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n511), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G651), .ZN(new_n621));
  AOI21_X1  g196(.A(KEYINPUT10), .B1(new_n512), .B2(G92), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT10), .ZN(new_n623));
  INV_X1    g198(.A(G92), .ZN(new_n624));
  NOR4_X1   g199(.A1(new_n505), .A2(new_n623), .A3(new_n624), .A4(new_n511), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n617), .B(new_n621), .C1(new_n622), .C2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(G868), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(G171), .B2(new_n627), .ZN(G284));
  OAI21_X1  g204(.A(new_n628), .B1(G171), .B2(new_n627), .ZN(G321));
  NAND2_X1  g205(.A1(G299), .A2(new_n627), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(new_n627), .B2(G168), .ZN(G297));
  XOR2_X1   g207(.A(G297), .B(KEYINPUT80), .Z(G280));
  INV_X1    g208(.A(new_n626), .ZN(new_n634));
  INV_X1    g209(.A(G559), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n634), .B1(new_n635), .B2(G860), .ZN(G148));
  NAND3_X1  g211(.A1(new_n634), .A2(KEYINPUT81), .A3(new_n635), .ZN(new_n637));
  INV_X1    g212(.A(KEYINPUT81), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(new_n626), .B2(G559), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n627), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n572), .A2(G868), .ZN(new_n641));
  OAI21_X1  g216(.A(KEYINPUT82), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(KEYINPUT82), .B2(new_n640), .ZN(G323));
  XNOR2_X1  g218(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g219(.A(KEYINPUT83), .B(KEYINPUT12), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(new_n470), .B2(new_n487), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT83), .B(KEYINPUT12), .Z(new_n647));
  NAND4_X1  g222(.A1(new_n647), .A2(new_n460), .A3(new_n467), .A4(new_n469), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT13), .Z(new_n650));
  NAND2_X1  g225(.A1(KEYINPUT84), .A2(G2100), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n478), .A2(G135), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n460), .A2(G123), .A3(G2105), .ZN(new_n654));
  OR2_X1    g229(.A1(G99), .A2(G2105), .ZN(new_n655));
  OAI211_X1 g230(.A(new_n655), .B(G2104), .C1(G111), .C2(new_n462), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n653), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(G2096), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  OAI211_X1 g234(.A(new_n652), .B(new_n659), .C1(KEYINPUT84), .C2(G2100), .ZN(G156));
  XNOR2_X1  g235(.A(G2451), .B(G2454), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT16), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2443), .B(G2446), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1341), .B(G1348), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n664), .B(new_n665), .Z(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT15), .B(G2430), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G2435), .ZN(new_n668));
  XOR2_X1   g243(.A(G2427), .B(G2438), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(KEYINPUT14), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n666), .B(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(G14), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(G401));
  XNOR2_X1  g249(.A(G2072), .B(G2078), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT17), .Z(new_n676));
  XOR2_X1   g251(.A(G2067), .B(G2678), .Z(new_n677));
  XOR2_X1   g252(.A(G2084), .B(G2090), .Z(new_n678));
  NAND3_X1  g253(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT85), .Z(new_n680));
  NOR2_X1   g255(.A1(new_n676), .A2(new_n677), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n681), .A2(new_n678), .ZN(new_n682));
  INV_X1    g257(.A(new_n677), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n682), .B1(new_n683), .B2(new_n675), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n683), .A2(new_n675), .A3(new_n678), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT18), .Z(new_n686));
  NAND3_X1  g261(.A1(new_n680), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(new_n658), .ZN(new_n688));
  INV_X1    g263(.A(G2100), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(G227));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1971), .B(G1976), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT86), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT19), .ZN(new_n696));
  XOR2_X1   g271(.A(G1956), .B(G2474), .Z(new_n697));
  XOR2_X1   g272(.A(G1961), .B(G1966), .Z(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n696), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(KEYINPUT20), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n697), .A2(new_n698), .ZN(new_n703));
  OR3_X1    g278(.A1(new_n696), .A2(new_n700), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n696), .A2(new_n700), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT20), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n696), .A2(new_n703), .ZN(new_n708));
  NAND4_X1  g283(.A1(new_n702), .A2(new_n704), .A3(new_n707), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(G1991), .B(G1996), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  XOR2_X1   g287(.A(G1981), .B(G1986), .Z(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n701), .A2(KEYINPUT20), .B1(new_n696), .B2(new_n703), .ZN(new_n715));
  NAND4_X1  g290(.A1(new_n715), .A2(new_n710), .A3(new_n704), .A4(new_n707), .ZN(new_n716));
  AND3_X1   g291(.A1(new_n712), .A2(new_n714), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n714), .B1(new_n712), .B2(new_n716), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n693), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n712), .A2(new_n716), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(new_n713), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n712), .A2(new_n714), .A3(new_n716), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n721), .A2(new_n692), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n719), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(G229));
  XNOR2_X1  g300(.A(KEYINPUT87), .B(G29), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n727), .A2(KEYINPUT28), .A3(G26), .ZN(new_n728));
  OAI211_X1 g303(.A(G140), .B(new_n462), .C1(new_n485), .C2(new_n486), .ZN(new_n729));
  OAI211_X1 g304(.A(G128), .B(G2105), .C1(new_n485), .C2(new_n486), .ZN(new_n730));
  INV_X1    g305(.A(G116), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G2105), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n732), .B(G2104), .C1(G104), .C2(G2105), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n729), .A2(new_n730), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(KEYINPUT93), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT93), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n729), .A2(new_n730), .A3(new_n733), .A4(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G29), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n728), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(KEYINPUT28), .B1(new_n727), .B2(G26), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G2067), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n727), .A2(G35), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n482), .B2(new_n726), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT29), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G2090), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n727), .A2(G27), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G164), .B2(new_n727), .ZN(new_n751));
  INV_X1    g326(.A(G2078), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G160), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT24), .B(G34), .Z(new_n755));
  OAI22_X1  g330(.A1(new_n754), .A2(new_n740), .B1(new_n726), .B2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(G2084), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n740), .A2(G33), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n490), .A2(KEYINPUT25), .A3(G103), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT25), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(G127), .B1(new_n485), .B2(new_n486), .ZN(new_n766));
  NAND2_X1  g341(.A1(G115), .A2(G2104), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n462), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI211_X1 g343(.A(G139), .B(new_n462), .C1(new_n485), .C2(new_n486), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  NOR3_X1   g345(.A1(new_n765), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n759), .B1(new_n771), .B2(new_n740), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G2072), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n758), .A2(new_n773), .ZN(new_n774));
  AND4_X1   g349(.A1(new_n744), .A2(new_n749), .A3(new_n753), .A4(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n748), .A2(G2090), .ZN(new_n776));
  OAI21_X1  g351(.A(KEYINPUT90), .B1(G4), .B2(G16), .ZN(new_n777));
  OR3_X1    g352(.A1(KEYINPUT90), .A2(G4), .A3(G16), .ZN(new_n778));
  INV_X1    g353(.A(G16), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n777), .B(new_n778), .C1(new_n626), .C2(new_n779), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT91), .B(G1348), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n780), .A2(new_n782), .ZN(new_n784));
  NOR3_X1   g359(.A1(new_n776), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n779), .A2(G20), .ZN(new_n786));
  AND4_X1   g361(.A1(new_n584), .A2(new_n583), .A3(new_n588), .A4(new_n592), .ZN(new_n787));
  OAI211_X1 g362(.A(KEYINPUT23), .B(new_n786), .C1(new_n787), .C2(new_n779), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(KEYINPUT23), .B2(new_n786), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G1956), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n775), .A2(new_n785), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n779), .A2(G21), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G168), .B2(new_n779), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G1966), .ZN(new_n794));
  INV_X1    g369(.A(G28), .ZN(new_n795));
  AOI21_X1  g370(.A(G29), .B1(new_n795), .B2(KEYINPUT30), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(KEYINPUT30), .B2(new_n795), .ZN(new_n797));
  OR2_X1    g372(.A1(G29), .A2(G32), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n460), .A2(G141), .A3(new_n462), .ZN(new_n799));
  NAND3_X1  g374(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT26), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n460), .A2(G129), .A3(G2105), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n467), .A2(new_n469), .A3(G105), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n799), .A2(new_n802), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n798), .B1(new_n805), .B2(new_n740), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT27), .B(G1996), .ZN(new_n807));
  OAI221_X1 g382(.A(new_n797), .B1(new_n657), .B2(new_n727), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n806), .B2(new_n807), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n779), .A2(G19), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n572), .B2(new_n779), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT92), .B(G1341), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n809), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(new_n811), .B2(new_n812), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT31), .B(G11), .ZN(new_n815));
  OAI21_X1  g390(.A(KEYINPUT94), .B1(G5), .B2(G16), .ZN(new_n816));
  OR3_X1    g391(.A1(KEYINPUT94), .A2(G5), .A3(G16), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n816), .B(new_n817), .C1(G301), .C2(new_n779), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT95), .B(G1961), .Z(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n818), .A2(new_n819), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n814), .A2(new_n815), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  NOR3_X1   g397(.A1(new_n791), .A2(new_n794), .A3(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT96), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT34), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n779), .A2(G23), .ZN(new_n826));
  AND3_X1   g401(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n827), .B2(new_n779), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT33), .Z(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(G1976), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n779), .A2(G22), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(G166), .B2(new_n779), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(G1971), .ZN(new_n833));
  INV_X1    g408(.A(G1971), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n834), .B(new_n831), .C1(G166), .C2(new_n779), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n779), .A2(G6), .ZN(new_n836));
  INV_X1    g411(.A(G305), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n836), .B1(new_n837), .B2(new_n779), .ZN(new_n838));
  XOR2_X1   g413(.A(KEYINPUT32), .B(G1981), .Z(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n833), .A2(new_n835), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n825), .B1(new_n830), .B2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(G1976), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n829), .B(new_n843), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n833), .A2(new_n840), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n844), .A2(KEYINPUT34), .A3(new_n835), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n842), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n727), .A2(G25), .ZN(new_n848));
  OR2_X1    g423(.A1(G95), .A2(G2105), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n849), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n850));
  OAI211_X1 g425(.A(G131), .B(new_n462), .C1(new_n485), .C2(new_n486), .ZN(new_n851));
  OAI211_X1 g426(.A(G119), .B(G2105), .C1(new_n485), .C2(new_n486), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n848), .B1(new_n854), .B2(new_n727), .ZN(new_n855));
  XNOR2_X1  g430(.A(KEYINPUT35), .B(G1991), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n855), .B(new_n857), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n615), .B(KEYINPUT88), .Z(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(G16), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(G16), .B2(G24), .ZN(new_n861));
  INV_X1    g436(.A(G1986), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n847), .A2(new_n858), .A3(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT89), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n866), .A2(KEYINPUT36), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n863), .B1(new_n842), .B2(new_n846), .ZN(new_n869));
  INV_X1    g444(.A(new_n867), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n869), .A2(new_n870), .A3(new_n858), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n866), .A2(KEYINPUT36), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n824), .B1(new_n872), .B2(new_n873), .ZN(G311));
  INV_X1    g449(.A(new_n871), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n870), .B1(new_n869), .B2(new_n858), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n873), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n824), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(G150));
  NAND2_X1  g454(.A1(G80), .A2(G543), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n881), .B1(new_n535), .B2(G67), .ZN(new_n882));
  OAI21_X1  g457(.A(KEYINPUT97), .B1(new_n882), .B2(new_n541), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n542), .A2(G55), .A3(G543), .A4(new_n500), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n542), .A2(G93), .A3(new_n543), .A4(new_n500), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(G67), .B1(new_n551), .B2(new_n552), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n880), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT97), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n888), .A2(new_n889), .A3(new_n504), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n883), .A2(new_n886), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(G860), .ZN(new_n892));
  XOR2_X1   g467(.A(new_n892), .B(KEYINPUT37), .Z(new_n893));
  NOR2_X1   g468(.A1(new_n626), .A2(new_n635), .ZN(new_n894));
  XNOR2_X1  g469(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n894), .B(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n889), .B1(new_n888), .B2(new_n504), .ZN(new_n897));
  AOI211_X1 g472(.A(KEYINPUT97), .B(new_n541), .C1(new_n887), .C2(new_n880), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT98), .ZN(new_n900));
  INV_X1    g475(.A(G43), .ZN(new_n901));
  INV_X1    g476(.A(G81), .ZN(new_n902));
  OAI22_X1  g477(.A1(new_n901), .A2(new_n581), .B1(new_n612), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(G56), .B1(new_n551), .B2(new_n552), .ZN(new_n904));
  INV_X1    g479(.A(new_n569), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n541), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n900), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n564), .A2(new_n565), .A3(new_n570), .A4(KEYINPUT98), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n899), .A2(new_n907), .A3(new_n908), .A4(new_n886), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n891), .A2(new_n900), .A3(new_n571), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n896), .B(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n893), .B1(new_n912), .B2(G860), .ZN(G145));
  XNOR2_X1  g488(.A(new_n482), .B(new_n754), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(new_n657), .ZN(new_n915));
  AOI22_X1  g490(.A1(new_n460), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n769), .B(new_n764), .C1(new_n916), .C2(new_n462), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n917), .A2(new_n491), .A3(new_n496), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n917), .B1(new_n491), .B2(new_n496), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n735), .A2(new_n805), .A3(new_n737), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n805), .B1(new_n735), .B2(new_n737), .ZN(new_n922));
  OAI22_X1  g497(.A1(new_n919), .A2(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n460), .A2(G130), .A3(G2105), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT99), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT99), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n460), .A2(new_n926), .A3(G130), .A4(G2105), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n929));
  OR2_X1    g504(.A1(new_n929), .A2(KEYINPUT100), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(KEYINPUT100), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n930), .B(new_n931), .C1(G118), .C2(new_n462), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n478), .A2(G142), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n928), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n853), .A2(new_n646), .A3(new_n648), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n853), .B1(new_n646), .B2(new_n648), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n649), .A2(new_n854), .ZN(new_n939));
  AOI22_X1  g514(.A1(new_n925), .A2(new_n927), .B1(new_n478), .B2(G142), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n939), .A2(new_n940), .A3(new_n932), .A4(new_n935), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n497), .A2(new_n771), .ZN(new_n943));
  INV_X1    g518(.A(new_n805), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n738), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n735), .A2(new_n805), .A3(new_n737), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n943), .A2(new_n945), .A3(new_n918), .A4(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n923), .A2(new_n942), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT101), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT101), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n923), .A2(new_n942), .A3(new_n947), .A4(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n949), .A2(KEYINPUT102), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n923), .A2(new_n947), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n953), .A2(new_n941), .A3(new_n938), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT102), .B1(new_n949), .B2(new_n951), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n915), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT103), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT103), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n959), .B(new_n915), .C1(new_n955), .C2(new_n956), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n657), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n914), .B(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n949), .A2(new_n951), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n963), .A2(new_n954), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G37), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n961), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT104), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n961), .A2(KEYINPUT104), .A3(new_n968), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n973), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g549(.A(KEYINPUT42), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n637), .A2(new_n639), .ZN(new_n976));
  OR2_X1    g551(.A1(new_n976), .A2(new_n911), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n911), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n787), .A2(new_n626), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n623), .B1(new_n612), .B2(new_n624), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n587), .A2(KEYINPUT10), .A3(G92), .A4(new_n543), .ZN(new_n982));
  AOI22_X1  g557(.A1(new_n981), .A2(new_n982), .B1(G651), .B2(new_n620), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n983), .A2(G299), .A3(new_n617), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n980), .A2(KEYINPUT105), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT105), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n634), .A2(new_n986), .A3(G299), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n979), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT41), .B1(new_n980), .B2(new_n984), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n992), .B1(new_n988), .B2(KEYINPUT41), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n979), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n975), .B1(new_n991), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(G303), .A2(new_n837), .ZN(new_n996));
  OAI221_X1 g571(.A(G305), .B1(new_n524), .B2(new_n525), .C1(new_n515), .C2(new_n518), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n827), .B1(new_n610), .B2(new_n614), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT106), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n615), .A2(G288), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n999), .B1(new_n998), .B2(new_n1000), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n996), .B(new_n997), .C1(new_n1002), .C2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n996), .A2(new_n997), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n1001), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n1008), .A2(KEYINPUT107), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n990), .B(KEYINPUT42), .C1(new_n979), .C2(new_n993), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n995), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1009), .B1(new_n995), .B2(new_n1010), .ZN(new_n1012));
  OAI21_X1  g587(.A(G868), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n891), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1013), .B1(G868), .B2(new_n1014), .ZN(G295));
  OAI21_X1  g590(.A(new_n1013), .B1(G868), .B2(new_n1014), .ZN(G331));
  AND3_X1   g591(.A1(new_n556), .A2(G168), .A3(new_n561), .ZN(new_n1017));
  AOI21_X1  g592(.A(G168), .B1(new_n556), .B2(new_n561), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(new_n911), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n909), .B(new_n910), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n989), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1020), .A2(KEYINPUT108), .A3(new_n1021), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT108), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1019), .A2(new_n911), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1022), .B1(new_n1026), .B2(new_n993), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT109), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1004), .A2(new_n1006), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1029), .B(new_n1022), .C1(new_n1026), .C2(new_n993), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1031), .A2(new_n966), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT43), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1007), .B(new_n1022), .C1(new_n1026), .C2(new_n993), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n1036), .A2(new_n966), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT41), .ZN(new_n1038));
  AOI22_X1  g613(.A1(new_n1020), .A2(new_n1021), .B1(new_n988), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n980), .A2(new_n984), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(KEYINPUT41), .ZN(new_n1041));
  AOI22_X1  g616(.A1(new_n1026), .A2(new_n989), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT110), .B1(new_n1042), .B2(new_n1007), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT110), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n988), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1044), .B(new_n1008), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1037), .A2(new_n1043), .A3(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1035), .B1(new_n1048), .B2(new_n1034), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT44), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1037), .A2(new_n1043), .A3(new_n1047), .A4(new_n1034), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1033), .A2(KEYINPUT43), .ZN(new_n1052));
  AND2_X1   g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1050), .B1(KEYINPUT44), .B2(new_n1053), .ZN(G397));
  INV_X1    g629(.A(G1384), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n497), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT45), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(G160), .A2(G40), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(G1384), .B1(new_n491), .B2(new_n496), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT45), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1058), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g638(.A(KEYINPUT56), .B(G2072), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g640(.A(G299), .B(KEYINPUT57), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  OR2_X1    g642(.A1(new_n1061), .A2(KEYINPUT50), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1061), .A2(KEYINPUT50), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1059), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1065), .B(new_n1067), .C1(G1956), .C2(new_n1070), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1061), .A2(KEYINPUT50), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1061), .A2(KEYINPUT50), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1060), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G2067), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n1074), .A2(new_n782), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1077), .A2(new_n626), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT118), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1058), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1064), .ZN(new_n1081));
  OAI22_X1  g656(.A1(new_n1070), .A2(G1956), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(new_n1066), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1079), .A2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1078), .A2(KEYINPUT118), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1071), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT120), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1088));
  OAI22_X1  g663(.A1(new_n1070), .A2(new_n781), .B1(G2067), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT60), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1087), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1077), .A2(KEYINPUT120), .A3(KEYINPUT60), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1091), .A2(new_n634), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1087), .B(new_n626), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1071), .A2(new_n1083), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT61), .ZN(new_n1098));
  XOR2_X1   g673(.A(KEYINPUT58), .B(G1341), .Z(new_n1099));
  NAND2_X1  g674(.A1(new_n1088), .A2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1100), .B1(new_n1080), .B2(G1996), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT119), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT119), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1100), .B(new_n1103), .C1(new_n1080), .C2(G1996), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1102), .A2(new_n572), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT59), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1097), .A2(new_n1098), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  OR2_X1    g682(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1096), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1086), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1063), .A2(KEYINPUT53), .A3(new_n752), .ZN(new_n1112));
  INV_X1    g687(.A(G1961), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1074), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT53), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(new_n1080), .B2(G2078), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1112), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(G171), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1112), .A2(G301), .A3(new_n1116), .A4(new_n1114), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1118), .A2(KEYINPUT123), .A3(new_n1119), .ZN(new_n1120));
  OR2_X1    g695(.A1(new_n1119), .A2(KEYINPUT123), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(G8), .ZN(new_n1124));
  NOR2_X1   g699(.A1(G168), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT122), .ZN(new_n1126));
  OAI21_X1  g701(.A(KEYINPUT51), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(G1966), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n1070), .A2(new_n757), .B1(new_n1080), .B2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1129), .A2(new_n1124), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1127), .B1(new_n1130), .B2(new_n1125), .ZN(new_n1131));
  OAI22_X1  g706(.A1(new_n1063), .A2(G1966), .B1(new_n1074), .B2(G2084), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(G8), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1125), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1133), .A2(new_n1126), .A3(KEYINPUT51), .A4(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1136), .B1(new_n1129), .B2(new_n1134), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1132), .A2(KEYINPUT121), .A3(new_n1125), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1131), .A2(new_n1135), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1123), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT52), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1076), .A2(new_n1124), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n827), .A2(G1976), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1142), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1143), .ZN(new_n1146));
  NAND2_X1  g721(.A1(G305), .A2(G1981), .ZN(new_n1147));
  INV_X1    g722(.A(G1981), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n605), .A2(new_n606), .A3(new_n607), .A4(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1147), .A2(KEYINPUT49), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(KEYINPUT115), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT115), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1147), .A2(new_n1152), .A3(KEYINPUT49), .A4(new_n1149), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1146), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1155));
  XNOR2_X1  g730(.A(KEYINPUT114), .B(KEYINPUT49), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1145), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g733(.A(KEYINPUT113), .B(G1976), .ZN(new_n1159));
  AOI21_X1  g734(.A(KEYINPUT52), .B1(G288), .B2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1143), .A2(new_n1144), .A3(new_n1160), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n1158), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(G2090), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1070), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1080), .A2(new_n834), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1124), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1167));
  AND3_X1   g742(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1166), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1168), .A2(new_n1167), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT117), .ZN(new_n1171));
  AOI21_X1  g746(.A(G2090), .B1(new_n1074), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1070), .A2(KEYINPUT117), .ZN(new_n1173));
  AOI22_X1  g748(.A1(new_n1172), .A2(new_n1173), .B1(new_n834), .B2(new_n1080), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1170), .B1(new_n1174), .B2(new_n1124), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1118), .A2(KEYINPUT54), .A3(new_n1119), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1162), .A2(new_n1169), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1141), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1111), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1180), .A2(new_n843), .A3(new_n827), .ZN(new_n1181));
  XOR2_X1   g756(.A(new_n1149), .B(KEYINPUT116), .Z(new_n1182));
  AOI21_X1  g757(.A(new_n1146), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1175), .A2(new_n1169), .A3(new_n1158), .A4(new_n1161), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1184), .B1(KEYINPUT62), .B2(new_n1140), .ZN(new_n1185));
  AND3_X1   g760(.A1(new_n1131), .A2(new_n1135), .A3(new_n1139), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT62), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1118), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1183), .B1(new_n1185), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(new_n1170), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1162), .A2(new_n1190), .A3(new_n1166), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1130), .A2(G168), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1184), .A2(new_n1192), .ZN(new_n1193));
  OR2_X1    g768(.A1(new_n1190), .A2(new_n1166), .ZN(new_n1194));
  NAND4_X1  g769(.A1(new_n1162), .A2(new_n1194), .A3(KEYINPUT63), .A4(new_n1169), .ZN(new_n1195));
  OAI22_X1  g770(.A1(new_n1193), .A2(KEYINPUT63), .B1(new_n1195), .B2(new_n1192), .ZN(new_n1196));
  NAND4_X1  g771(.A1(new_n1179), .A2(new_n1189), .A3(new_n1191), .A4(new_n1196), .ZN(new_n1197));
  NOR2_X1   g772(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1198), .A2(G1996), .A3(new_n805), .ZN(new_n1199));
  XNOR2_X1  g774(.A(new_n1199), .B(KEYINPUT111), .ZN(new_n1200));
  INV_X1    g775(.A(new_n1198), .ZN(new_n1201));
  OR2_X1    g776(.A1(new_n1201), .A2(G1996), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1202), .A2(new_n805), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n1200), .A2(new_n1203), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n738), .B(G2067), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1198), .A2(new_n1205), .ZN(new_n1206));
  XNOR2_X1  g781(.A(new_n1206), .B(KEYINPUT112), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1204), .A2(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n853), .B(new_n856), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1208), .B1(new_n1198), .B2(new_n1209), .ZN(new_n1210));
  XNOR2_X1  g785(.A(new_n615), .B(new_n862), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1211), .A2(new_n1198), .ZN(new_n1212));
  AND2_X1   g787(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1197), .A2(new_n1213), .ZN(new_n1214));
  NAND4_X1  g789(.A1(new_n1204), .A2(new_n857), .A3(new_n854), .A4(new_n1207), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n739), .A2(new_n1075), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1201), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(KEYINPUT124), .A2(KEYINPUT46), .ZN(new_n1218));
  XNOR2_X1  g793(.A(new_n1202), .B(new_n1218), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1198), .B1(new_n805), .B2(new_n1205), .ZN(new_n1220));
  OAI21_X1  g795(.A(new_n1220), .B1(KEYINPUT124), .B2(KEYINPUT46), .ZN(new_n1221));
  NOR2_X1   g796(.A1(new_n1219), .A2(new_n1221), .ZN(new_n1222));
  XNOR2_X1  g797(.A(KEYINPUT125), .B(KEYINPUT47), .ZN(new_n1223));
  XNOR2_X1  g798(.A(new_n1222), .B(new_n1223), .ZN(new_n1224));
  NAND3_X1  g799(.A1(new_n1198), .A2(new_n862), .A3(new_n615), .ZN(new_n1225));
  XNOR2_X1  g800(.A(new_n1225), .B(KEYINPUT48), .ZN(new_n1226));
  AOI211_X1 g801(.A(new_n1217), .B(new_n1224), .C1(new_n1210), .C2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1214), .A2(new_n1227), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g803(.A(KEYINPUT126), .ZN(new_n1230));
  NAND4_X1  g804(.A1(new_n724), .A2(G319), .A3(new_n673), .A4(new_n690), .ZN(new_n1231));
  INV_X1    g805(.A(new_n1231), .ZN(new_n1232));
  AOI21_X1  g806(.A(KEYINPUT104), .B1(new_n961), .B2(new_n968), .ZN(new_n1233));
  AOI211_X1 g807(.A(new_n970), .B(new_n967), .C1(new_n958), .C2(new_n960), .ZN(new_n1234));
  OAI21_X1  g808(.A(new_n1232), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  OAI21_X1  g809(.A(new_n1230), .B1(new_n1053), .B2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g810(.A(new_n1231), .B1(new_n971), .B2(new_n972), .ZN(new_n1237));
  NAND2_X1  g811(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1238));
  NAND3_X1  g812(.A1(new_n1237), .A2(KEYINPUT126), .A3(new_n1238), .ZN(new_n1239));
  NAND2_X1  g813(.A1(new_n1236), .A2(new_n1239), .ZN(G308));
  NAND2_X1  g814(.A1(new_n1237), .A2(new_n1238), .ZN(G225));
endmodule


