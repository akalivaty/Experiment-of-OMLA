//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 0 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n795, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003;
  INV_X1    g000(.A(G120gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G113gat), .ZN(new_n203));
  INV_X1    g002(.A(G113gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G120gat), .ZN(new_n205));
  AOI21_X1  g004(.A(KEYINPUT1), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G127gat), .B(G134gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(KEYINPUT71), .A2(G127gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(KEYINPUT71), .A2(G127gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n210), .A2(G134gat), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT72), .ZN(new_n213));
  AND2_X1   g012(.A1(KEYINPUT71), .A2(G127gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(KEYINPUT71), .A2(G127gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT72), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(new_n217), .A3(G134gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT70), .ZN(new_n219));
  INV_X1    g018(.A(G127gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n219), .B1(new_n220), .B2(G134gat), .ZN(new_n221));
  INV_X1    g020(.A(G134gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n222), .A2(KEYINPUT70), .A3(G127gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n213), .A2(new_n218), .A3(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n206), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n209), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT24), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n228), .B(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(G183gat), .A2(G190gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(G169gat), .A2(G176gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT67), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n233), .B(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT25), .ZN(new_n236));
  NOR2_X1   g035(.A1(G169gat), .A2(G176gat), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n236), .B1(new_n237), .B2(KEYINPUT23), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n240), .B1(new_n237), .B2(KEYINPUT23), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT23), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n242), .B(KEYINPUT65), .C1(G169gat), .C2(G176gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NOR3_X1   g044(.A1(new_n232), .A2(new_n239), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n230), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n231), .B(KEYINPUT64), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n233), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n250), .B1(KEYINPUT23), .B2(new_n237), .ZN(new_n251));
  AND3_X1   g050(.A1(new_n244), .A2(KEYINPUT66), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT66), .B1(new_n244), .B2(new_n251), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n249), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n246), .B1(new_n254), .B2(new_n236), .ZN(new_n255));
  XNOR2_X1  g054(.A(KEYINPUT27), .B(G183gat), .ZN(new_n256));
  INV_X1    g055(.A(G190gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  XOR2_X1   g057(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT26), .ZN(new_n261));
  OAI21_X1  g060(.A(KEYINPUT69), .B1(new_n237), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n237), .A2(new_n261), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n264), .B(new_n233), .C1(new_n265), .C2(new_n263), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n260), .A2(new_n266), .A3(new_n228), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n227), .B1(new_n255), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n224), .B1(new_n212), .B2(KEYINPUT72), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n217), .B1(new_n216), .B2(G134gat), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n226), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(new_n208), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n244), .A2(new_n251), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT66), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n244), .A2(KEYINPUT66), .A3(new_n251), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT25), .B1(new_n278), .B2(new_n249), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n273), .B(new_n267), .C1(new_n279), .C2(new_n246), .ZN(new_n280));
  INV_X1    g079(.A(G227gat), .ZN(new_n281));
  INV_X1    g080(.A(G233gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n269), .A2(new_n280), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT32), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT33), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  XOR2_X1   g086(.A(G15gat), .B(G43gat), .Z(new_n288));
  XNOR2_X1  g087(.A(G71gat), .B(G99gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n285), .A2(new_n287), .A3(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n290), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n284), .B(KEYINPUT32), .C1(new_n286), .C2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n283), .B1(new_n269), .B2(new_n280), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT34), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI211_X1 g096(.A(KEYINPUT34), .B(new_n283), .C1(new_n269), .C2(new_n280), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT36), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n297), .A2(new_n298), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n302), .A2(new_n291), .A3(new_n293), .ZN(new_n303));
  AND3_X1   g102(.A1(new_n300), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n301), .B1(new_n300), .B2(new_n303), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT6), .ZN(new_n307));
  XNOR2_X1  g106(.A(G1gat), .B(G29gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n308), .B(KEYINPUT0), .ZN(new_n309));
  XNOR2_X1  g108(.A(G57gat), .B(G85gat), .ZN(new_n310));
  XOR2_X1   g109(.A(new_n309), .B(new_n310), .Z(new_n311));
  NAND2_X1  g110(.A1(G155gat), .A2(G162gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT2), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT78), .ZN(new_n314));
  NAND2_X1  g113(.A1(G141gat), .A2(G148gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(G141gat), .A2(G148gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT78), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n312), .A2(new_n319), .A3(KEYINPUT2), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n314), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  AND3_X1   g120(.A1(KEYINPUT77), .A2(G155gat), .A3(G162gat), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT77), .B1(G155gat), .B2(G162gat), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n322), .B1(new_n312), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n317), .ZN(new_n325));
  AND3_X1   g124(.A1(new_n325), .A2(new_n313), .A3(new_n315), .ZN(new_n326));
  XNOR2_X1  g125(.A(G155gat), .B(G162gat), .ZN(new_n327));
  AOI22_X1  g126(.A1(new_n321), .A2(new_n324), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n272), .A2(new_n328), .A3(new_n208), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT80), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT80), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n227), .A2(new_n331), .A3(new_n328), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT4), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n330), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G225gat), .A2(G233gat), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n329), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n336), .B1(new_n337), .B2(KEYINPUT4), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n324), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n326), .A2(new_n327), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT3), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT3), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n342), .A2(new_n273), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT79), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI22_X1  g146(.A1(new_n341), .A2(KEYINPUT3), .B1(new_n272), .B2(new_n208), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT79), .B1(new_n348), .B2(new_n344), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n334), .B(new_n338), .C1(new_n347), .C2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT5), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n273), .A2(new_n341), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n330), .A2(new_n332), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n351), .B1(new_n353), .B2(new_n336), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n350), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n345), .A2(new_n346), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n348), .A2(KEYINPUT79), .A3(new_n344), .ZN(new_n357));
  AOI22_X1  g156(.A1(new_n356), .A2(new_n357), .B1(new_n333), .B2(new_n329), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n333), .B1(new_n330), .B2(new_n332), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n336), .A2(KEYINPUT5), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n358), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  AOI211_X1 g161(.A(new_n307), .B(new_n311), .C1(new_n355), .C2(new_n362), .ZN(new_n363));
  AND2_X1   g162(.A1(new_n355), .A2(new_n362), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT6), .B1(new_n364), .B2(new_n311), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n311), .B1(new_n355), .B2(new_n362), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n363), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(G226gat), .A2(G233gat), .ZN(new_n369));
  INV_X1    g168(.A(new_n246), .ZN(new_n370));
  AOI22_X1  g169(.A1(new_n276), .A2(new_n277), .B1(new_n247), .B2(new_n248), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n370), .B1(new_n371), .B2(KEYINPUT25), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n369), .B1(new_n372), .B2(new_n267), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT29), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n374), .B1(new_n255), .B2(new_n268), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n373), .B1(new_n375), .B2(new_n369), .ZN(new_n376));
  INV_X1    g175(.A(G204gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(G197gat), .ZN(new_n378));
  INV_X1    g177(.A(G197gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(G204gat), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT73), .ZN(new_n381));
  AND3_X1   g180(.A1(new_n378), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n381), .B1(new_n378), .B2(new_n380), .ZN(new_n383));
  INV_X1    g182(.A(G211gat), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT74), .ZN(new_n385));
  INV_X1    g184(.A(G218gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(KEYINPUT74), .A2(G218gat), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n384), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI22_X1  g188(.A1(new_n382), .A2(new_n383), .B1(new_n389), .B2(KEYINPUT22), .ZN(new_n390));
  XOR2_X1   g189(.A(G211gat), .B(G218gat), .Z(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n379), .A2(G204gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n377), .A2(G197gat), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT73), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n380), .A3(new_n381), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n388), .ZN(new_n398));
  NOR2_X1   g197(.A1(KEYINPUT74), .A2(G218gat), .ZN(new_n399));
  OAI21_X1  g198(.A(G211gat), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT22), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n391), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n397), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n392), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n376), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(KEYINPUT75), .B(KEYINPUT29), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n408), .B1(new_n255), .B2(new_n268), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n369), .ZN(new_n410));
  INV_X1    g209(.A(new_n369), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n411), .B1(new_n255), .B2(new_n268), .ZN(new_n412));
  AOI211_X1 g211(.A(KEYINPUT76), .B(new_n405), .C1(new_n410), .C2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT76), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n407), .B1(new_n372), .B2(new_n267), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n412), .B1(new_n415), .B2(new_n411), .ZN(new_n416));
  INV_X1    g215(.A(new_n405), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n414), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n406), .B1(new_n413), .B2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(G8gat), .B(G36gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(G64gat), .B(G92gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n420), .B(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n422), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n406), .B(new_n424), .C1(new_n413), .C2(new_n418), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n423), .A2(KEYINPUT30), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n373), .B1(new_n369), .B2(new_n409), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT76), .B1(new_n427), .B2(new_n405), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n416), .A2(new_n414), .A3(new_n417), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT30), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n430), .A2(new_n431), .A3(new_n406), .A4(new_n424), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n368), .B1(new_n426), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT82), .ZN(new_n434));
  NAND2_X1  g233(.A1(G228gat), .A2(G233gat), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n407), .B1(new_n392), .B2(new_n404), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n341), .B1(new_n437), .B2(KEYINPUT3), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n344), .A2(new_n408), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n417), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n436), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n390), .A2(new_n391), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n403), .B1(new_n397), .B2(new_n402), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n374), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n328), .B1(new_n444), .B2(new_n343), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n407), .B1(new_n328), .B2(new_n343), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n436), .B1(new_n446), .B2(new_n405), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n434), .B(G22gat), .C1(new_n441), .C2(new_n448), .ZN(new_n449));
  XNOR2_X1  g248(.A(G78gat), .B(G106gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(KEYINPUT31), .B(G50gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n450), .B(new_n451), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(G22gat), .B1(new_n441), .B2(new_n448), .ZN(new_n454));
  NOR3_X1   g253(.A1(new_n441), .A2(new_n448), .A3(G22gat), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n454), .B1(new_n455), .B2(KEYINPUT82), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n452), .ZN(new_n458));
  INV_X1    g257(.A(G22gat), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n408), .B1(new_n442), .B2(new_n443), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n328), .B1(new_n460), .B2(new_n343), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n446), .A2(new_n405), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n435), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT29), .B1(new_n392), .B2(new_n404), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n341), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n465), .A2(new_n440), .A3(new_n436), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n459), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n458), .B1(new_n455), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT81), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n463), .A2(new_n459), .A3(new_n466), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n452), .B1(new_n454), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT81), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n457), .A2(new_n470), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT83), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n457), .A2(new_n470), .A3(KEYINPUT83), .A4(new_n473), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n306), .B1(new_n433), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n363), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n355), .A2(new_n362), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT85), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n355), .A2(new_n362), .A3(KEYINPUT85), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n311), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n311), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n307), .B1(new_n481), .B2(new_n486), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n480), .B(new_n425), .C1(new_n485), .C2(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(KEYINPUT87), .B(KEYINPUT37), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n430), .A2(new_n406), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT37), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n492), .B1(new_n376), .B2(new_n417), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n416), .A2(new_n405), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT38), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AND3_X1   g294(.A1(new_n491), .A2(new_n495), .A3(new_n422), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n488), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n491), .A2(new_n422), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n492), .B1(new_n430), .B2(new_n406), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT38), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n497), .A2(new_n500), .B1(new_n476), .B2(new_n477), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT40), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n335), .B1(new_n358), .B2(new_n360), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT39), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  OR2_X1    g305(.A1(new_n353), .A2(new_n336), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT39), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n311), .B1(new_n503), .B2(new_n508), .ZN(new_n509));
  OAI211_X1 g308(.A(KEYINPUT84), .B(new_n502), .C1(new_n506), .C2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n484), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT85), .B1(new_n355), .B2(new_n362), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n486), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n503), .A2(new_n508), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n502), .A2(KEYINPUT84), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n514), .A2(new_n311), .A3(new_n505), .A4(new_n515), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n510), .A2(new_n513), .A3(new_n516), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n517), .A2(KEYINPUT86), .A3(new_n426), .A4(new_n432), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT86), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n425), .A2(KEYINPUT30), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n424), .B1(new_n430), .B2(new_n406), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n432), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n510), .A2(new_n513), .A3(new_n516), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n519), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n479), .B1(new_n501), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT89), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n300), .A2(new_n303), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n527), .B1(new_n478), .B2(new_n529), .ZN(new_n530));
  AOI211_X1 g329(.A(KEYINPUT89), .B(new_n528), .C1(new_n476), .C2(new_n477), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n433), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(KEYINPUT35), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT88), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n472), .A2(KEYINPUT81), .ZN(new_n535));
  AOI211_X1 g334(.A(new_n469), .B(new_n452), .C1(new_n454), .C2(new_n471), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT83), .B1(new_n537), .B2(new_n457), .ZN(new_n538));
  AND4_X1   g337(.A1(KEYINPUT83), .A2(new_n457), .A3(new_n470), .A4(new_n473), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n529), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT35), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n480), .B1(new_n485), .B2(new_n487), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n522), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n534), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n542), .A2(new_n541), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n528), .B1(new_n476), .B2(new_n477), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n545), .A2(new_n546), .A3(KEYINPUT88), .A4(new_n522), .ZN(new_n547));
  AND2_X1   g346(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n526), .B1(new_n533), .B2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G113gat), .B(G141gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT11), .ZN(new_n551));
  INV_X1    g350(.A(G169gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(G197gat), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n554), .B(KEYINPUT12), .Z(new_n555));
  INV_X1    g354(.A(KEYINPUT90), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n556), .A2(G8gat), .ZN(new_n557));
  XOR2_X1   g356(.A(G15gat), .B(G22gat), .Z(new_n558));
  INV_X1    g357(.A(G1gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(G15gat), .B(G22gat), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT16), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n561), .B1(new_n562), .B2(G1gat), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n557), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n556), .A2(G8gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G43gat), .B(G50gat), .ZN(new_n568));
  OR3_X1    g367(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n569));
  OAI21_X1  g368(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n570));
  AOI22_X1  g369(.A1(new_n569), .A2(new_n570), .B1(G29gat), .B2(G36gat), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n568), .B1(new_n571), .B2(KEYINPUT15), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(KEYINPUT15), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n567), .A2(new_n574), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n572), .B(new_n573), .Z(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(new_n566), .ZN(new_n577));
  NAND2_X1  g376(.A1(G229gat), .A2(G233gat), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n578), .B(KEYINPUT13), .Z(new_n579));
  NAND3_X1  g378(.A1(new_n575), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT92), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n574), .A2(KEYINPUT17), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT91), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n566), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(KEYINPUT17), .B1(new_n567), .B2(KEYINPUT91), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n584), .B1(new_n585), .B2(new_n576), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n586), .A2(KEYINPUT18), .A3(new_n578), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT18), .B1(new_n586), .B2(new_n578), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n555), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n589), .ZN(new_n591));
  INV_X1    g390(.A(new_n555), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n591), .A2(new_n581), .A3(new_n587), .A4(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n549), .A2(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(G183gat), .B(G211gat), .Z(new_n597));
  XNOR2_X1  g396(.A(G57gat), .B(G64gat), .ZN(new_n598));
  AOI21_X1  g397(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n599));
  OR2_X1    g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(G71gat), .B(G78gat), .Z(new_n601));
  OR2_X1    g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n601), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT21), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(G231gat), .A2(G233gat), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n606), .B(new_n607), .Z(new_n608));
  XOR2_X1   g407(.A(G127gat), .B(G155gat), .Z(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT20), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n608), .B(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT94), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n604), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n567), .B1(KEYINPUT21), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  OR2_X1    g417(.A1(new_n608), .A2(new_n610), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n608), .A2(new_n610), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n619), .A2(new_n613), .A3(new_n620), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n615), .A2(new_n618), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n618), .B1(new_n615), .B2(new_n621), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n597), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n615), .A2(new_n621), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(new_n617), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n615), .A2(new_n618), .A3(new_n621), .ZN(new_n627));
  INV_X1    g426(.A(new_n597), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G85gat), .A2(G92gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT7), .ZN(new_n632));
  INV_X1    g431(.A(G99gat), .ZN(new_n633));
  INV_X1    g432(.A(G106gat), .ZN(new_n634));
  OAI21_X1  g433(.A(KEYINPUT8), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI211_X1 g434(.A(new_n632), .B(new_n635), .C1(G85gat), .C2(G92gat), .ZN(new_n636));
  XOR2_X1   g435(.A(G99gat), .B(G106gat), .Z(new_n637));
  OR2_X1    g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT97), .ZN(new_n641));
  AND2_X1   g440(.A1(new_n574), .A2(KEYINPUT17), .ZN(new_n642));
  OR3_X1    g441(.A1(new_n641), .A2(new_n582), .A3(new_n642), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n638), .A2(new_n639), .ZN(new_n644));
  AND2_X1   g443(.A1(G232gat), .A2(G233gat), .ZN(new_n645));
  AOI22_X1  g444(.A1(new_n576), .A2(new_n644), .B1(KEYINPUT41), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(G190gat), .B(G218gat), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n648), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n643), .A2(new_n646), .A3(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n645), .A2(KEYINPUT41), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT95), .ZN(new_n653));
  XNOR2_X1  g452(.A(G134gat), .B(G162gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n649), .A2(new_n651), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT98), .ZN(new_n658));
  OR2_X1    g457(.A1(new_n651), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n651), .A2(new_n658), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n659), .A2(new_n660), .A3(new_n649), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n655), .B(KEYINPUT96), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n657), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n630), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(G230gat), .A2(G233gat), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(KEYINPUT99), .Z(new_n666));
  NAND2_X1  g465(.A1(new_n644), .A2(new_n616), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT10), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n640), .A2(new_n604), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n644), .A2(KEYINPUT10), .A3(new_n616), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n666), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n666), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n673), .B1(new_n667), .B2(new_n669), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(G120gat), .B(G148gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(G176gat), .B(G204gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  OR3_X1    g478(.A1(new_n672), .A2(new_n674), .A3(new_n678), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n679), .A2(KEYINPUT100), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT100), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n675), .A2(new_n682), .A3(new_n678), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n664), .A2(new_n685), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n596), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n368), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(G1gat), .ZN(G1324gat));
  INV_X1    g488(.A(new_n522), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT16), .B(G8gat), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OR2_X1    g492(.A1(new_n693), .A2(KEYINPUT42), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(KEYINPUT42), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n691), .A2(G8gat), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n696), .A2(KEYINPUT101), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n696), .A2(KEYINPUT101), .ZN(new_n698));
  OAI211_X1 g497(.A(new_n694), .B(new_n695), .C1(new_n697), .C2(new_n698), .ZN(G1325gat));
  AOI21_X1  g498(.A(G15gat), .B1(new_n687), .B2(new_n529), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT102), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  INV_X1    g502(.A(new_n306), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n687), .A2(G15gat), .A3(new_n704), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(G1326gat));
  INV_X1    g505(.A(new_n478), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n687), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT43), .B(G22gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1327gat));
  NOR3_X1   g509(.A1(new_n630), .A2(new_n663), .A3(new_n685), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n596), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(G29gat), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n368), .A2(new_n713), .ZN(new_n714));
  OR3_X1    g513(.A1(new_n712), .A2(KEYINPUT103), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(KEYINPUT103), .B1(new_n712), .B2(new_n714), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n715), .A2(KEYINPUT45), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(KEYINPUT45), .B1(new_n715), .B2(new_n716), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n720));
  INV_X1    g519(.A(new_n433), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n540), .A2(KEYINPUT89), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n546), .A2(new_n527), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n544), .B(new_n547), .C1(new_n724), .C2(new_n541), .ZN(new_n725));
  INV_X1    g524(.A(new_n526), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n663), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n720), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  OAI211_X1 g528(.A(KEYINPUT105), .B(KEYINPUT44), .C1(new_n549), .C2(new_n663), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n727), .A2(new_n728), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n630), .A2(new_n685), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n594), .A2(KEYINPUT104), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT104), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n590), .A2(new_n593), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n734), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n733), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n368), .ZN(new_n743));
  OAI21_X1  g542(.A(G29gat), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n719), .A2(new_n744), .ZN(G1328gat));
  INV_X1    g544(.A(G36gat), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n690), .A2(new_n746), .ZN(new_n747));
  OR2_X1    g546(.A1(new_n712), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT106), .ZN(new_n749));
  OR3_X1    g548(.A1(new_n748), .A2(new_n749), .A3(KEYINPUT46), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(new_n748), .B2(KEYINPUT46), .ZN(new_n751));
  AOI22_X1  g550(.A1(new_n750), .A2(new_n751), .B1(KEYINPUT46), .B2(new_n748), .ZN(new_n752));
  OAI21_X1  g551(.A(G36gat), .B1(new_n742), .B2(new_n522), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(G1329gat));
  INV_X1    g553(.A(G43gat), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n755), .B1(new_n712), .B2(new_n528), .ZN(new_n756));
  XOR2_X1   g555(.A(KEYINPUT107), .B(KEYINPUT47), .Z(new_n757));
  NOR2_X1   g556(.A1(new_n306), .A2(new_n755), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n756), .B(new_n757), .C1(new_n742), .C2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT47), .ZN(new_n761));
  INV_X1    g560(.A(new_n756), .ZN(new_n762));
  AOI22_X1  g561(.A1(new_n729), .A2(new_n730), .B1(new_n728), .B2(new_n727), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n763), .A2(new_n740), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n762), .B1(new_n764), .B2(new_n758), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n760), .B1(new_n761), .B2(new_n765), .ZN(G1330gat));
  INV_X1    g565(.A(G50gat), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n596), .A2(new_n767), .A3(new_n707), .A4(new_n711), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n763), .A2(new_n478), .A3(new_n740), .ZN(new_n769));
  OAI211_X1 g568(.A(KEYINPUT48), .B(new_n768), .C1(new_n769), .C2(new_n767), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT108), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n768), .B(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n733), .A2(new_n707), .A3(new_n741), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n772), .B1(new_n773), .B2(G50gat), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n770), .B1(new_n774), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g574(.A1(new_n630), .A2(new_n663), .A3(new_n685), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n549), .A2(new_n739), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n368), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n690), .ZN(new_n780));
  NOR2_X1   g579(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n781));
  AND2_X1   g580(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n783), .B1(new_n781), .B2(new_n780), .ZN(G1333gat));
  NAND2_X1  g583(.A1(new_n777), .A2(new_n529), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT109), .ZN(new_n786));
  AOI21_X1  g585(.A(G71gat), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n787), .B1(new_n786), .B2(new_n785), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n777), .A2(G71gat), .A3(new_n704), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT50), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT50), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n788), .A2(new_n792), .A3(new_n789), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(G1334gat));
  NAND2_X1  g593(.A1(new_n777), .A2(new_n707), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(G78gat), .ZN(G1335gat));
  INV_X1    g595(.A(new_n663), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n624), .A2(new_n629), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n798), .A2(KEYINPUT110), .A3(new_n738), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT110), .B1(new_n798), .B2(new_n738), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n544), .A2(new_n547), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n803), .B1(KEYINPUT35), .B2(new_n532), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n797), .B(new_n802), .C1(new_n804), .C2(new_n526), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT51), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n727), .A2(KEYINPUT51), .A3(new_n802), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n684), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(G85gat), .B1(new_n809), .B2(new_n368), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n802), .A2(new_n685), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n811), .B1(new_n731), .B2(new_n732), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n368), .A2(G85gat), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n810), .B1(new_n812), .B2(new_n814), .ZN(G1336gat));
  INV_X1    g614(.A(G92gat), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n816), .B1(new_n812), .B2(new_n690), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT111), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n690), .A2(new_n816), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n818), .B1(new_n809), .B2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(KEYINPUT52), .B1(new_n817), .B2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n763), .A2(new_n522), .A3(new_n811), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n824), .B(new_n821), .C1(new_n825), .C2(new_n816), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n823), .A2(new_n826), .ZN(G1337gat));
  AOI21_X1  g626(.A(G99gat), .B1(new_n809), .B2(new_n529), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n306), .A2(new_n633), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n828), .B1(new_n812), .B2(new_n829), .ZN(G1338gat));
  AOI21_X1  g629(.A(new_n634), .B1(new_n812), .B2(new_n707), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n478), .A2(G106gat), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT51), .B1(new_n727), .B2(new_n802), .ZN(new_n833));
  NOR4_X1   g632(.A1(new_n549), .A2(new_n806), .A3(new_n663), .A4(new_n801), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n685), .B(new_n832), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(KEYINPUT112), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n807), .A2(new_n808), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT112), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n837), .A2(new_n838), .A3(new_n685), .A4(new_n832), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(KEYINPUT53), .B1(new_n831), .B2(new_n840), .ZN(new_n841));
  XNOR2_X1  g640(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n763), .A2(new_n478), .A3(new_n811), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n835), .B(new_n842), .C1(new_n843), .C2(new_n634), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n841), .A2(new_n844), .ZN(G1339gat));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n672), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n670), .A2(new_n671), .A3(new_n666), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n678), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n850), .B1(new_n672), .B2(new_n846), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT55), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n849), .A2(KEYINPUT55), .A3(new_n851), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n854), .A2(new_n680), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n856), .A2(new_n735), .A3(new_n737), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n575), .A2(new_n577), .ZN(new_n858));
  OAI22_X1  g657(.A1(new_n586), .A2(new_n578), .B1(new_n858), .B2(new_n579), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n554), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n593), .A2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n685), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n797), .B1(new_n857), .B2(new_n863), .ZN(new_n864));
  AND3_X1   g663(.A1(new_n797), .A2(new_n856), .A3(new_n862), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n798), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n686), .A2(new_n738), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n540), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n690), .A2(new_n743), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n870), .A2(new_n204), .A3(new_n595), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n743), .B1(new_n866), .B2(new_n867), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n722), .A2(new_n723), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n874), .A2(new_n690), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n739), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n871), .B1(new_n876), .B2(new_n204), .ZN(G1340gat));
  NOR3_X1   g676(.A1(new_n870), .A2(new_n202), .A3(new_n684), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n875), .A2(new_n685), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n878), .B1(new_n879), .B2(new_n202), .ZN(G1341gat));
  NAND3_X1  g679(.A1(new_n875), .A2(new_n216), .A3(new_n630), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n870), .A2(new_n798), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n881), .B1(new_n216), .B2(new_n882), .ZN(G1342gat));
  NAND2_X1  g682(.A1(new_n797), .A2(new_n522), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n884), .B(KEYINPUT114), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n874), .A2(G134gat), .A3(new_n885), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT56), .ZN(new_n887));
  OAI21_X1  g686(.A(G134gat), .B1(new_n870), .B2(new_n663), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(G1343gat));
  INV_X1    g688(.A(G141gat), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n869), .A2(new_n306), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT57), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n856), .A2(new_n594), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n797), .B1(new_n893), .B2(new_n863), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n798), .B1(new_n865), .B2(new_n894), .ZN(new_n895));
  AOI211_X1 g694(.A(new_n892), .B(new_n478), .C1(new_n895), .C2(new_n867), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n478), .B1(new_n866), .B2(new_n867), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n897), .A2(KEYINPUT57), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n896), .B1(new_n898), .B2(KEYINPUT115), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT115), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n900), .B1(new_n897), .B2(KEYINPUT57), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n891), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n890), .B1(new_n902), .B2(new_n739), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n707), .A2(new_n306), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(KEYINPUT116), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n595), .A2(G141gat), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n872), .A2(new_n522), .A3(new_n905), .A4(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(KEYINPUT58), .B1(new_n903), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n866), .A2(new_n867), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(new_n707), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(KEYINPUT115), .A3(new_n892), .ZN(new_n912));
  INV_X1    g711(.A(new_n896), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n912), .A2(new_n913), .A3(new_n901), .ZN(new_n914));
  INV_X1    g713(.A(new_n891), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n914), .A2(new_n594), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(G141gat), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n908), .A2(KEYINPUT117), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT117), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n907), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(KEYINPUT58), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  AND3_X1   g721(.A1(new_n917), .A2(new_n918), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n918), .B1(new_n917), .B2(new_n922), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n909), .B1(new_n923), .B2(new_n924), .ZN(G1344gat));
  NAND3_X1  g724(.A1(new_n872), .A2(new_n522), .A3(new_n905), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(G148gat), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n927), .A2(new_n928), .A3(new_n685), .ZN(new_n929));
  AOI211_X1 g728(.A(KEYINPUT59), .B(new_n928), .C1(new_n902), .C2(new_n685), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT59), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n893), .A2(new_n863), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n663), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n797), .A2(new_n856), .A3(new_n862), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n630), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n664), .A2(new_n594), .A3(new_n685), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n892), .B(new_n707), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n891), .A2(new_n684), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n937), .B(new_n938), .C1(new_n897), .C2(new_n892), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n931), .B1(new_n939), .B2(G148gat), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n929), .B1(new_n930), .B2(new_n940), .ZN(G1345gat));
  AOI21_X1  g740(.A(G155gat), .B1(new_n927), .B2(new_n630), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n630), .A2(G155gat), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT119), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n942), .B1(new_n902), .B2(new_n944), .ZN(G1346gat));
  NAND2_X1  g744(.A1(new_n902), .A2(new_n797), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(G162gat), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n872), .A2(new_n905), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n948), .A2(G162gat), .A3(new_n885), .ZN(new_n949));
  XOR2_X1   g748(.A(new_n949), .B(KEYINPUT120), .Z(new_n950));
  NAND2_X1  g749(.A1(new_n947), .A2(new_n950), .ZN(G1347gat));
  NAND2_X1  g750(.A1(new_n690), .A2(new_n743), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  AND3_X1   g752(.A1(new_n910), .A2(new_n873), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g753(.A(G169gat), .B1(new_n954), .B2(new_n739), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n868), .A2(new_n953), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n956), .A2(new_n552), .A3(new_n595), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n955), .A2(new_n957), .ZN(G1348gat));
  INV_X1    g757(.A(G176gat), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n954), .A2(new_n959), .A3(new_n685), .ZN(new_n960));
  OAI21_X1  g759(.A(G176gat), .B1(new_n956), .B2(new_n684), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(G1349gat));
  AND2_X1   g761(.A1(new_n630), .A2(new_n256), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n954), .A2(new_n963), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT60), .ZN(new_n965));
  OAI21_X1  g764(.A(KEYINPUT121), .B1(new_n956), .B2(new_n798), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(G183gat), .ZN(new_n967));
  NOR3_X1   g766(.A1(new_n956), .A2(KEYINPUT121), .A3(new_n798), .ZN(new_n968));
  OAI221_X1 g767(.A(new_n964), .B1(KEYINPUT122), .B2(new_n965), .C1(new_n967), .C2(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n965), .A2(KEYINPUT122), .ZN(new_n970));
  XNOR2_X1  g769(.A(new_n969), .B(new_n970), .ZN(G1350gat));
  OAI21_X1  g770(.A(G190gat), .B1(new_n956), .B2(new_n663), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT61), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n954), .A2(new_n257), .A3(new_n797), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n974), .ZN(G1351gat));
  NOR2_X1   g774(.A1(new_n952), .A2(new_n704), .ZN(new_n976));
  AND2_X1   g775(.A1(new_n897), .A2(new_n976), .ZN(new_n977));
  XOR2_X1   g776(.A(KEYINPUT123), .B(G197gat), .Z(new_n978));
  NOR2_X1   g777(.A1(new_n738), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g779(.A(new_n980), .B(KEYINPUT124), .ZN(new_n981));
  OAI211_X1 g780(.A(new_n937), .B(new_n976), .C1(new_n897), .C2(new_n892), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n978), .B1(new_n982), .B2(new_n595), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n981), .A2(new_n983), .ZN(G1352gat));
  NAND3_X1  g783(.A1(new_n977), .A2(new_n377), .A3(new_n685), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT62), .ZN(new_n986));
  XNOR2_X1  g785(.A(new_n985), .B(new_n986), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT125), .ZN(new_n988));
  OR3_X1    g787(.A1(new_n982), .A2(new_n988), .A3(new_n684), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n988), .B1(new_n982), .B2(new_n684), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n989), .A2(G204gat), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n987), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n992), .A2(KEYINPUT126), .ZN(new_n993));
  INV_X1    g792(.A(KEYINPUT126), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n987), .A2(new_n991), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n993), .A2(new_n995), .ZN(G1353gat));
  OAI21_X1  g795(.A(G211gat), .B1(new_n982), .B2(new_n798), .ZN(new_n997));
  XOR2_X1   g796(.A(new_n997), .B(KEYINPUT63), .Z(new_n998));
  NAND3_X1  g797(.A1(new_n977), .A2(new_n384), .A3(new_n630), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n998), .A2(new_n999), .ZN(G1354gat));
  AND2_X1   g799(.A1(new_n977), .A2(new_n797), .ZN(new_n1001));
  OAI21_X1  g800(.A(new_n797), .B1(new_n399), .B2(new_n398), .ZN(new_n1002));
  OAI22_X1  g801(.A1(new_n1001), .A2(G218gat), .B1(new_n982), .B2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g802(.A(new_n1003), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


