

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X1 U323 ( .A(n435), .B(KEYINPUT65), .ZN(n566) );
  AND2_X1 U324 ( .A1(n434), .A2(n550), .ZN(n435) );
  XNOR2_X1 U325 ( .A(KEYINPUT48), .B(n409), .ZN(n548) );
  XNOR2_X1 U326 ( .A(n301), .B(n300), .ZN(n312) );
  AND2_X1 U327 ( .A1(G232GAT), .A2(G233GAT), .ZN(n291) );
  XOR2_X1 U328 ( .A(G204GAT), .B(G64GAT), .Z(n292) );
  AND2_X1 U329 ( .A1(n568), .A2(n555), .ZN(n363) );
  XNOR2_X1 U330 ( .A(KEYINPUT113), .B(KEYINPUT47), .ZN(n400) );
  XNOR2_X1 U331 ( .A(KEYINPUT119), .B(KEYINPUT54), .ZN(n411) );
  XNOR2_X1 U332 ( .A(n388), .B(n291), .ZN(n389) );
  XNOR2_X1 U333 ( .A(n299), .B(n298), .ZN(n301) );
  XNOR2_X1 U334 ( .A(n390), .B(n389), .ZN(n394) );
  XOR2_X1 U335 ( .A(n559), .B(n402), .Z(n579) );
  XNOR2_X1 U336 ( .A(n312), .B(n311), .ZN(n572) );
  XOR2_X1 U337 ( .A(n398), .B(n397), .Z(n559) );
  XNOR2_X1 U338 ( .A(n459), .B(KEYINPUT122), .ZN(n460) );
  XNOR2_X1 U339 ( .A(n461), .B(n460), .ZN(G1351GAT) );
  XNOR2_X1 U340 ( .A(G71GAT), .B(G57GAT), .ZN(n293) );
  XNOR2_X1 U341 ( .A(n293), .B(KEYINPUT13), .ZN(n377) );
  XOR2_X1 U342 ( .A(G148GAT), .B(KEYINPUT76), .Z(n295) );
  XNOR2_X1 U343 ( .A(G106GAT), .B(G78GAT), .ZN(n294) );
  XNOR2_X1 U344 ( .A(n295), .B(n294), .ZN(n437) );
  XOR2_X1 U345 ( .A(n377), .B(n437), .Z(n299) );
  XOR2_X1 U346 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n297) );
  XNOR2_X1 U347 ( .A(G120GAT), .B(KEYINPUT79), .ZN(n296) );
  XOR2_X1 U348 ( .A(n297), .B(n296), .Z(n298) );
  XOR2_X1 U349 ( .A(G99GAT), .B(G85GAT), .Z(n383) );
  XOR2_X1 U350 ( .A(n383), .B(KEYINPUT31), .Z(n300) );
  XNOR2_X1 U351 ( .A(G176GAT), .B(G92GAT), .ZN(n302) );
  XNOR2_X1 U352 ( .A(n292), .B(n302), .ZN(n338) );
  INV_X1 U353 ( .A(KEYINPUT77), .ZN(n303) );
  XNOR2_X1 U354 ( .A(n338), .B(n303), .ZN(n307) );
  INV_X1 U355 ( .A(n307), .ZN(n305) );
  NAND2_X1 U356 ( .A1(G230GAT), .A2(G233GAT), .ZN(n306) );
  INV_X1 U357 ( .A(n306), .ZN(n304) );
  NAND2_X1 U358 ( .A1(n305), .A2(n304), .ZN(n309) );
  NAND2_X1 U359 ( .A1(n307), .A2(n306), .ZN(n308) );
  NAND2_X1 U360 ( .A1(n309), .A2(n308), .ZN(n310) );
  XNOR2_X1 U361 ( .A(n310), .B(KEYINPUT78), .ZN(n311) );
  XOR2_X1 U362 ( .A(KEYINPUT41), .B(KEYINPUT64), .Z(n313) );
  XNOR2_X1 U363 ( .A(n572), .B(n313), .ZN(n555) );
  XOR2_X1 U364 ( .A(KEYINPUT85), .B(KEYINPUT17), .Z(n315) );
  XNOR2_X1 U365 ( .A(KEYINPUT19), .B(G183GAT), .ZN(n314) );
  XNOR2_X1 U366 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U367 ( .A(KEYINPUT18), .B(n316), .ZN(n341) );
  XOR2_X1 U368 ( .A(KEYINPUT20), .B(KEYINPUT67), .Z(n318) );
  XNOR2_X1 U369 ( .A(G169GAT), .B(G71GAT), .ZN(n317) );
  XNOR2_X1 U370 ( .A(n318), .B(n317), .ZN(n330) );
  XOR2_X1 U371 ( .A(G15GAT), .B(G127GAT), .Z(n366) );
  XOR2_X1 U372 ( .A(G176GAT), .B(G190GAT), .Z(n320) );
  XNOR2_X1 U373 ( .A(G43GAT), .B(G99GAT), .ZN(n319) );
  XNOR2_X1 U374 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U375 ( .A(n366), .B(n321), .Z(n323) );
  NAND2_X1 U376 ( .A1(G227GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U377 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U378 ( .A(n324), .B(KEYINPUT86), .Z(n328) );
  XOR2_X1 U379 ( .A(KEYINPUT0), .B(G120GAT), .Z(n326) );
  XNOR2_X1 U380 ( .A(G113GAT), .B(G134GAT), .ZN(n325) );
  XNOR2_X1 U381 ( .A(n326), .B(n325), .ZN(n424) );
  XNOR2_X1 U382 ( .A(n424), .B(KEYINPUT84), .ZN(n327) );
  XNOR2_X1 U383 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U384 ( .A(n330), .B(n329), .Z(n331) );
  XOR2_X1 U385 ( .A(n341), .B(n331), .Z(n535) );
  INV_X1 U386 ( .A(n535), .ZN(n467) );
  XOR2_X1 U387 ( .A(G169GAT), .B(G8GAT), .Z(n346) );
  XOR2_X1 U388 ( .A(KEYINPUT92), .B(n346), .Z(n333) );
  NAND2_X1 U389 ( .A1(G226GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U390 ( .A(n333), .B(n332), .ZN(n336) );
  XOR2_X1 U391 ( .A(KEYINPUT21), .B(G211GAT), .Z(n335) );
  XNOR2_X1 U392 ( .A(G197GAT), .B(G218GAT), .ZN(n334) );
  XNOR2_X1 U393 ( .A(n335), .B(n334), .ZN(n441) );
  XOR2_X1 U394 ( .A(n336), .B(n441), .Z(n340) );
  XNOR2_X1 U395 ( .A(G36GAT), .B(G190GAT), .ZN(n337) );
  XNOR2_X1 U396 ( .A(n337), .B(KEYINPUT81), .ZN(n395) );
  XNOR2_X1 U397 ( .A(n395), .B(n338), .ZN(n339) );
  XNOR2_X1 U398 ( .A(n340), .B(n339), .ZN(n342) );
  XNOR2_X1 U399 ( .A(n342), .B(n341), .ZN(n524) );
  XNOR2_X1 U400 ( .A(KEYINPUT118), .B(n524), .ZN(n410) );
  XOR2_X1 U401 ( .A(G113GAT), .B(G22GAT), .Z(n344) );
  XNOR2_X1 U402 ( .A(G197GAT), .B(G15GAT), .ZN(n343) );
  XNOR2_X1 U403 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U404 ( .A(n345), .B(G36GAT), .Z(n348) );
  XNOR2_X1 U405 ( .A(n346), .B(G50GAT), .ZN(n347) );
  XNOR2_X1 U406 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U407 ( .A(KEYINPUT74), .B(KEYINPUT75), .Z(n350) );
  XNOR2_X1 U408 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n349) );
  XNOR2_X1 U409 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U410 ( .A(n352), .B(n351), .Z(n357) );
  XOR2_X1 U411 ( .A(G29GAT), .B(G43GAT), .Z(n354) );
  XNOR2_X1 U412 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n353) );
  XNOR2_X1 U413 ( .A(n354), .B(n353), .ZN(n396) );
  XNOR2_X1 U414 ( .A(G1GAT), .B(KEYINPUT72), .ZN(n355) );
  XNOR2_X1 U415 ( .A(n355), .B(KEYINPUT73), .ZN(n378) );
  XNOR2_X1 U416 ( .A(n396), .B(n378), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n357), .B(n356), .ZN(n362) );
  XOR2_X1 U418 ( .A(G141GAT), .B(KEYINPUT70), .Z(n359) );
  NAND2_X1 U419 ( .A1(G229GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U420 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U421 ( .A(KEYINPUT71), .B(n360), .Z(n361) );
  XOR2_X1 U422 ( .A(n362), .B(n361), .Z(n506) );
  INV_X1 U423 ( .A(n506), .ZN(n568) );
  XNOR2_X1 U424 ( .A(n363), .B(KEYINPUT46), .ZN(n381) );
  XOR2_X1 U425 ( .A(G78GAT), .B(KEYINPUT83), .Z(n365) );
  XNOR2_X1 U426 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n364) );
  XNOR2_X1 U427 ( .A(n365), .B(n364), .ZN(n370) );
  XOR2_X1 U428 ( .A(G22GAT), .B(G155GAT), .Z(n445) );
  XOR2_X1 U429 ( .A(G211GAT), .B(n445), .Z(n368) );
  XNOR2_X1 U430 ( .A(G183GAT), .B(n366), .ZN(n367) );
  XNOR2_X1 U431 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U432 ( .A(n370), .B(n369), .Z(n372) );
  NAND2_X1 U433 ( .A1(G231GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U434 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U435 ( .A(KEYINPUT82), .B(KEYINPUT12), .Z(n374) );
  XNOR2_X1 U436 ( .A(G8GAT), .B(G64GAT), .ZN(n373) );
  XNOR2_X1 U437 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U438 ( .A(n376), .B(n375), .Z(n380) );
  XNOR2_X1 U439 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U440 ( .A(n380), .B(n379), .ZN(n575) );
  NOR2_X1 U441 ( .A1(n381), .A2(n575), .ZN(n382) );
  XNOR2_X1 U442 ( .A(KEYINPUT112), .B(n382), .ZN(n399) );
  XOR2_X1 U443 ( .A(KEYINPUT11), .B(G218GAT), .Z(n385) );
  XOR2_X1 U444 ( .A(G50GAT), .B(G162GAT), .Z(n436) );
  XNOR2_X1 U445 ( .A(n383), .B(n436), .ZN(n384) );
  XNOR2_X1 U446 ( .A(n385), .B(n384), .ZN(n390) );
  XOR2_X1 U447 ( .A(KEYINPUT9), .B(KEYINPUT80), .Z(n387) );
  XNOR2_X1 U448 ( .A(KEYINPUT66), .B(G106GAT), .ZN(n386) );
  XNOR2_X1 U449 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U450 ( .A(KEYINPUT68), .B(KEYINPUT10), .Z(n392) );
  XNOR2_X1 U451 ( .A(G134GAT), .B(G92GAT), .ZN(n391) );
  XNOR2_X1 U452 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U453 ( .A(n394), .B(n393), .Z(n398) );
  XNOR2_X1 U454 ( .A(n396), .B(n395), .ZN(n397) );
  INV_X1 U455 ( .A(n559), .ZN(n463) );
  NAND2_X1 U456 ( .A1(n399), .A2(n463), .ZN(n401) );
  XNOR2_X1 U457 ( .A(n401), .B(n400), .ZN(n408) );
  XOR2_X1 U458 ( .A(KEYINPUT69), .B(KEYINPUT45), .Z(n404) );
  XNOR2_X1 U459 ( .A(KEYINPUT36), .B(KEYINPUT99), .ZN(n402) );
  NAND2_X1 U460 ( .A1(n579), .A2(n575), .ZN(n403) );
  XNOR2_X1 U461 ( .A(n404), .B(n403), .ZN(n405) );
  NOR2_X1 U462 ( .A1(n405), .A2(n568), .ZN(n406) );
  INV_X1 U463 ( .A(n572), .ZN(n462) );
  NAND2_X1 U464 ( .A1(n406), .A2(n462), .ZN(n407) );
  NAND2_X1 U465 ( .A1(n408), .A2(n407), .ZN(n409) );
  NAND2_X1 U466 ( .A1(n410), .A2(n548), .ZN(n412) );
  XNOR2_X1 U467 ( .A(n412), .B(n411), .ZN(n434) );
  XOR2_X1 U468 ( .A(G148GAT), .B(G155GAT), .Z(n414) );
  XNOR2_X1 U469 ( .A(G1GAT), .B(G57GAT), .ZN(n413) );
  XNOR2_X1 U470 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U471 ( .A(KEYINPUT4), .B(KEYINPUT89), .Z(n416) );
  XNOR2_X1 U472 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n415) );
  XNOR2_X1 U473 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U474 ( .A(n418), .B(n417), .Z(n423) );
  XOR2_X1 U475 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n420) );
  NAND2_X1 U476 ( .A1(G225GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U477 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U478 ( .A(KEYINPUT5), .B(n421), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n423), .B(n422), .ZN(n428) );
  XOR2_X1 U480 ( .A(G162GAT), .B(G85GAT), .Z(n426) );
  XNOR2_X1 U481 ( .A(n424), .B(G127GAT), .ZN(n425) );
  XNOR2_X1 U482 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U483 ( .A(n428), .B(n427), .Z(n433) );
  XOR2_X1 U484 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n430) );
  XNOR2_X1 U485 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n429) );
  XNOR2_X1 U486 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U487 ( .A(KEYINPUT2), .B(n431), .Z(n449) );
  XNOR2_X1 U488 ( .A(G29GAT), .B(n449), .ZN(n432) );
  XOR2_X1 U489 ( .A(n433), .B(n432), .Z(n550) );
  XOR2_X1 U490 ( .A(n437), .B(n436), .Z(n439) );
  NAND2_X1 U491 ( .A1(G228GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U492 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U493 ( .A(n440), .B(KEYINPUT23), .Z(n443) );
  XNOR2_X1 U494 ( .A(n441), .B(KEYINPUT22), .ZN(n442) );
  XNOR2_X1 U495 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U496 ( .A(n444), .B(KEYINPUT24), .Z(n447) );
  XNOR2_X1 U497 ( .A(n445), .B(G204GAT), .ZN(n446) );
  XNOR2_X1 U498 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U499 ( .A(n449), .B(n448), .ZN(n473) );
  NOR2_X1 U500 ( .A1(n566), .A2(n473), .ZN(n450) );
  XNOR2_X1 U501 ( .A(n450), .B(KEYINPUT55), .ZN(n451) );
  NOR2_X1 U502 ( .A1(n467), .A2(n451), .ZN(n452) );
  XNOR2_X1 U503 ( .A(n452), .B(KEYINPUT120), .ZN(n564) );
  NAND2_X1 U504 ( .A1(n555), .A2(n564), .ZN(n456) );
  XOR2_X1 U505 ( .A(G176GAT), .B(KEYINPUT121), .Z(n454) );
  XOR2_X1 U506 ( .A(KEYINPUT57), .B(KEYINPUT56), .Z(n453) );
  XNOR2_X1 U507 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U508 ( .A(n456), .B(n455), .ZN(G1349GAT) );
  NAND2_X1 U509 ( .A1(n564), .A2(n559), .ZN(n461) );
  XOR2_X1 U510 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n458) );
  XNOR2_X1 U511 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n457) );
  XNOR2_X1 U512 ( .A(n458), .B(n457), .ZN(n459) );
  XOR2_X1 U513 ( .A(KEYINPUT34), .B(KEYINPUT96), .Z(n482) );
  NAND2_X1 U514 ( .A1(n462), .A2(n568), .ZN(n495) );
  NAND2_X1 U515 ( .A1(n463), .A2(n575), .ZN(n464) );
  XOR2_X1 U516 ( .A(KEYINPUT16), .B(n464), .Z(n479) );
  INV_X1 U517 ( .A(n550), .ZN(n522) );
  AND2_X1 U518 ( .A1(n535), .A2(n524), .ZN(n465) );
  NOR2_X1 U519 ( .A1(n473), .A2(n465), .ZN(n466) );
  XOR2_X1 U520 ( .A(KEYINPUT25), .B(n466), .Z(n471) );
  XOR2_X1 U521 ( .A(KEYINPUT93), .B(KEYINPUT26), .Z(n469) );
  NAND2_X1 U522 ( .A1(n467), .A2(n473), .ZN(n468) );
  XNOR2_X1 U523 ( .A(n469), .B(n468), .ZN(n567) );
  XOR2_X1 U524 ( .A(n524), .B(KEYINPUT27), .Z(n474) );
  NOR2_X1 U525 ( .A1(n567), .A2(n474), .ZN(n547) );
  XNOR2_X1 U526 ( .A(n547), .B(KEYINPUT94), .ZN(n470) );
  NOR2_X1 U527 ( .A1(n471), .A2(n470), .ZN(n472) );
  NOR2_X1 U528 ( .A1(n522), .A2(n472), .ZN(n477) );
  XNOR2_X1 U529 ( .A(KEYINPUT28), .B(n473), .ZN(n531) );
  NOR2_X1 U530 ( .A1(n474), .A2(n531), .ZN(n475) );
  NAND2_X1 U531 ( .A1(n522), .A2(n475), .ZN(n537) );
  NOR2_X1 U532 ( .A1(n537), .A2(n535), .ZN(n476) );
  NOR2_X1 U533 ( .A1(n477), .A2(n476), .ZN(n491) );
  INV_X1 U534 ( .A(n491), .ZN(n478) );
  NAND2_X1 U535 ( .A1(n479), .A2(n478), .ZN(n507) );
  NOR2_X1 U536 ( .A1(n495), .A2(n507), .ZN(n480) );
  XOR2_X1 U537 ( .A(KEYINPUT95), .B(n480), .Z(n489) );
  NAND2_X1 U538 ( .A1(n489), .A2(n522), .ZN(n481) );
  XNOR2_X1 U539 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U540 ( .A(G1GAT), .B(n483), .Z(G1324GAT) );
  NAND2_X1 U541 ( .A1(n489), .A2(n524), .ZN(n484) );
  XNOR2_X1 U542 ( .A(n484), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U543 ( .A(KEYINPUT35), .B(KEYINPUT98), .Z(n486) );
  NAND2_X1 U544 ( .A1(n489), .A2(n535), .ZN(n485) );
  XNOR2_X1 U545 ( .A(n486), .B(n485), .ZN(n488) );
  XOR2_X1 U546 ( .A(G15GAT), .B(KEYINPUT97), .Z(n487) );
  XNOR2_X1 U547 ( .A(n488), .B(n487), .ZN(G1326GAT) );
  NAND2_X1 U548 ( .A1(n489), .A2(n531), .ZN(n490) );
  XNOR2_X1 U549 ( .A(n490), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U550 ( .A(G29GAT), .B(KEYINPUT39), .Z(n498) );
  XOR2_X1 U551 ( .A(KEYINPUT37), .B(KEYINPUT100), .Z(n494) );
  NOR2_X1 U552 ( .A1(n575), .A2(n491), .ZN(n492) );
  NAND2_X1 U553 ( .A1(n579), .A2(n492), .ZN(n493) );
  XNOR2_X1 U554 ( .A(n494), .B(n493), .ZN(n521) );
  NOR2_X1 U555 ( .A1(n495), .A2(n521), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n496), .B(KEYINPUT38), .ZN(n503) );
  NAND2_X1 U557 ( .A1(n522), .A2(n503), .ZN(n497) );
  XNOR2_X1 U558 ( .A(n498), .B(n497), .ZN(G1328GAT) );
  XOR2_X1 U559 ( .A(G36GAT), .B(KEYINPUT101), .Z(n500) );
  NAND2_X1 U560 ( .A1(n524), .A2(n503), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(G1329GAT) );
  NAND2_X1 U562 ( .A1(n503), .A2(n535), .ZN(n501) );
  XNOR2_X1 U563 ( .A(n501), .B(KEYINPUT40), .ZN(n502) );
  XNOR2_X1 U564 ( .A(G43GAT), .B(n502), .ZN(G1330GAT) );
  NAND2_X1 U565 ( .A1(n503), .A2(n531), .ZN(n504) );
  XNOR2_X1 U566 ( .A(n504), .B(KEYINPUT102), .ZN(n505) );
  XNOR2_X1 U567 ( .A(G50GAT), .B(n505), .ZN(G1331GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT42), .B(KEYINPUT103), .Z(n509) );
  NAND2_X1 U569 ( .A1(n506), .A2(n555), .ZN(n520) );
  NOR2_X1 U570 ( .A1(n507), .A2(n520), .ZN(n516) );
  NAND2_X1 U571 ( .A1(n516), .A2(n522), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U573 ( .A(G57GAT), .B(n510), .ZN(G1332GAT) );
  NAND2_X1 U574 ( .A1(n516), .A2(n524), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n511), .B(KEYINPUT104), .ZN(n512) );
  XNOR2_X1 U576 ( .A(G64GAT), .B(n512), .ZN(G1333GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n514) );
  NAND2_X1 U578 ( .A1(n516), .A2(n535), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U580 ( .A(G71GAT), .B(n515), .ZN(G1334GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n518) );
  NAND2_X1 U582 ( .A1(n516), .A2(n531), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U584 ( .A(G78GAT), .B(n519), .Z(G1335GAT) );
  NOR2_X1 U585 ( .A1(n521), .A2(n520), .ZN(n532) );
  NAND2_X1 U586 ( .A1(n522), .A2(n532), .ZN(n523) );
  XNOR2_X1 U587 ( .A(G85GAT), .B(n523), .ZN(G1336GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n526) );
  NAND2_X1 U589 ( .A1(n532), .A2(n524), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U591 ( .A(G92GAT), .B(n527), .ZN(G1337GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n529) );
  NAND2_X1 U593 ( .A1(n532), .A2(n535), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U595 ( .A(G99GAT), .B(n530), .ZN(G1338GAT) );
  NAND2_X1 U596 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U597 ( .A(n533), .B(KEYINPUT44), .ZN(n534) );
  XNOR2_X1 U598 ( .A(G106GAT), .B(n534), .ZN(G1339GAT) );
  NAND2_X1 U599 ( .A1(n548), .A2(n535), .ZN(n536) );
  NOR2_X1 U600 ( .A1(n537), .A2(n536), .ZN(n543) );
  NAND2_X1 U601 ( .A1(n568), .A2(n543), .ZN(n538) );
  XNOR2_X1 U602 ( .A(n538), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U603 ( .A(G120GAT), .B(KEYINPUT49), .Z(n540) );
  NAND2_X1 U604 ( .A1(n543), .A2(n555), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(G1341GAT) );
  NAND2_X1 U606 ( .A1(n543), .A2(n575), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n541), .B(KEYINPUT50), .ZN(n542) );
  XNOR2_X1 U608 ( .A(G127GAT), .B(n542), .ZN(G1342GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n545) );
  NAND2_X1 U610 ( .A1(n543), .A2(n559), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U612 ( .A(G134GAT), .B(n546), .ZN(G1343GAT) );
  NAND2_X1 U613 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U614 ( .A1(n550), .A2(n549), .ZN(n560) );
  NAND2_X1 U615 ( .A1(n560), .A2(n568), .ZN(n551) );
  XNOR2_X1 U616 ( .A(G141GAT), .B(n551), .ZN(G1344GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT116), .B(KEYINPUT53), .Z(n553) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U620 ( .A(KEYINPUT115), .B(n554), .Z(n557) );
  NAND2_X1 U621 ( .A1(n560), .A2(n555), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(G1345GAT) );
  NAND2_X1 U623 ( .A1(n560), .A2(n575), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U625 ( .A(G162GAT), .B(KEYINPUT117), .Z(n562) );
  NAND2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(G1347GAT) );
  NAND2_X1 U628 ( .A1(n564), .A2(n568), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G169GAT), .B(n563), .ZN(G1348GAT) );
  NAND2_X1 U630 ( .A1(n564), .A2(n575), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(G183GAT), .ZN(G1350GAT) );
  NOR2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n580) );
  NAND2_X1 U633 ( .A1(n568), .A2(n580), .ZN(n571) );
  XOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT60), .Z(n569) );
  XNOR2_X1 U635 ( .A(KEYINPUT59), .B(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .Z(n574) );
  NAND2_X1 U638 ( .A1(n580), .A2(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n577) );
  NAND2_X1 U641 ( .A1(n580), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G211GAT), .B(n578), .ZN(G1354GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n582) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

