

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592;

  XOR2_X1 U324 ( .A(KEYINPUT54), .B(n418), .Z(n292) );
  XNOR2_X1 U325 ( .A(n403), .B(n402), .ZN(n540) );
  XNOR2_X1 U326 ( .A(KEYINPUT48), .B(KEYINPUT116), .ZN(n402) );
  NOR2_X1 U327 ( .A1(n454), .A2(n543), .ZN(n578) );
  XOR2_X1 U328 ( .A(n453), .B(n452), .Z(n533) );
  XOR2_X2 U329 ( .A(n373), .B(n372), .Z(n582) );
  XOR2_X1 U330 ( .A(G50GAT), .B(G162GAT), .Z(n420) );
  INV_X1 U331 ( .A(KEYINPUT9), .ZN(n340) );
  XNOR2_X1 U332 ( .A(n341), .B(n340), .ZN(n352) );
  XNOR2_X1 U333 ( .A(n355), .B(KEYINPUT105), .ZN(n356) );
  XNOR2_X1 U334 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U335 ( .A(n568), .B(n356), .ZN(n589) );
  INV_X1 U336 ( .A(G190GAT), .ZN(n455) );
  XOR2_X1 U337 ( .A(n475), .B(KEYINPUT28), .Z(n535) );
  XNOR2_X1 U338 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U339 ( .A(n458), .B(n457), .ZN(G1351GAT) );
  XOR2_X1 U340 ( .A(KEYINPUT55), .B(KEYINPUT122), .Z(n435) );
  XOR2_X1 U341 ( .A(KEYINPUT90), .B(G57GAT), .Z(n294) );
  XNOR2_X1 U342 ( .A(G127GAT), .B(G148GAT), .ZN(n293) );
  XNOR2_X1 U343 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U344 ( .A(G85GAT), .B(G162GAT), .Z(n296) );
  XNOR2_X1 U345 ( .A(G29GAT), .B(G155GAT), .ZN(n295) );
  XNOR2_X1 U346 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U347 ( .A(n298), .B(n297), .ZN(n316) );
  XOR2_X1 U348 ( .A(KEYINPUT5), .B(KEYINPUT88), .Z(n300) );
  XNOR2_X1 U349 ( .A(KEYINPUT91), .B(KEYINPUT89), .ZN(n299) );
  XNOR2_X1 U350 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U351 ( .A(KEYINPUT92), .B(KEYINPUT6), .Z(n302) );
  XNOR2_X1 U352 ( .A(G1GAT), .B(KEYINPUT4), .ZN(n301) );
  XNOR2_X1 U353 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U354 ( .A(n304), .B(n303), .Z(n314) );
  XOR2_X1 U355 ( .A(KEYINPUT86), .B(KEYINPUT2), .Z(n306) );
  XNOR2_X1 U356 ( .A(KEYINPUT3), .B(KEYINPUT87), .ZN(n305) );
  XNOR2_X1 U357 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U358 ( .A(G141GAT), .B(n307), .Z(n424) );
  XOR2_X1 U359 ( .A(G120GAT), .B(KEYINPUT0), .Z(n309) );
  XNOR2_X1 U360 ( .A(G113GAT), .B(G134GAT), .ZN(n308) );
  XNOR2_X1 U361 ( .A(n309), .B(n308), .ZN(n449) );
  XOR2_X1 U362 ( .A(n449), .B(KEYINPUT1), .Z(n311) );
  NAND2_X1 U363 ( .A1(G225GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U364 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U365 ( .A(n424), .B(n312), .ZN(n313) );
  XNOR2_X1 U366 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U367 ( .A(n316), .B(n315), .ZN(n527) );
  XNOR2_X1 U368 ( .A(G1GAT), .B(G64GAT), .ZN(n317) );
  XOR2_X1 U369 ( .A(G15GAT), .B(G127GAT), .Z(n439) );
  XOR2_X1 U370 ( .A(n317), .B(n439), .Z(n330) );
  XNOR2_X1 U371 ( .A(G22GAT), .B(G155GAT), .ZN(n318) );
  XNOR2_X1 U372 ( .A(n318), .B(G78GAT), .ZN(n429) );
  XOR2_X1 U373 ( .A(KEYINPUT77), .B(n429), .Z(n320) );
  NAND2_X1 U374 ( .A1(G231GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U375 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U376 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n322) );
  XNOR2_X1 U377 ( .A(KEYINPUT12), .B(KEYINPUT78), .ZN(n321) );
  XNOR2_X1 U378 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U379 ( .A(n324), .B(n323), .Z(n328) );
  XOR2_X1 U380 ( .A(G71GAT), .B(G57GAT), .Z(n325) );
  XOR2_X1 U381 ( .A(KEYINPUT13), .B(n325), .Z(n373) );
  XNOR2_X1 U382 ( .A(G8GAT), .B(G183GAT), .ZN(n326) );
  XOR2_X1 U383 ( .A(n326), .B(G211GAT), .Z(n416) );
  XOR2_X1 U384 ( .A(n373), .B(n416), .Z(n327) );
  XNOR2_X1 U385 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U386 ( .A(n330), .B(n329), .Z(n587) );
  INV_X1 U387 ( .A(n587), .ZN(n565) );
  XOR2_X1 U388 ( .A(KEYINPUT11), .B(KEYINPUT65), .Z(n332) );
  XNOR2_X1 U389 ( .A(G92GAT), .B(KEYINPUT64), .ZN(n331) );
  XNOR2_X1 U390 ( .A(n332), .B(n331), .ZN(n337) );
  XOR2_X1 U391 ( .A(G36GAT), .B(G190GAT), .Z(n404) );
  XNOR2_X1 U392 ( .A(G99GAT), .B(G85GAT), .ZN(n333) );
  XNOR2_X1 U393 ( .A(n333), .B(KEYINPUT72), .ZN(n358) );
  XOR2_X1 U394 ( .A(n404), .B(n358), .Z(n335) );
  NAND2_X1 U395 ( .A1(G232GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U396 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U397 ( .A(n337), .B(n336), .ZN(n354) );
  XOR2_X1 U398 ( .A(G29GAT), .B(G43GAT), .Z(n339) );
  XNOR2_X1 U399 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n338) );
  XNOR2_X1 U400 ( .A(n339), .B(n338), .ZN(n387) );
  XNOR2_X1 U401 ( .A(n387), .B(G134GAT), .ZN(n341) );
  INV_X1 U402 ( .A(KEYINPUT74), .ZN(n342) );
  NAND2_X1 U403 ( .A1(KEYINPUT76), .A2(n342), .ZN(n345) );
  INV_X1 U404 ( .A(KEYINPUT76), .ZN(n343) );
  NAND2_X1 U405 ( .A1(n343), .A2(KEYINPUT74), .ZN(n344) );
  NAND2_X1 U406 ( .A1(n345), .A2(n344), .ZN(n347) );
  XNOR2_X1 U407 ( .A(G218GAT), .B(KEYINPUT75), .ZN(n346) );
  XNOR2_X1 U408 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U409 ( .A(n348), .B(KEYINPUT10), .ZN(n350) );
  XOR2_X1 U410 ( .A(G106GAT), .B(n420), .Z(n349) );
  XNOR2_X1 U411 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U412 ( .A(n354), .B(n353), .Z(n568) );
  INV_X1 U413 ( .A(KEYINPUT36), .ZN(n355) );
  NOR2_X1 U414 ( .A1(n565), .A2(n589), .ZN(n357) );
  XNOR2_X1 U415 ( .A(KEYINPUT45), .B(n357), .ZN(n393) );
  INV_X1 U416 ( .A(KEYINPUT33), .ZN(n359) );
  XNOR2_X1 U417 ( .A(n359), .B(n358), .ZN(n361) );
  NAND2_X1 U418 ( .A1(G230GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U419 ( .A(n361), .B(n360), .ZN(n365) );
  XOR2_X1 U420 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n363) );
  XNOR2_X1 U421 ( .A(G120GAT), .B(G78GAT), .ZN(n362) );
  XNOR2_X1 U422 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U423 ( .A(n365), .B(n364), .ZN(n371) );
  XOR2_X1 U424 ( .A(G148GAT), .B(KEYINPUT70), .Z(n367) );
  XNOR2_X1 U425 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n366) );
  XNOR2_X1 U426 ( .A(n367), .B(n366), .ZN(n428) );
  XOR2_X1 U427 ( .A(G64GAT), .B(G92GAT), .Z(n369) );
  XNOR2_X1 U428 ( .A(G176GAT), .B(G204GAT), .ZN(n368) );
  XNOR2_X1 U429 ( .A(n369), .B(n368), .ZN(n407) );
  XOR2_X1 U430 ( .A(n428), .B(n407), .Z(n370) );
  XNOR2_X1 U431 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U432 ( .A(KEYINPUT30), .B(G1GAT), .Z(n375) );
  XNOR2_X1 U433 ( .A(G169GAT), .B(G15GAT), .ZN(n374) );
  XNOR2_X1 U434 ( .A(n375), .B(n374), .ZN(n391) );
  XOR2_X1 U435 ( .A(G8GAT), .B(KEYINPUT69), .Z(n377) );
  XNOR2_X1 U436 ( .A(KEYINPUT29), .B(KEYINPUT68), .ZN(n376) );
  XNOR2_X1 U437 ( .A(n377), .B(n376), .ZN(n385) );
  NAND2_X1 U438 ( .A1(G229GAT), .A2(G233GAT), .ZN(n383) );
  XOR2_X1 U439 ( .A(G113GAT), .B(G197GAT), .Z(n379) );
  XNOR2_X1 U440 ( .A(G22GAT), .B(G141GAT), .ZN(n378) );
  XNOR2_X1 U441 ( .A(n379), .B(n378), .ZN(n381) );
  XOR2_X1 U442 ( .A(G36GAT), .B(G50GAT), .Z(n380) );
  XNOR2_X1 U443 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U444 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U445 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U446 ( .A(n386), .B(KEYINPUT67), .Z(n389) );
  XNOR2_X1 U447 ( .A(n387), .B(KEYINPUT66), .ZN(n388) );
  XNOR2_X1 U448 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U449 ( .A(n391), .B(n390), .ZN(n558) );
  INV_X1 U450 ( .A(n558), .ZN(n571) );
  AND2_X1 U451 ( .A1(n582), .A2(n558), .ZN(n392) );
  AND2_X1 U452 ( .A1(n393), .A2(n392), .ZN(n394) );
  XOR2_X1 U453 ( .A(n394), .B(KEYINPUT115), .Z(n401) );
  INV_X1 U454 ( .A(n568), .ZN(n553) );
  XNOR2_X1 U455 ( .A(KEYINPUT41), .B(n582), .ZN(n574) );
  NAND2_X1 U456 ( .A1(n571), .A2(n574), .ZN(n396) );
  XNOR2_X1 U457 ( .A(KEYINPUT114), .B(KEYINPUT46), .ZN(n395) );
  XNOR2_X1 U458 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U459 ( .A(KEYINPUT113), .B(n565), .Z(n580) );
  NAND2_X1 U460 ( .A1(n397), .A2(n580), .ZN(n398) );
  NOR2_X1 U461 ( .A1(n553), .A2(n398), .ZN(n399) );
  XOR2_X1 U462 ( .A(KEYINPUT47), .B(n399), .Z(n400) );
  NOR2_X1 U463 ( .A1(n401), .A2(n400), .ZN(n403) );
  XOR2_X1 U464 ( .A(KEYINPUT93), .B(n404), .Z(n406) );
  NAND2_X1 U465 ( .A1(G226GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U466 ( .A(n406), .B(n405), .ZN(n408) );
  XOR2_X1 U467 ( .A(n408), .B(n407), .Z(n414) );
  XOR2_X1 U468 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n410) );
  XNOR2_X1 U469 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n409) );
  XNOR2_X1 U470 ( .A(n410), .B(n409), .ZN(n448) );
  XOR2_X1 U471 ( .A(KEYINPUT85), .B(KEYINPUT21), .Z(n412) );
  XNOR2_X1 U472 ( .A(G197GAT), .B(G218GAT), .ZN(n411) );
  XNOR2_X1 U473 ( .A(n412), .B(n411), .ZN(n419) );
  XNOR2_X1 U474 ( .A(n448), .B(n419), .ZN(n413) );
  XNOR2_X1 U475 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U476 ( .A(n416), .B(n415), .Z(n473) );
  BUF_X1 U477 ( .A(n473), .Z(n531) );
  XNOR2_X1 U478 ( .A(KEYINPUT121), .B(n531), .ZN(n417) );
  NOR2_X1 U479 ( .A1(n540), .A2(n417), .ZN(n418) );
  NOR2_X1 U480 ( .A1(n527), .A2(n292), .ZN(n461) );
  XOR2_X1 U481 ( .A(n419), .B(G204GAT), .Z(n422) );
  XNOR2_X1 U482 ( .A(n420), .B(G211GAT), .ZN(n421) );
  XNOR2_X1 U483 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U484 ( .A(n424), .B(n423), .ZN(n433) );
  XOR2_X1 U485 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n426) );
  NAND2_X1 U486 ( .A1(G228GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U487 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U488 ( .A(n427), .B(KEYINPUT22), .Z(n431) );
  XNOR2_X1 U489 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U490 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U491 ( .A(n433), .B(n432), .ZN(n475) );
  NAND2_X1 U492 ( .A1(n461), .A2(n475), .ZN(n434) );
  XNOR2_X1 U493 ( .A(n435), .B(n434), .ZN(n454) );
  XOR2_X1 U494 ( .A(KEYINPUT83), .B(G99GAT), .Z(n437) );
  XNOR2_X1 U495 ( .A(G43GAT), .B(G190GAT), .ZN(n436) );
  XNOR2_X1 U496 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U497 ( .A(n439), .B(n438), .Z(n441) );
  NAND2_X1 U498 ( .A1(G227GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U499 ( .A(n441), .B(n440), .ZN(n453) );
  XOR2_X1 U500 ( .A(G176GAT), .B(KEYINPUT84), .Z(n443) );
  XNOR2_X1 U501 ( .A(KEYINPUT20), .B(G183GAT), .ZN(n442) );
  XNOR2_X1 U502 ( .A(n443), .B(n442), .ZN(n447) );
  XOR2_X1 U503 ( .A(KEYINPUT82), .B(KEYINPUT80), .Z(n445) );
  XNOR2_X1 U504 ( .A(KEYINPUT81), .B(G71GAT), .ZN(n444) );
  XNOR2_X1 U505 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U506 ( .A(n447), .B(n446), .Z(n451) );
  XNOR2_X1 U507 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U508 ( .A(n451), .B(n450), .ZN(n452) );
  INV_X1 U509 ( .A(n533), .ZN(n543) );
  NAND2_X1 U510 ( .A1(n578), .A2(n553), .ZN(n458) );
  XOR2_X1 U511 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n456) );
  XNOR2_X1 U512 ( .A(KEYINPUT26), .B(KEYINPUT94), .ZN(n460) );
  NOR2_X1 U513 ( .A1(n533), .A2(n475), .ZN(n459) );
  XNOR2_X1 U514 ( .A(n460), .B(n459), .ZN(n557) );
  NAND2_X1 U515 ( .A1(n461), .A2(n557), .ZN(n462) );
  XOR2_X1 U516 ( .A(KEYINPUT125), .B(n462), .Z(n590) );
  INV_X1 U517 ( .A(n590), .ZN(n586) );
  NAND2_X1 U518 ( .A1(n586), .A2(n571), .ZN(n464) );
  XOR2_X1 U519 ( .A(KEYINPUT127), .B(KEYINPUT60), .Z(n463) );
  XNOR2_X1 U520 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U521 ( .A(n465), .B(KEYINPUT59), .ZN(n467) );
  XOR2_X1 U522 ( .A(G197GAT), .B(KEYINPUT126), .Z(n466) );
  XNOR2_X1 U523 ( .A(n467), .B(n466), .ZN(G1352GAT) );
  XOR2_X1 U524 ( .A(KEYINPUT34), .B(KEYINPUT102), .Z(n491) );
  XNOR2_X1 U525 ( .A(KEYINPUT16), .B(KEYINPUT79), .ZN(n469) );
  NOR2_X1 U526 ( .A1(n553), .A2(n565), .ZN(n468) );
  XNOR2_X1 U527 ( .A(n469), .B(n468), .ZN(n486) );
  XNOR2_X1 U528 ( .A(n531), .B(KEYINPUT27), .ZN(n471) );
  NAND2_X1 U529 ( .A1(n527), .A2(n471), .ZN(n539) );
  INV_X1 U530 ( .A(n535), .ZN(n542) );
  NAND2_X1 U531 ( .A1(n543), .A2(n542), .ZN(n470) );
  NOR2_X1 U532 ( .A1(n539), .A2(n470), .ZN(n484) );
  NAND2_X1 U533 ( .A1(n557), .A2(n471), .ZN(n472) );
  XNOR2_X1 U534 ( .A(KEYINPUT95), .B(n472), .ZN(n481) );
  XOR2_X1 U535 ( .A(KEYINPUT98), .B(KEYINPUT25), .Z(n478) );
  AND2_X1 U536 ( .A1(n473), .A2(n533), .ZN(n474) );
  XOR2_X1 U537 ( .A(KEYINPUT96), .B(n474), .Z(n476) );
  NAND2_X1 U538 ( .A1(n476), .A2(n475), .ZN(n477) );
  XNOR2_X1 U539 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U540 ( .A(n479), .B(KEYINPUT97), .ZN(n480) );
  NOR2_X1 U541 ( .A1(n481), .A2(n480), .ZN(n482) );
  NOR2_X1 U542 ( .A1(n527), .A2(n482), .ZN(n483) );
  NOR2_X1 U543 ( .A1(n484), .A2(n483), .ZN(n485) );
  XOR2_X1 U544 ( .A(KEYINPUT99), .B(n485), .Z(n499) );
  NOR2_X1 U545 ( .A1(n486), .A2(n499), .ZN(n487) );
  XNOR2_X1 U546 ( .A(n487), .B(KEYINPUT100), .ZN(n517) );
  NAND2_X1 U547 ( .A1(n582), .A2(n571), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n488), .B(KEYINPUT73), .ZN(n504) );
  NAND2_X1 U549 ( .A1(n517), .A2(n504), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n489), .B(KEYINPUT101), .ZN(n497) );
  NAND2_X1 U551 ( .A1(n497), .A2(n527), .ZN(n490) );
  XNOR2_X1 U552 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U553 ( .A(G1GAT), .B(n492), .Z(G1324GAT) );
  XOR2_X1 U554 ( .A(G8GAT), .B(KEYINPUT103), .Z(n494) );
  NAND2_X1 U555 ( .A1(n497), .A2(n531), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n494), .B(n493), .ZN(G1325GAT) );
  XOR2_X1 U557 ( .A(G15GAT), .B(KEYINPUT35), .Z(n496) );
  NAND2_X1 U558 ( .A1(n497), .A2(n533), .ZN(n495) );
  XNOR2_X1 U559 ( .A(n496), .B(n495), .ZN(G1326GAT) );
  NAND2_X1 U560 ( .A1(n535), .A2(n497), .ZN(n498) );
  XNOR2_X1 U561 ( .A(G22GAT), .B(n498), .ZN(G1327GAT) );
  NOR2_X1 U562 ( .A1(n589), .A2(n499), .ZN(n500) );
  NAND2_X1 U563 ( .A1(n565), .A2(n500), .ZN(n501) );
  XNOR2_X1 U564 ( .A(KEYINPUT106), .B(n501), .ZN(n503) );
  XOR2_X1 U565 ( .A(KEYINPUT107), .B(KEYINPUT37), .Z(n502) );
  XNOR2_X1 U566 ( .A(n503), .B(n502), .ZN(n526) );
  NAND2_X1 U567 ( .A1(n504), .A2(n526), .ZN(n505) );
  XOR2_X1 U568 ( .A(KEYINPUT38), .B(n505), .Z(n514) );
  NAND2_X1 U569 ( .A1(n514), .A2(n527), .ZN(n509) );
  XOR2_X1 U570 ( .A(KEYINPUT104), .B(KEYINPUT39), .Z(n507) );
  XNOR2_X1 U571 ( .A(G29GAT), .B(KEYINPUT108), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n509), .B(n508), .ZN(G1328GAT) );
  XOR2_X1 U574 ( .A(G36GAT), .B(KEYINPUT109), .Z(n511) );
  NAND2_X1 U575 ( .A1(n514), .A2(n531), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(G1329GAT) );
  NAND2_X1 U577 ( .A1(n514), .A2(n533), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n512), .B(KEYINPUT40), .ZN(n513) );
  XNOR2_X1 U579 ( .A(G43GAT), .B(n513), .ZN(G1330GAT) );
  NAND2_X1 U580 ( .A1(n514), .A2(n535), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n515), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U582 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n519) );
  NAND2_X1 U583 ( .A1(n574), .A2(n558), .ZN(n516) );
  XOR2_X1 U584 ( .A(KEYINPUT110), .B(n516), .Z(n525) );
  AND2_X1 U585 ( .A1(n517), .A2(n525), .ZN(n522) );
  NAND2_X1 U586 ( .A1(n527), .A2(n522), .ZN(n518) );
  XNOR2_X1 U587 ( .A(n519), .B(n518), .ZN(G1332GAT) );
  NAND2_X1 U588 ( .A1(n531), .A2(n522), .ZN(n520) );
  XNOR2_X1 U589 ( .A(n520), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U590 ( .A1(n522), .A2(n533), .ZN(n521) );
  XNOR2_X1 U591 ( .A(n521), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U592 ( .A(G78GAT), .B(KEYINPUT43), .Z(n524) );
  NAND2_X1 U593 ( .A1(n522), .A2(n535), .ZN(n523) );
  XNOR2_X1 U594 ( .A(n524), .B(n523), .ZN(G1335GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n529) );
  AND2_X1 U596 ( .A1(n526), .A2(n525), .ZN(n536) );
  NAND2_X1 U597 ( .A1(n536), .A2(n527), .ZN(n528) );
  XNOR2_X1 U598 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U599 ( .A(G85GAT), .B(n530), .ZN(G1336GAT) );
  NAND2_X1 U600 ( .A1(n531), .A2(n536), .ZN(n532) );
  XNOR2_X1 U601 ( .A(n532), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U602 ( .A1(n536), .A2(n533), .ZN(n534) );
  XNOR2_X1 U603 ( .A(n534), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U604 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U605 ( .A(n537), .B(KEYINPUT44), .ZN(n538) );
  XNOR2_X1 U606 ( .A(G106GAT), .B(n538), .ZN(G1339GAT) );
  NOR2_X1 U607 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U608 ( .A(KEYINPUT117), .B(n541), .Z(n556) );
  NAND2_X1 U609 ( .A1(n556), .A2(n542), .ZN(n544) );
  NOR2_X1 U610 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U611 ( .A(n545), .B(KEYINPUT118), .Z(n549) );
  INV_X1 U612 ( .A(n549), .ZN(n552) );
  NAND2_X1 U613 ( .A1(n552), .A2(n571), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n546), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U615 ( .A(G120GAT), .B(KEYINPUT49), .Z(n548) );
  NAND2_X1 U616 ( .A1(n552), .A2(n574), .ZN(n547) );
  XNOR2_X1 U617 ( .A(n548), .B(n547), .ZN(G1341GAT) );
  NOR2_X1 U618 ( .A1(n580), .A2(n549), .ZN(n550) );
  XOR2_X1 U619 ( .A(KEYINPUT50), .B(n550), .Z(n551) );
  XNOR2_X1 U620 ( .A(G127GAT), .B(n551), .ZN(G1342GAT) );
  XOR2_X1 U621 ( .A(G134GAT), .B(KEYINPUT51), .Z(n555) );
  NAND2_X1 U622 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(G1343GAT) );
  NAND2_X1 U624 ( .A1(n557), .A2(n556), .ZN(n567) );
  NOR2_X1 U625 ( .A1(n558), .A2(n567), .ZN(n559) );
  XOR2_X1 U626 ( .A(G141GAT), .B(n559), .Z(G1344GAT) );
  INV_X1 U627 ( .A(n574), .ZN(n560) );
  NOR2_X1 U628 ( .A1(n567), .A2(n560), .ZN(n564) );
  XOR2_X1 U629 ( .A(KEYINPUT53), .B(KEYINPUT119), .Z(n562) );
  XNOR2_X1 U630 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n561) );
  XNOR2_X1 U631 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U632 ( .A(n564), .B(n563), .ZN(G1345GAT) );
  NOR2_X1 U633 ( .A1(n565), .A2(n567), .ZN(n566) );
  XOR2_X1 U634 ( .A(G155GAT), .B(n566), .Z(G1346GAT) );
  NOR2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U636 ( .A(G162GAT), .B(n569), .Z(n570) );
  XNOR2_X1 U637 ( .A(KEYINPUT120), .B(n570), .ZN(G1347GAT) );
  XOR2_X1 U638 ( .A(G169GAT), .B(KEYINPUT123), .Z(n573) );
  NAND2_X1 U639 ( .A1(n578), .A2(n571), .ZN(n572) );
  XNOR2_X1 U640 ( .A(n573), .B(n572), .ZN(G1348GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n576) );
  NAND2_X1 U642 ( .A1(n578), .A2(n574), .ZN(n575) );
  XNOR2_X1 U643 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U644 ( .A(G176GAT), .B(n577), .ZN(G1349GAT) );
  INV_X1 U645 ( .A(n578), .ZN(n579) );
  NOR2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U647 ( .A(G183GAT), .B(n581), .Z(G1350GAT) );
  XOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT61), .Z(n585) );
  INV_X1 U649 ( .A(n582), .ZN(n583) );
  NAND2_X1 U650 ( .A1(n586), .A2(n583), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n585), .B(n584), .ZN(G1353GAT) );
  NAND2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n588), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U655 ( .A(KEYINPUT62), .B(n591), .Z(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

