//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 0 0 0 0 1 0 0 1 1 1 0 0 1 1 1 1 0 0 0 0 1 1 1 0 1 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 0 1 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n806, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1026,
    new_n1027;
  XNOR2_X1  g000(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT96), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G155gat), .ZN(new_n204));
  XOR2_X1   g003(.A(G183gat), .B(G211gat), .Z(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT95), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT93), .ZN(new_n209));
  INV_X1    g008(.A(G57gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n209), .B1(new_n210), .B2(G64gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(G64gat), .ZN(new_n212));
  INV_X1    g011(.A(G64gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n213), .A2(KEYINPUT93), .A3(G57gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n211), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT94), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT94), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n211), .A2(new_n214), .A3(new_n217), .A4(new_n212), .ZN(new_n218));
  NAND2_X1  g017(.A1(G71gat), .A2(G78gat), .ZN(new_n219));
  OR2_X1    g018(.A1(G71gat), .A2(G78gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT9), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AND3_X1   g021(.A1(new_n216), .A2(new_n218), .A3(new_n222), .ZN(new_n223));
  XOR2_X1   g022(.A(G71gat), .B(G78gat), .Z(new_n224));
  XNOR2_X1  g023(.A(G57gat), .B(G64gat), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n224), .B(KEYINPUT92), .C1(new_n221), .C2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT92), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n213), .A2(G57gat), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n221), .B1(new_n228), .B2(new_n212), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n220), .A2(new_n219), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n227), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n226), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n208), .B1(new_n223), .B2(new_n232), .ZN(new_n233));
  AND2_X1   g032(.A1(new_n226), .A2(new_n231), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n216), .A2(new_n218), .A3(new_n222), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n234), .A2(KEYINPUT95), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  OR2_X1    g036(.A1(new_n237), .A2(KEYINPUT21), .ZN(new_n238));
  NAND2_X1  g037(.A1(G231gat), .A2(G233gat), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n238), .B(new_n239), .Z(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G127gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n238), .B(new_n239), .ZN(new_n242));
  INV_X1    g041(.A(G127gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n237), .A2(KEYINPUT21), .ZN(new_n245));
  XNOR2_X1  g044(.A(G15gat), .B(G22gat), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT16), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT88), .B1(new_n247), .B2(G1gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NOR3_X1   g048(.A1(new_n247), .A2(KEYINPUT88), .A3(G1gat), .ZN(new_n250));
  OAI22_X1  g049(.A1(new_n249), .A2(new_n250), .B1(G1gat), .B2(new_n246), .ZN(new_n251));
  OAI21_X1  g050(.A(KEYINPUT89), .B1(new_n246), .B2(G1gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(G8gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n251), .B(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n245), .A2(new_n254), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n241), .A2(new_n244), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n255), .B1(new_n241), .B2(new_n244), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n207), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n244), .ZN(new_n259));
  INV_X1    g058(.A(new_n255), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n241), .A2(new_n244), .A3(new_n255), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n261), .A2(new_n262), .A3(new_n206), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n258), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G190gat), .B(G218gat), .ZN(new_n265));
  OR2_X1    g064(.A1(new_n265), .A2(KEYINPUT99), .ZN(new_n266));
  NAND2_X1  g065(.A1(G85gat), .A2(G92gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n267), .B(KEYINPUT7), .ZN(new_n268));
  OR2_X1    g067(.A1(KEYINPUT98), .A2(G85gat), .ZN(new_n269));
  INV_X1    g068(.A(G92gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(KEYINPUT98), .A2(G85gat), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(G99gat), .A2(G106gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT8), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n268), .A2(new_n272), .A3(new_n274), .ZN(new_n275));
  XOR2_X1   g074(.A(G99gat), .B(G106gat), .Z(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n276), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n278), .A2(new_n268), .A3(new_n272), .A4(new_n274), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT17), .ZN(new_n282));
  XNOR2_X1  g081(.A(KEYINPUT86), .B(G50gat), .ZN(new_n283));
  INV_X1    g082(.A(G43gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OR2_X1    g084(.A1(new_n285), .A2(KEYINPUT87), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n284), .A2(G50gat), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n287), .B1(new_n285), .B2(KEYINPUT87), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT15), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  NOR2_X1   g088(.A1(G29gat), .A2(G36gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n290), .B(KEYINPUT14), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n291), .B1(G29gat), .B2(G36gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT15), .ZN(new_n293));
  XNOR2_X1  g092(.A(G43gat), .B(G50gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT84), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n296), .B1(new_n295), .B2(new_n294), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n289), .A2(new_n298), .ZN(new_n299));
  AND2_X1   g098(.A1(new_n291), .A2(KEYINPUT85), .ZN(new_n300));
  NAND2_X1  g099(.A1(G29gat), .A2(G36gat), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n301), .B1(new_n291), .B2(KEYINPUT85), .ZN(new_n302));
  OAI221_X1 g101(.A(new_n296), .B1(new_n295), .B2(new_n294), .C1(new_n300), .C2(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n282), .B1(new_n299), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n303), .B(new_n282), .C1(new_n289), .C2(new_n298), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n281), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n299), .A2(new_n303), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(new_n281), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT41), .ZN(new_n310));
  NAND2_X1  g109(.A1(G232gat), .A2(G233gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n266), .B1(new_n307), .B2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(G134gat), .B(G162gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n311), .A2(new_n310), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n316), .B(KEYINPUT97), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n265), .A2(KEYINPUT99), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n317), .B(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n314), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n266), .B(new_n320), .C1(new_n307), .C2(new_n312), .ZN(new_n321));
  AND3_X1   g120(.A1(new_n315), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n319), .B1(new_n315), .B2(new_n321), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G120gat), .B(G148gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(G176gat), .B(G204gat), .ZN(new_n326));
  XOR2_X1   g125(.A(new_n325), .B(new_n326), .Z(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n237), .A2(new_n280), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n280), .B1(new_n235), .B2(new_n234), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT10), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n237), .A2(KEYINPUT10), .A3(new_n281), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(G230gat), .A2(G233gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n330), .B1(new_n237), .B2(new_n280), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(new_n337), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n328), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT100), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n343), .B1(new_n332), .B2(new_n334), .ZN(new_n344));
  OAI211_X1 g143(.A(KEYINPUT100), .B(new_n333), .C1(new_n339), .C2(KEYINPUT10), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n344), .A2(new_n336), .A3(new_n345), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n341), .A2(new_n328), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n342), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n264), .A2(new_n324), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT101), .ZN(new_n351));
  OR2_X1    g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n351), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G197gat), .B(G204gat), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT22), .ZN(new_n356));
  INV_X1    g155(.A(G211gat), .ZN(new_n357));
  INV_X1    g156(.A(G218gat), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(G211gat), .B(G218gat), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n361), .A2(new_n355), .A3(new_n359), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT69), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n363), .A2(KEYINPUT69), .A3(new_n364), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(G226gat), .A2(G233gat), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n371), .A2(KEYINPUT29), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT25), .ZN(new_n373));
  NOR2_X1   g172(.A1(G183gat), .A2(G190gat), .ZN(new_n374));
  AND2_X1   g173(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n374), .B1(new_n375), .B2(G190gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(G183gat), .A2(G190gat), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT24), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT65), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n377), .A2(KEYINPUT65), .A3(new_n378), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n376), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(G169gat), .A2(G176gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(G169gat), .A2(G176gat), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n384), .B1(new_n385), .B2(KEYINPUT23), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT23), .ZN(new_n387));
  NOR3_X1   g186(.A1(new_n387), .A2(G169gat), .A3(G176gat), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n373), .B1(new_n383), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT27), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n391), .A2(G183gat), .ZN(new_n392));
  INV_X1    g191(.A(G183gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n393), .A2(KEYINPUT27), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT66), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(KEYINPUT27), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n391), .A2(G183gat), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT66), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT28), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n400), .A2(G190gat), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n395), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(G190gat), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n396), .A2(new_n397), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n400), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT67), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n385), .A2(new_n407), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n408), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n409));
  NOR4_X1   g208(.A1(KEYINPUT67), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n409), .A2(new_n411), .B1(G183gat), .B2(G190gat), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n390), .B1(new_n406), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT64), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n414), .B1(new_n386), .B2(new_n388), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n385), .A2(KEYINPUT23), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n387), .B1(G169gat), .B2(G176gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n414), .A2(new_n373), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n416), .A2(new_n417), .A3(new_n384), .A4(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n376), .A2(new_n379), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n415), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n372), .B1(new_n413), .B2(new_n421), .ZN(new_n422));
  NOR3_X1   g221(.A1(KEYINPUT67), .A2(G169gat), .A3(G176gat), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT26), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n384), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n377), .B1(new_n425), .B2(new_n410), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n426), .B1(new_n405), .B2(new_n402), .ZN(new_n427));
  AND3_X1   g226(.A1(new_n415), .A2(new_n419), .A3(new_n420), .ZN(new_n428));
  NOR4_X1   g227(.A1(new_n427), .A2(new_n428), .A3(new_n390), .A4(new_n371), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n369), .B1(new_n422), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n367), .A2(new_n368), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n406), .A2(new_n412), .ZN(new_n432));
  INV_X1    g231(.A(new_n390), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n432), .A2(new_n433), .A3(new_n421), .A4(new_n370), .ZN(new_n434));
  NOR3_X1   g233(.A1(new_n427), .A2(new_n428), .A3(new_n390), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n431), .B(new_n434), .C1(new_n435), .C2(new_n372), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n430), .A2(KEYINPUT70), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT70), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n438), .B(new_n369), .C1(new_n422), .C2(new_n429), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G8gat), .B(G36gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(G64gat), .B(G92gat), .ZN(new_n442));
  XOR2_X1   g241(.A(new_n441), .B(new_n442), .Z(new_n443));
  NAND2_X1  g242(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n443), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n437), .A2(new_n445), .A3(new_n439), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n444), .A2(KEYINPUT30), .A3(new_n446), .ZN(new_n447));
  AOI211_X1 g246(.A(KEYINPUT30), .B(new_n445), .C1(new_n437), .C2(new_n439), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(G225gat), .A2(G233gat), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT1), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT68), .ZN(new_n454));
  INV_X1    g253(.A(G113gat), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n454), .A2(new_n455), .A3(G120gat), .ZN(new_n456));
  INV_X1    g255(.A(G134gat), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(G127gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n243), .A2(G134gat), .ZN(new_n459));
  AND4_X1   g258(.A1(new_n453), .A2(new_n456), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(G113gat), .B(G120gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT68), .ZN(new_n462));
  INV_X1    g261(.A(G120gat), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(G113gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n455), .A2(G120gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(new_n453), .ZN(new_n467));
  XNOR2_X1  g266(.A(G127gat), .B(G134gat), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  AOI22_X1  g268(.A1(new_n460), .A2(new_n462), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(G155gat), .ZN(new_n471));
  INV_X1    g270(.A(G162gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(G155gat), .A2(G162gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(KEYINPUT2), .ZN(new_n477));
  XNOR2_X1  g276(.A(G141gat), .B(G148gat), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT71), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(G148gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(G141gat), .ZN(new_n482));
  INV_X1    g281(.A(G141gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(G148gat), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n482), .A2(new_n484), .A3(new_n479), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n476), .B1(new_n480), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n483), .A2(KEYINPUT72), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT72), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(G141gat), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(new_n490), .A3(G148gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n482), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n474), .B1(new_n473), .B2(KEYINPUT2), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n487), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n470), .B1(new_n495), .B2(KEYINPUT3), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n483), .A2(G148gat), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n481), .A2(G141gat), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT71), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n499), .A2(new_n485), .A3(new_n477), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n500), .A2(new_n476), .B1(new_n492), .B2(new_n493), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT3), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n452), .B1(new_n496), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n470), .A2(new_n487), .A3(new_n494), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT76), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT4), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n501), .A2(new_n508), .A3(new_n470), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n506), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT5), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n505), .A2(KEYINPUT76), .A3(KEYINPUT4), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n504), .A2(new_n510), .A3(new_n511), .A4(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT73), .ZN(new_n514));
  AND3_X1   g313(.A1(new_n506), .A2(new_n514), .A3(new_n509), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n501), .A2(KEYINPUT73), .A3(new_n508), .A4(new_n470), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n466), .A2(new_n454), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n468), .A2(new_n453), .A3(new_n456), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n461), .A2(KEYINPUT1), .ZN(new_n519));
  OAI22_X1  g318(.A1(new_n517), .A2(new_n518), .B1(new_n519), .B2(new_n468), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n520), .B1(new_n501), .B2(new_n502), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n474), .A2(KEYINPUT2), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n482), .A2(new_n484), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n522), .B1(new_n523), .B2(KEYINPUT71), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n475), .B1(new_n524), .B2(new_n485), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n475), .A2(new_n477), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n526), .B1(new_n482), .B2(new_n491), .ZN(new_n527));
  NOR3_X1   g326(.A1(new_n525), .A2(new_n527), .A3(KEYINPUT3), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n451), .B(new_n516), .C1(new_n521), .C2(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n515), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n520), .B1(new_n525), .B2(new_n527), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT74), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(new_n505), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n495), .A2(KEYINPUT74), .A3(new_n520), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n533), .A2(new_n452), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT5), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n513), .B1(new_n530), .B2(new_n536), .ZN(new_n537));
  XOR2_X1   g336(.A(G1gat), .B(G29gat), .Z(new_n538));
  XNOR2_X1  g337(.A(KEYINPUT75), .B(KEYINPUT0), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G57gat), .B(G85gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n537), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n542), .B(new_n513), .C1(new_n530), .C2(new_n536), .ZN(new_n545));
  XNOR2_X1  g344(.A(KEYINPUT77), .B(KEYINPUT6), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n546), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n537), .A2(new_n543), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n450), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT29), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n431), .B1(new_n552), .B2(new_n503), .ZN(new_n553));
  INV_X1    g352(.A(G228gat), .ZN(new_n554));
  INV_X1    g353(.A(G233gat), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n363), .A2(KEYINPUT78), .A3(new_n364), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n361), .B1(new_n359), .B2(new_n355), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT78), .ZN(new_n560));
  AOI21_X1  g359(.A(KEYINPUT29), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT3), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n557), .B1(new_n562), .B2(new_n501), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n553), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT29), .B1(new_n363), .B2(new_n364), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n502), .B1(new_n566), .B2(KEYINPUT79), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(KEYINPUT79), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n501), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n556), .B1(new_n570), .B2(new_n553), .ZN(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT31), .B(G50gat), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n565), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G78gat), .B(G106gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(G22gat), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n369), .B1(KEYINPUT29), .B2(new_n528), .ZN(new_n577));
  INV_X1    g376(.A(new_n569), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n495), .B1(new_n578), .B2(new_n567), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n557), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n572), .B1(new_n580), .B2(new_n564), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n574), .A2(new_n576), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n576), .B1(new_n574), .B2(new_n581), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n551), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT36), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n432), .A2(new_n433), .A3(new_n421), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(new_n520), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n413), .A2(new_n470), .A3(new_n421), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G227gat), .A2(G233gat), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g392(.A(KEYINPUT34), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT34), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n589), .A2(new_n590), .A3(new_n595), .A4(new_n592), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(G15gat), .B(G43gat), .Z(new_n598));
  XNOR2_X1  g397(.A(G71gat), .B(G99gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n591), .A2(new_n593), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT33), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n597), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n602), .A2(KEYINPUT32), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n592), .B1(new_n589), .B2(new_n590), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n600), .B1(new_n608), .B2(KEYINPUT33), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n609), .A2(new_n594), .A3(new_n596), .ZN(new_n610));
  AND3_X1   g409(.A1(new_n605), .A2(new_n607), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n607), .B1(new_n605), .B2(new_n610), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n587), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n605), .A2(new_n610), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(new_n606), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n605), .A2(new_n607), .A3(new_n610), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n615), .A2(KEYINPUT36), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n586), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT81), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT40), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n533), .A2(new_n534), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(new_n451), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT80), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n623), .A2(new_n624), .A3(KEYINPUT39), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n496), .A2(new_n503), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n510), .A2(new_n626), .A3(new_n512), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(new_n452), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n452), .B1(new_n533), .B2(new_n534), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT39), .ZN(new_n630));
  OAI21_X1  g429(.A(KEYINPUT80), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AND3_X1   g430(.A1(new_n625), .A2(new_n628), .A3(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n627), .A2(new_n630), .A3(new_n452), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(new_n542), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n621), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n625), .A2(new_n628), .A3(new_n631), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n636), .A2(KEYINPUT40), .A3(new_n542), .A4(new_n633), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n635), .A2(new_n544), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n446), .A2(KEYINPUT30), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n445), .B1(new_n437), .B2(new_n439), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n641), .A2(new_n448), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n620), .B1(new_n638), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n635), .A2(new_n544), .A3(new_n637), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n644), .A2(new_n450), .A3(KEYINPUT81), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n547), .A2(new_n549), .A3(new_n444), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT37), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n440), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT82), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n440), .A2(KEYINPUT82), .A3(new_n648), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n443), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n430), .A2(new_n436), .ZN(new_n654));
  AOI21_X1  g453(.A(KEYINPUT38), .B1(new_n654), .B2(KEYINPUT37), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n647), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n437), .A2(KEYINPUT37), .A3(new_n439), .ZN(new_n657));
  AOI21_X1  g456(.A(KEYINPUT82), .B1(new_n440), .B2(new_n648), .ZN(new_n658));
  AOI211_X1 g457(.A(new_n650), .B(KEYINPUT37), .C1(new_n437), .C2(new_n439), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n445), .B(new_n657), .C1(new_n658), .C2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(KEYINPUT38), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n585), .B1(new_n656), .B2(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n619), .B1(new_n646), .B2(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n611), .A2(new_n612), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n664), .A2(new_n550), .A3(new_n584), .A4(new_n450), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(KEYINPUT35), .ZN(new_n666));
  AND3_X1   g465(.A1(new_n584), .A2(new_n615), .A3(new_n616), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT35), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n667), .A2(new_n668), .A3(new_n550), .A4(new_n450), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(KEYINPUT83), .B1(new_n663), .B2(new_n670), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n445), .B(new_n655), .C1(new_n658), .C2(new_n659), .ZN(new_n672));
  INV_X1    g471(.A(new_n647), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n661), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT81), .B1(new_n644), .B2(new_n450), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n636), .A2(new_n542), .A3(new_n633), .ZN(new_n676));
  AOI22_X1  g475(.A1(new_n676), .A2(new_n621), .B1(new_n543), .B2(new_n537), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n642), .A2(new_n620), .A3(new_n637), .A4(new_n677), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n674), .A2(new_n584), .A3(new_n675), .A4(new_n678), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n586), .A2(new_n618), .ZN(new_n680));
  AOI22_X1  g479(.A1(new_n679), .A2(new_n680), .B1(new_n666), .B2(new_n669), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT83), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n671), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT90), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n254), .B(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n306), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n686), .B1(new_n687), .B2(new_n304), .ZN(new_n688));
  NAND2_X1  g487(.A1(G229gat), .A2(G233gat), .ZN(new_n689));
  INV_X1    g488(.A(new_n254), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n308), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n688), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT18), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n308), .B(new_n690), .ZN(new_n694));
  XOR2_X1   g493(.A(new_n689), .B(KEYINPUT13), .Z(new_n695));
  AOI22_X1  g494(.A1(new_n692), .A2(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(G113gat), .B(G141gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(G197gat), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT11), .B(G169gat), .Z(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XOR2_X1   g499(.A(new_n700), .B(KEYINPUT12), .Z(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n688), .A2(KEYINPUT18), .A3(new_n689), .A4(new_n691), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n696), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n702), .B1(new_n696), .B2(new_n703), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n684), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT91), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n684), .A2(KEYINPUT91), .A3(new_n708), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n354), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n550), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT102), .B(G1gat), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1324gat));
  NAND2_X1  g516(.A1(new_n713), .A2(new_n642), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT42), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(KEYINPUT103), .ZN(new_n720));
  XOR2_X1   g519(.A(KEYINPUT16), .B(G8gat), .Z(new_n721));
  MUX2_X1   g520(.A(KEYINPUT103), .B(new_n720), .S(new_n721), .Z(new_n722));
  NOR2_X1   g521(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n718), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n719), .B1(new_n724), .B2(new_n721), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n718), .A2(G8gat), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n723), .B1(new_n725), .B2(new_n726), .ZN(G1325gat));
  INV_X1    g526(.A(G15gat), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n713), .A2(new_n728), .A3(new_n664), .ZN(new_n729));
  INV_X1    g528(.A(new_n618), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n713), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n729), .B1(new_n731), .B2(new_n728), .ZN(G1326gat));
  AOI211_X1 g531(.A(new_n584), .B(new_n354), .C1(new_n711), .C2(new_n712), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT43), .B(G22gat), .Z(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(G1327gat));
  INV_X1    g534(.A(new_n349), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n264), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n324), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n739), .B1(new_n711), .B2(new_n712), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n550), .A2(G29gat), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OR2_X1    g541(.A1(new_n742), .A2(KEYINPUT45), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(KEYINPUT45), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n324), .B1(new_n671), .B2(new_n683), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT44), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n679), .A2(new_n680), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n666), .A2(new_n669), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT104), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n681), .A2(KEYINPUT104), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n324), .A2(KEYINPUT44), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  OAI22_X1  g554(.A1(new_n745), .A2(new_n746), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n737), .A2(new_n708), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(G29gat), .B1(new_n759), .B2(new_n550), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n743), .A2(new_n744), .A3(new_n760), .ZN(G1328gat));
  INV_X1    g560(.A(G36gat), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n740), .A2(new_n762), .A3(new_n642), .ZN(new_n763));
  OR2_X1    g562(.A1(new_n763), .A2(KEYINPUT46), .ZN(new_n764));
  OAI21_X1  g563(.A(G36gat), .B1(new_n759), .B2(new_n450), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(KEYINPUT46), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(G1329gat));
  NOR2_X1   g566(.A1(new_n618), .A2(new_n284), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n756), .A2(new_n758), .A3(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT47), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n769), .B1(KEYINPUT105), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n740), .A2(new_n664), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n771), .B1(new_n284), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n770), .A2(KEYINPUT105), .ZN(new_n774));
  XOR2_X1   g573(.A(new_n774), .B(KEYINPUT106), .Z(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n773), .B(new_n776), .ZN(G1330gat));
  INV_X1    g576(.A(new_n759), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n778), .A2(new_n283), .A3(new_n585), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n740), .A2(new_n585), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n779), .B1(new_n780), .B2(new_n283), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g581(.A1(new_n264), .A2(new_n324), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n783), .A2(new_n708), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n736), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(KEYINPUT107), .ZN(new_n786));
  INV_X1    g585(.A(new_n753), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(new_n550), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(new_n210), .ZN(G1332gat));
  NOR2_X1   g589(.A1(new_n788), .A2(new_n450), .ZN(new_n791));
  NOR2_X1   g590(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n792));
  AND2_X1   g591(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n794), .B1(new_n791), .B2(new_n792), .ZN(G1333gat));
  INV_X1    g594(.A(G71gat), .ZN(new_n796));
  INV_X1    g595(.A(new_n664), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n796), .B1(new_n788), .B2(new_n797), .ZN(new_n798));
  NOR4_X1   g597(.A1(new_n788), .A2(KEYINPUT108), .A3(new_n796), .A4(new_n618), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT108), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n786), .A2(new_n787), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n618), .A2(new_n796), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n798), .B1(new_n799), .B2(new_n803), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n804), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g604(.A1(new_n801), .A2(new_n585), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g606(.A1(new_n269), .A2(new_n271), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n264), .A2(new_n708), .A3(new_n349), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n756), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n808), .B1(new_n810), .B2(new_n550), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n258), .A2(new_n263), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n813), .A2(new_n738), .A3(new_n707), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n812), .B1(new_n681), .B2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT109), .ZN(new_n816));
  INV_X1    g615(.A(new_n814), .ZN(new_n817));
  OAI211_X1 g616(.A(KEYINPUT51), .B(new_n817), .C1(new_n663), .C2(new_n670), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n815), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  OAI211_X1 g618(.A(KEYINPUT109), .B(new_n812), .C1(new_n681), .C2(new_n814), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n821), .A2(new_n349), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n822), .A2(new_n714), .A3(new_n269), .A4(new_n271), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n811), .A2(new_n823), .ZN(G1336gat));
  NOR3_X1   g623(.A1(new_n349), .A2(G92gat), .A3(new_n450), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n819), .A2(new_n820), .A3(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT111), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n819), .A2(KEYINPUT111), .A3(new_n820), .A4(new_n825), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT52), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT112), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n756), .A2(new_n833), .A3(new_n642), .A4(new_n809), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n756), .A2(new_n642), .A3(new_n809), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n270), .B1(new_n835), .B2(KEYINPUT112), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n832), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n815), .A2(new_n818), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n825), .ZN(new_n839));
  XOR2_X1   g638(.A(new_n839), .B(KEYINPUT110), .Z(new_n840));
  NAND2_X1  g639(.A1(new_n835), .A2(G92gat), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n831), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(KEYINPUT113), .B1(new_n837), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n835), .A2(KEYINPUT112), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n844), .A2(new_n834), .A3(G92gat), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT52), .B1(new_n828), .B2(new_n829), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n840), .A2(new_n841), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(KEYINPUT52), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT113), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n847), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n843), .A2(new_n851), .ZN(G1337gat));
  OAI21_X1  g651(.A(G99gat), .B1(new_n810), .B2(new_n618), .ZN(new_n853));
  OR3_X1    g652(.A1(new_n797), .A2(G99gat), .A3(new_n349), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n853), .B1(new_n821), .B2(new_n854), .ZN(G1338gat));
  XNOR2_X1  g654(.A(KEYINPUT114), .B(G106gat), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n856), .B1(new_n810), .B2(new_n584), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n584), .A2(G106gat), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n838), .A2(new_n736), .A3(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT53), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT115), .ZN(new_n862));
  AOI21_X1  g661(.A(KEYINPUT53), .B1(new_n822), .B2(new_n859), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n857), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n862), .B1(new_n857), .B2(new_n863), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n861), .B1(new_n864), .B2(new_n865), .ZN(G1339gat));
  INV_X1    g665(.A(KEYINPUT55), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n868));
  AOI211_X1 g667(.A(new_n867), .B(new_n327), .C1(new_n338), .C2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n868), .B1(new_n335), .B2(new_n337), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT116), .ZN(new_n871));
  AND3_X1   g670(.A1(new_n346), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n871), .B1(new_n346), .B2(new_n870), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n869), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT117), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n869), .B(KEYINPUT117), .C1(new_n872), .C2(new_n873), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n327), .B1(new_n338), .B2(new_n868), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n879), .B1(new_n872), .B2(new_n873), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n867), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n878), .A2(new_n708), .A3(new_n348), .A4(new_n881), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n694), .A2(new_n695), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n689), .B1(new_n688), .B2(new_n691), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n700), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n704), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n886), .A2(new_n349), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n738), .B1(new_n882), .B2(new_n888), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n704), .B(new_n885), .C1(new_n322), .C2(new_n323), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n890), .B1(new_n867), .B2(new_n880), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n348), .A3(new_n878), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n813), .B1(new_n889), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n784), .A2(new_n349), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n550), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n896), .A2(new_n450), .A3(new_n667), .ZN(new_n897));
  AOI21_X1  g696(.A(G113gat), .B1(new_n897), .B2(new_n708), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n585), .B1(new_n894), .B2(new_n895), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n899), .A2(new_n714), .A3(new_n450), .A4(new_n664), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n900), .A2(new_n455), .A3(new_n707), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n898), .A2(new_n901), .ZN(G1340gat));
  NAND3_X1  g701(.A1(new_n897), .A2(new_n463), .A3(new_n736), .ZN(new_n903));
  OAI21_X1  g702(.A(G120gat), .B1(new_n900), .B2(new_n349), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT118), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n904), .A2(new_n905), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n903), .B1(new_n906), .B2(new_n907), .ZN(G1341gat));
  NAND3_X1  g707(.A1(new_n897), .A2(new_n243), .A3(new_n264), .ZN(new_n909));
  OAI21_X1  g708(.A(G127gat), .B1(new_n900), .B2(new_n813), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(G1342gat));
  OAI21_X1  g710(.A(G134gat), .B1(new_n900), .B2(new_n324), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n897), .A2(new_n457), .A3(new_n738), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n913), .A2(KEYINPUT119), .A3(KEYINPUT56), .ZN(new_n914));
  AOI21_X1  g713(.A(KEYINPUT119), .B1(new_n913), .B2(KEYINPUT56), .ZN(new_n915));
  OAI221_X1 g714(.A(new_n912), .B1(KEYINPUT56), .B2(new_n913), .C1(new_n914), .C2(new_n915), .ZN(G1343gat));
  NOR2_X1   g715(.A1(new_n730), .A2(new_n584), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n896), .A2(new_n450), .A3(new_n917), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n918), .A2(new_n483), .A3(new_n708), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n919), .A2(KEYINPUT58), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n488), .A2(new_n490), .ZN(new_n921));
  INV_X1    g720(.A(new_n895), .ZN(new_n922));
  INV_X1    g721(.A(new_n348), .ZN(new_n923));
  AOI211_X1 g722(.A(new_n923), .B(new_n707), .C1(new_n876), .C2(new_n877), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT120), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n880), .A2(new_n925), .ZN(new_n926));
  OAI211_X1 g725(.A(KEYINPUT120), .B(new_n879), .C1(new_n872), .C2(new_n873), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n926), .A2(new_n867), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n887), .B1(new_n924), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n892), .B1(new_n929), .B2(new_n738), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n922), .B1(new_n930), .B2(new_n813), .ZN(new_n931));
  OAI21_X1  g730(.A(KEYINPUT57), .B1(new_n931), .B2(new_n584), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n894), .A2(new_n895), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT57), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n933), .A2(new_n934), .A3(new_n585), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n730), .A2(new_n550), .A3(new_n642), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n932), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n921), .B1(new_n937), .B2(new_n707), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n920), .A2(new_n938), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n928), .A2(new_n878), .A3(new_n708), .A4(new_n348), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n738), .B1(new_n940), .B2(new_n888), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n813), .B1(new_n941), .B2(new_n893), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n584), .B1(new_n942), .B2(new_n895), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n936), .B1(new_n943), .B2(new_n934), .ZN(new_n944));
  AOI211_X1 g743(.A(KEYINPUT57), .B(new_n584), .C1(new_n894), .C2(new_n895), .ZN(new_n945));
  OAI21_X1  g744(.A(KEYINPUT121), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT121), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n932), .A2(new_n947), .A3(new_n935), .A4(new_n936), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n946), .A2(new_n708), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n919), .B1(new_n949), .B2(new_n921), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT58), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n939), .B1(new_n950), .B2(new_n951), .ZN(G1344gat));
  NAND3_X1  g751(.A1(new_n946), .A2(new_n736), .A3(new_n948), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n481), .A2(KEYINPUT59), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n352), .A2(new_n707), .A3(new_n353), .ZN(new_n956));
  AOI211_X1 g755(.A(KEYINPUT57), .B(new_n584), .C1(new_n942), .C2(new_n956), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n934), .B1(new_n933), .B2(new_n585), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n936), .A2(new_n736), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  OAI21_X1  g759(.A(KEYINPUT59), .B1(new_n960), .B2(new_n481), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n955), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n918), .A2(new_n481), .A3(new_n736), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(G1345gat));
  AOI21_X1  g763(.A(G155gat), .B1(new_n918), .B2(new_n264), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n946), .A2(new_n948), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n813), .A2(new_n471), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n967), .B(KEYINPUT122), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n965), .B1(new_n966), .B2(new_n968), .ZN(G1346gat));
  AOI21_X1  g768(.A(G162gat), .B1(new_n918), .B2(new_n738), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n324), .A2(new_n472), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n970), .B1(new_n966), .B2(new_n971), .ZN(G1347gat));
  AOI21_X1  g771(.A(new_n714), .B1(new_n894), .B2(new_n895), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n973), .A2(new_n642), .A3(new_n667), .ZN(new_n974));
  AOI21_X1  g773(.A(G169gat), .B1(new_n974), .B2(new_n708), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n714), .A2(new_n450), .ZN(new_n976));
  AND3_X1   g775(.A1(new_n899), .A2(new_n664), .A3(new_n976), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n708), .A2(G169gat), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n975), .B1(new_n977), .B2(new_n978), .ZN(G1348gat));
  AOI21_X1  g778(.A(G176gat), .B1(new_n974), .B2(new_n736), .ZN(new_n980));
  AND2_X1   g779(.A1(new_n736), .A2(G176gat), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n980), .B1(new_n977), .B2(new_n981), .ZN(G1349gat));
  NAND2_X1  g781(.A1(new_n977), .A2(new_n264), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n983), .A2(G183gat), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT123), .ZN(new_n985));
  NAND4_X1  g784(.A1(new_n974), .A2(new_n395), .A3(new_n399), .A4(new_n264), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n987), .A2(KEYINPUT60), .ZN(new_n988));
  INV_X1    g787(.A(KEYINPUT60), .ZN(new_n989));
  NAND4_X1  g788(.A1(new_n984), .A2(new_n985), .A3(new_n989), .A4(new_n986), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n988), .A2(new_n990), .ZN(G1350gat));
  NAND3_X1  g790(.A1(new_n974), .A2(new_n403), .A3(new_n738), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n738), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n993), .A2(G190gat), .ZN(new_n994));
  AND2_X1   g793(.A1(new_n994), .A2(KEYINPUT61), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n994), .A2(KEYINPUT61), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n992), .B1(new_n995), .B2(new_n996), .ZN(G1351gat));
  NAND2_X1  g796(.A1(new_n917), .A2(new_n642), .ZN(new_n998));
  XOR2_X1   g797(.A(new_n998), .B(KEYINPUT124), .Z(new_n999));
  AND2_X1   g798(.A1(new_n973), .A2(new_n999), .ZN(new_n1000));
  XOR2_X1   g799(.A(KEYINPUT125), .B(G197gat), .Z(new_n1001));
  NAND3_X1  g800(.A1(new_n1000), .A2(new_n708), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n618), .A2(new_n976), .ZN(new_n1003));
  OR3_X1    g802(.A1(new_n957), .A2(new_n958), .A3(new_n1003), .ZN(new_n1004));
  NOR2_X1   g803(.A1(new_n1004), .A2(new_n707), .ZN(new_n1005));
  OAI21_X1  g804(.A(new_n1002), .B1(new_n1005), .B2(new_n1001), .ZN(G1352gat));
  OAI21_X1  g805(.A(G204gat), .B1(new_n1004), .B2(new_n349), .ZN(new_n1007));
  INV_X1    g806(.A(KEYINPUT126), .ZN(new_n1008));
  AOI211_X1 g807(.A(G204gat), .B(new_n349), .C1(new_n1008), .C2(KEYINPUT62), .ZN(new_n1009));
  NAND3_X1  g808(.A1(new_n973), .A2(new_n999), .A3(new_n1009), .ZN(new_n1010));
  NOR2_X1   g809(.A1(new_n1008), .A2(KEYINPUT62), .ZN(new_n1011));
  XNOR2_X1  g810(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  NAND3_X1  g811(.A1(new_n1007), .A2(new_n1012), .A3(KEYINPUT127), .ZN(new_n1013));
  INV_X1    g812(.A(KEYINPUT127), .ZN(new_n1014));
  INV_X1    g813(.A(new_n1012), .ZN(new_n1015));
  INV_X1    g814(.A(G204gat), .ZN(new_n1016));
  NOR3_X1   g815(.A1(new_n957), .A2(new_n958), .A3(new_n1003), .ZN(new_n1017));
  AOI21_X1  g816(.A(new_n1016), .B1(new_n1017), .B2(new_n736), .ZN(new_n1018));
  OAI21_X1  g817(.A(new_n1014), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n1013), .A2(new_n1019), .ZN(G1353gat));
  NAND3_X1  g819(.A1(new_n1000), .A2(new_n357), .A3(new_n264), .ZN(new_n1021));
  NAND2_X1  g820(.A1(new_n1017), .A2(new_n264), .ZN(new_n1022));
  AND3_X1   g821(.A1(new_n1022), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1023));
  AOI21_X1  g822(.A(KEYINPUT63), .B1(new_n1022), .B2(G211gat), .ZN(new_n1024));
  OAI21_X1  g823(.A(new_n1021), .B1(new_n1023), .B2(new_n1024), .ZN(G1354gat));
  OAI21_X1  g824(.A(G218gat), .B1(new_n1004), .B2(new_n324), .ZN(new_n1026));
  NAND3_X1  g825(.A1(new_n1000), .A2(new_n358), .A3(new_n738), .ZN(new_n1027));
  NAND2_X1  g826(.A1(new_n1026), .A2(new_n1027), .ZN(G1355gat));
endmodule


