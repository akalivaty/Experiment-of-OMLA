//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 0 1 1 0 0 0 1 1 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n546, new_n547, new_n548, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n564, new_n565, new_n566, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n611,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT66), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI21_X1  g033(.A(new_n457), .B1(new_n458), .B2(new_n453), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT67), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n463), .A2(new_n465), .A3(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n464), .A2(G2105), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n472), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n462), .A2(KEYINPUT68), .A3(G2104), .ZN(new_n474));
  NAND4_X1  g049(.A1(new_n473), .A2(new_n474), .A3(new_n461), .A4(new_n465), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G137), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n471), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  NAND4_X1  g054(.A1(new_n473), .A2(new_n474), .A3(G2105), .A4(new_n465), .ZN(new_n480));
  INV_X1    g055(.A(G124), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n461), .A2(G112), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  OAI22_X1  g058(.A1(new_n480), .A2(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n484), .B1(new_n476), .B2(G136), .ZN(G162));
  NOR2_X1   g060(.A1(new_n461), .A2(G114), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AND4_X1   g063(.A1(G2105), .A2(new_n473), .A3(new_n474), .A4(new_n465), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(G126), .ZN(new_n490));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n473), .A2(new_n474), .A3(new_n492), .A4(new_n465), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  XNOR2_X1  g069(.A(KEYINPUT3), .B(G2104), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT69), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT69), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n495), .A2(new_n492), .A3(new_n497), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n490), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  NAND2_X1  g078(.A1(KEYINPUT70), .A2(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g081(.A1(KEYINPUT70), .A2(KEYINPUT5), .A3(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G62), .ZN(new_n509));
  NAND2_X1  g084(.A1(G75), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G651), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n511), .A2(KEYINPUT71), .A3(G651), .ZN(new_n515));
  OR2_X1    g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n506), .A2(new_n507), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n505), .B1(new_n516), .B2(new_n517), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n518), .A2(G88), .B1(new_n519), .B2(G50), .ZN(new_n520));
  AND3_X1   g095(.A1(new_n514), .A2(new_n515), .A3(new_n520), .ZN(G166));
  NAND2_X1  g096(.A1(new_n519), .A2(G51), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n522), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n518), .A2(G89), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(G168));
  NAND2_X1  g103(.A1(new_n519), .A2(G52), .ZN(new_n529));
  INV_X1    g104(.A(new_n518), .ZN(new_n530));
  XNOR2_X1  g105(.A(KEYINPUT72), .B(G90), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G651), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n532), .A2(new_n535), .ZN(G171));
  XNOR2_X1  g111(.A(KEYINPUT73), .B(G43), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n518), .A2(G81), .B1(new_n519), .B2(new_n537), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT74), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(new_n534), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND4_X1  g122(.A1(G319), .A2(G483), .A3(G661), .A4(new_n547), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT75), .ZN(G188));
  NAND2_X1  g124(.A1(G78), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(new_n507), .ZN(new_n551));
  AOI21_X1  g126(.A(G543), .B1(KEYINPUT70), .B2(KEYINPUT5), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(G65), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n550), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n555), .A2(G651), .B1(G91), .B2(new_n518), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n519), .A2(G53), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(KEYINPUT9), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n519), .A2(new_n559), .A3(G53), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n556), .A2(new_n561), .ZN(G299));
  INV_X1    g137(.A(G171), .ZN(G301));
  INV_X1    g138(.A(KEYINPUT76), .ZN(new_n564));
  NOR2_X1   g139(.A1(G168), .A2(new_n564), .ZN(new_n565));
  NOR3_X1   g140(.A1(new_n526), .A2(new_n527), .A3(KEYINPUT76), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n565), .A2(new_n566), .ZN(G286));
  NAND3_X1  g142(.A1(new_n514), .A2(new_n515), .A3(new_n520), .ZN(G303));
  OR3_X1    g143(.A1(new_n551), .A2(G74), .A3(new_n552), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n569), .A2(G651), .B1(G49), .B2(new_n519), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT77), .ZN(new_n571));
  AND3_X1   g146(.A1(new_n518), .A2(new_n571), .A3(G87), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n571), .B1(new_n518), .B2(G87), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n570), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT78), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OAI211_X1 g151(.A(new_n570), .B(KEYINPUT78), .C1(new_n572), .C2(new_n573), .ZN(new_n577));
  AND2_X1   g152(.A1(new_n576), .A2(new_n577), .ZN(G288));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n579), .B1(new_n506), .B2(new_n507), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT79), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n584), .B1(new_n580), .B2(new_n581), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n518), .A2(G86), .B1(new_n519), .B2(G48), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G305));
  AOI22_X1  g163(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n589), .A2(new_n534), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n518), .A2(G85), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n519), .A2(G47), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(G301), .A2(G868), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n518), .A2(G92), .ZN(new_n597));
  XOR2_X1   g172(.A(new_n597), .B(KEYINPUT10), .Z(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n553), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n601), .A2(G651), .B1(G54), .B2(new_n519), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n596), .B1(new_n604), .B2(G868), .ZN(G321));
  XOR2_X1   g180(.A(G321), .B(KEYINPUT80), .Z(G284));
  NOR2_X1   g181(.A1(G299), .A2(G868), .ZN(new_n607));
  INV_X1    g182(.A(G286), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G297));
  AOI21_X1  g184(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G280));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n604), .B1(new_n611), .B2(G860), .ZN(G148));
  INV_X1    g187(.A(G868), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n542), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n603), .A2(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(new_n613), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g192(.A(G123), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT82), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(new_n461), .B2(G111), .ZN(new_n620));
  OR2_X1    g195(.A1(G99), .A2(G2105), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n620), .A2(G2104), .A3(new_n621), .ZN(new_n622));
  NOR3_X1   g197(.A1(new_n619), .A2(new_n461), .A3(G111), .ZN(new_n623));
  OAI22_X1  g198(.A1(new_n480), .A2(new_n618), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n624), .B1(new_n476), .B2(G135), .ZN(new_n625));
  INV_X1    g200(.A(G2096), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n629));
  NOR3_X1   g204(.A1(new_n462), .A2(new_n464), .A3(G2105), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(KEYINPUT13), .B(G2100), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n627), .A2(new_n628), .A3(new_n633), .ZN(G156));
  INV_X1    g209(.A(KEYINPUT14), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2427), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2430), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n635), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(new_n638), .B2(new_n637), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2451), .B(G2454), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1341), .B(G1348), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n640), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(G14), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT83), .ZN(G401));
  INV_X1    g225(.A(KEYINPUT18), .ZN(new_n651));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  XNOR2_X1  g227(.A(G2067), .B(G2678), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n654), .A2(KEYINPUT17), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n652), .A2(new_n653), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n651), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2100), .ZN(new_n658));
  XOR2_X1   g233(.A(G2072), .B(G2078), .Z(new_n659));
  AOI21_X1  g234(.A(new_n659), .B1(new_n654), .B2(KEYINPUT18), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2096), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n658), .B(new_n661), .ZN(G227));
  XOR2_X1   g237(.A(G1971), .B(G1976), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  XOR2_X1   g239(.A(G1956), .B(G2474), .Z(new_n665));
  XOR2_X1   g240(.A(G1961), .B(G1966), .Z(new_n666));
  AND2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT20), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n665), .A2(new_n666), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n664), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n671), .B1(new_n664), .B2(new_n670), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1991), .B(G1996), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT84), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n675), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1981), .B(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(G229));
  MUX2_X1   g255(.A(G23), .B(new_n574), .S(G16), .Z(new_n681));
  XOR2_X1   g256(.A(KEYINPUT33), .B(G1976), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  MUX2_X1   g258(.A(G6), .B(G305), .S(G16), .Z(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT32), .B(G1981), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n683), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n684), .A2(new_n685), .ZN(new_n687));
  INV_X1    g262(.A(G1971), .ZN(new_n688));
  NAND2_X1  g263(.A1(G166), .A2(G16), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(G16), .B2(G22), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n687), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n686), .B(new_n691), .C1(new_n688), .C2(new_n690), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n692), .A2(KEYINPUT34), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(KEYINPUT34), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT35), .B(G1991), .Z(new_n695));
  NAND2_X1  g270(.A1(new_n476), .A2(G131), .ZN(new_n696));
  INV_X1    g271(.A(G95), .ZN(new_n697));
  AND3_X1   g272(.A1(new_n697), .A2(new_n461), .A3(KEYINPUT85), .ZN(new_n698));
  AOI21_X1  g273(.A(KEYINPUT85), .B1(new_n697), .B2(new_n461), .ZN(new_n699));
  OAI221_X1 g274(.A(G2104), .B1(G107), .B2(new_n461), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G119), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n696), .B(new_n700), .C1(new_n701), .C2(new_n480), .ZN(new_n702));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(G25), .A2(G29), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n695), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G24), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(new_n594), .B2(new_n707), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G1986), .ZN(new_n710));
  NOR3_X1   g285(.A1(new_n704), .A2(new_n705), .A3(new_n695), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g287(.A1(new_n693), .A2(new_n694), .A3(new_n706), .A4(new_n712), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT86), .B(KEYINPUT36), .Z(new_n714));
  OR2_X1    g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n714), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n707), .A2(G4), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(new_n604), .B2(new_n707), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(G1348), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT91), .B(KEYINPUT23), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n707), .A2(G20), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G299), .B2(G16), .ZN(new_n723));
  INV_X1    g298(.A(G1956), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n719), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G34), .ZN(new_n727));
  AOI21_X1  g302(.A(G29), .B1(new_n727), .B2(KEYINPUT24), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(KEYINPUT24), .B2(new_n727), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(new_n478), .B2(new_n703), .ZN(new_n730));
  INV_X1    g305(.A(G2084), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n707), .A2(G21), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G168), .B2(new_n707), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n703), .A2(G33), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT25), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n495), .A2(G127), .ZN(new_n738));
  NAND2_X1  g313(.A1(G115), .A2(G2104), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n737), .B1(new_n740), .B2(G2105), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n476), .A2(G139), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n735), .B1(new_n743), .B2(G29), .ZN(new_n744));
  INV_X1    g319(.A(G2072), .ZN(new_n745));
  OAI221_X1 g320(.A(new_n732), .B1(G1966), .B2(new_n734), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n744), .A2(new_n745), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n734), .A2(G1966), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT30), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n749), .A2(G28), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n703), .B1(new_n749), .B2(G28), .ZN(new_n751));
  AND2_X1   g326(.A1(KEYINPUT31), .A2(G11), .ZN(new_n752));
  NOR2_X1   g327(.A1(KEYINPUT31), .A2(G11), .ZN(new_n753));
  OAI22_X1  g328(.A1(new_n750), .A2(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n625), .B2(G29), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n730), .A2(new_n731), .ZN(new_n756));
  NAND4_X1  g331(.A1(new_n747), .A2(new_n748), .A3(new_n755), .A4(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n746), .A2(new_n757), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT89), .B(KEYINPUT28), .Z(new_n759));
  NAND2_X1  g334(.A1(new_n703), .A2(G26), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(KEYINPUT88), .B1(G104), .B2(G2105), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  NOR3_X1   g338(.A1(KEYINPUT88), .A2(G104), .A3(G2105), .ZN(new_n764));
  OAI221_X1 g339(.A(G2104), .B1(G116), .B2(new_n461), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G128), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n765), .B1(new_n766), .B2(new_n480), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n476), .A2(G140), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n761), .B1(new_n769), .B2(new_n703), .ZN(new_n770));
  INV_X1    g345(.A(G2067), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n707), .A2(G5), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G171), .B2(new_n707), .ZN(new_n774));
  INV_X1    g349(.A(G1961), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(G27), .A2(G29), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G164), .B2(G29), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n776), .B1(G2078), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G2078), .B2(new_n778), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n726), .A2(new_n758), .A3(new_n772), .A4(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(G16), .A2(G19), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n543), .B2(G16), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT87), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G1341), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n703), .A2(G35), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G162), .B2(new_n703), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT29), .Z(new_n788));
  INV_X1    g363(.A(G2090), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n703), .A2(G32), .ZN(new_n791));
  NAND3_X1  g366(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT26), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n792), .A2(new_n793), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n794), .A2(new_n795), .B1(G105), .B2(new_n469), .ZN(new_n796));
  INV_X1    g371(.A(G129), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n480), .B2(new_n797), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n476), .A2(G141), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n791), .B1(new_n800), .B2(new_n703), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT90), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT27), .B(G1996), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n788), .A2(new_n789), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n802), .A2(new_n804), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n790), .A2(new_n805), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  NOR3_X1   g383(.A1(new_n781), .A2(new_n785), .A3(new_n808), .ZN(new_n809));
  AND3_X1   g384(.A1(new_n715), .A2(new_n716), .A3(new_n809), .ZN(G311));
  NAND3_X1  g385(.A1(new_n715), .A2(new_n716), .A3(new_n809), .ZN(G150));
  AND2_X1   g386(.A1(G80), .A2(G543), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n508), .B2(G67), .ZN(new_n813));
  OR3_X1    g388(.A1(new_n813), .A2(KEYINPUT92), .A3(new_n534), .ZN(new_n814));
  OAI21_X1  g389(.A(KEYINPUT92), .B1(new_n813), .B2(new_n534), .ZN(new_n815));
  AOI22_X1  g390(.A1(new_n518), .A2(G93), .B1(new_n519), .B2(G55), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT93), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(new_n818), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G860), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT94), .B(KEYINPUT37), .Z(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n604), .A2(G559), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT38), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n819), .A2(new_n542), .A3(new_n820), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n543), .A2(new_n817), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n826), .B(new_n829), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n830), .A2(KEYINPUT39), .ZN(new_n831));
  INV_X1    g406(.A(G860), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n830), .B2(KEYINPUT39), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n824), .B1(new_n831), .B2(new_n833), .ZN(G145));
  XNOR2_X1  g409(.A(new_n625), .B(new_n478), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(G162), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT95), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n502), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n490), .A2(new_n501), .A3(KEYINPUT95), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n769), .ZN(new_n841));
  OAI21_X1  g416(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n842));
  INV_X1    g417(.A(G118), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n842), .B1(new_n843), .B2(G2105), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(new_n476), .B2(G142), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT98), .ZN(new_n846));
  AND3_X1   g421(.A1(new_n489), .A2(new_n846), .A3(G130), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n846), .B1(new_n489), .B2(G130), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n845), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n841), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n769), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n840), .B(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n849), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n800), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n743), .A2(KEYINPUT96), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT97), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n743), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n855), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n856), .A2(new_n855), .A3(new_n858), .ZN(new_n861));
  INV_X1    g436(.A(new_n702), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(KEYINPUT99), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT99), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n702), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n863), .A2(new_n631), .A3(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n631), .B1(new_n863), .B2(new_n865), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n860), .B(new_n861), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n868), .ZN(new_n870));
  INV_X1    g445(.A(new_n861), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n866), .B(new_n870), .C1(new_n871), .C2(new_n859), .ZN(new_n872));
  NAND4_X1  g447(.A1(new_n850), .A2(new_n854), .A3(new_n869), .A4(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  AOI22_X1  g449(.A1(new_n850), .A2(new_n854), .B1(new_n869), .B2(new_n872), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n836), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(KEYINPUT100), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n850), .A2(new_n854), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n869), .A2(new_n872), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(new_n873), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT100), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n881), .A2(new_n882), .A3(new_n836), .ZN(new_n883));
  AOI21_X1  g458(.A(G37), .B1(new_n877), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n836), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n880), .A2(new_n885), .A3(new_n873), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT101), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n884), .A2(KEYINPUT40), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(KEYINPUT40), .B1(new_n884), .B2(new_n887), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(G395));
  INV_X1    g465(.A(KEYINPUT108), .ZN(new_n891));
  XNOR2_X1  g466(.A(G166), .B(new_n574), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT104), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n594), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(KEYINPUT104), .B1(new_n590), .B2(new_n593), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n897));
  NAND2_X1  g472(.A1(G305), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n586), .A2(KEYINPUT105), .A3(new_n587), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n896), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n896), .B1(new_n898), .B2(new_n899), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n892), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT107), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n898), .A2(new_n899), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n905), .A2(new_n895), .A3(new_n894), .ZN(new_n906));
  XNOR2_X1  g481(.A(G303), .B(new_n574), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(new_n907), .A3(new_n900), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n903), .A2(new_n904), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(KEYINPUT42), .B1(new_n909), .B2(KEYINPUT106), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT106), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n903), .A2(new_n912), .A3(new_n908), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n913), .B1(KEYINPUT106), .B2(new_n909), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT42), .ZN(new_n915));
  OAI211_X1 g490(.A(new_n891), .B(new_n911), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n909), .A2(KEYINPUT106), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n903), .A2(new_n912), .A3(new_n908), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT108), .B1(new_n919), .B2(new_n910), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n829), .B(new_n615), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT103), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n603), .A2(G299), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n598), .A2(new_n561), .A3(new_n556), .A4(new_n602), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n924), .A2(KEYINPUT41), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(KEYINPUT41), .B1(new_n924), .B2(new_n925), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n922), .A2(new_n923), .A3(new_n928), .ZN(new_n929));
  NOR3_X1   g504(.A1(new_n921), .A2(new_n927), .A3(new_n926), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n924), .A2(KEYINPUT102), .A3(new_n925), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT102), .B1(new_n924), .B2(new_n925), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT103), .B1(new_n921), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n929), .B1(new_n930), .B2(new_n934), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n916), .A2(new_n920), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n935), .B1(new_n916), .B2(new_n920), .ZN(new_n937));
  OAI21_X1  g512(.A(G868), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n821), .A2(new_n613), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(G295));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n939), .ZN(G331));
  INV_X1    g516(.A(KEYINPUT43), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT109), .ZN(new_n943));
  NOR2_X1   g518(.A1(G171), .A2(G168), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n945), .B1(G286), .B2(G301), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n827), .A2(new_n946), .A3(new_n828), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n946), .B1(new_n827), .B2(new_n828), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n928), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n946), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n829), .A2(new_n951), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n952), .A2(new_n924), .A3(new_n925), .A4(new_n947), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n903), .A2(new_n908), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n950), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(G37), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n933), .A2(new_n952), .A3(new_n947), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n954), .B1(new_n950), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n943), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n959), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n961), .A2(KEYINPUT109), .A3(new_n956), .A4(new_n955), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n942), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n954), .B1(new_n950), .B2(new_n953), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n957), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT44), .B1(new_n963), .B2(new_n966), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n961), .A2(new_n942), .A3(new_n956), .A4(new_n955), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n968), .B1(new_n965), .B2(new_n942), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT44), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n967), .A2(new_n971), .ZN(G397));
  INV_X1    g547(.A(G1384), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n838), .A2(new_n973), .A3(new_n839), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT45), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n471), .A2(G40), .A3(new_n477), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT110), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT110), .ZN(new_n979));
  INV_X1    g554(.A(G137), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n475), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G40), .ZN(new_n982));
  NOR4_X1   g557(.A1(new_n981), .A2(new_n468), .A3(new_n982), .A4(new_n470), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n974), .A2(new_n979), .A3(new_n975), .A4(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n769), .B(new_n771), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n978), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT111), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n986), .B(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n978), .A2(new_n855), .A3(new_n984), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n976), .A2(new_n977), .ZN(new_n990));
  INV_X1    g565(.A(G1996), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AOI22_X1  g567(.A1(new_n989), .A2(new_n992), .B1(new_n991), .B2(new_n855), .ZN(new_n993));
  OAI21_X1  g568(.A(KEYINPUT112), .B1(new_n988), .B2(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n986), .B(KEYINPUT111), .ZN(new_n995));
  INV_X1    g570(.A(new_n993), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n862), .A2(new_n695), .ZN(new_n999));
  AND2_X1   g574(.A1(new_n862), .A2(new_n695), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n978), .B(new_n984), .C1(new_n999), .C2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n994), .A2(new_n998), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1986), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n594), .B(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1002), .B1(new_n990), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(G1384), .B1(new_n490), .B2(new_n501), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n983), .B1(new_n1006), .B2(KEYINPUT45), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT119), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1010), .A2(G2078), .ZN(new_n1011));
  AND3_X1   g586(.A1(new_n492), .A2(new_n497), .A3(new_n499), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n495), .A2(new_n1012), .B1(new_n493), .B2(KEYINPUT4), .ZN(new_n1013));
  INV_X1    g588(.A(G126), .ZN(new_n1014));
  OAI22_X1  g589(.A1(new_n480), .A2(new_n1014), .B1(new_n486), .B2(new_n487), .ZN(new_n1015));
  OAI211_X1 g590(.A(KEYINPUT45), .B(new_n973), .C1(new_n1013), .C2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT120), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n502), .A2(KEYINPUT120), .A3(KEYINPUT45), .A4(new_n973), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g595(.A(KEYINPUT119), .B(new_n983), .C1(new_n1006), .C2(KEYINPUT45), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1009), .A2(new_n1011), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n973), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n977), .B1(new_n1023), .B2(KEYINPUT50), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT50), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1006), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(new_n775), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1022), .A2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n838), .A2(KEYINPUT45), .A3(new_n973), .A4(new_n839), .ZN(new_n1030));
  INV_X1    g605(.A(G2078), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n977), .B1(new_n1023), .B2(new_n975), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n1010), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT125), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT125), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1033), .A2(new_n1036), .A3(new_n1010), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1029), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT126), .B1(new_n1038), .B2(G301), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT126), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1033), .A2(new_n1036), .A3(new_n1010), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1036), .B1(new_n1033), .B2(new_n1010), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1040), .B(G171), .C1(new_n1043), .C2(new_n1029), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1030), .A2(new_n983), .A3(new_n1011), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n1046), .A2(new_n976), .B1(new_n775), .B2(new_n1027), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1045), .A2(G301), .A3(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1039), .A2(new_n1044), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1027), .A2(new_n724), .ZN(new_n1052));
  NAND2_X1  g627(.A1(KEYINPUT121), .A2(KEYINPUT57), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT121), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT57), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AND3_X1   g631(.A1(G299), .A2(new_n1053), .A3(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1056), .B1(G299), .B2(new_n1053), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g634(.A(KEYINPUT56), .B(G2072), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1030), .A2(new_n1032), .A3(new_n1060), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1052), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1059), .B1(new_n1052), .B2(new_n1061), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT61), .ZN(new_n1064));
  OAI22_X1  g639(.A1(new_n1062), .A2(new_n1063), .B1(KEYINPUT123), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(KEYINPUT123), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OAI211_X1 g642(.A(KEYINPUT123), .B(new_n1064), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1030), .A2(new_n991), .A3(new_n1032), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1006), .A2(new_n983), .ZN(new_n1071));
  XOR2_X1   g646(.A(KEYINPUT58), .B(G1341), .Z(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  AOI211_X1 g648(.A(new_n1069), .B(new_n542), .C1(new_n1070), .C2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT122), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1075), .B1(new_n1071), .B2(G2067), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1006), .A2(new_n983), .A3(KEYINPUT122), .A4(new_n771), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(G1348), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n604), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G1348), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1027), .A2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1082), .A2(new_n603), .A3(new_n1077), .A4(new_n1076), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1074), .B1(new_n1084), .B2(KEYINPUT60), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT59), .B1(new_n1086), .B2(new_n543), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n603), .A2(KEYINPUT60), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1087), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1067), .A2(new_n1068), .A3(new_n1085), .A4(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1062), .A2(new_n1080), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1092), .A2(new_n1063), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1009), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1095));
  INV_X1    g670(.A(G1966), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1027), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n1095), .A2(new_n1096), .B1(new_n1097), .B2(new_n731), .ZN(new_n1098));
  INV_X1    g673(.A(G8), .ZN(new_n1099));
  NOR2_X1   g674(.A1(G168), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(KEYINPUT51), .B1(new_n1100), .B2(KEYINPUT124), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1097), .A2(new_n731), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(G168), .ZN(new_n1108));
  OAI211_X1 g683(.A(G8), .B(new_n1104), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1101), .B(new_n1103), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1102), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n688), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1114), .B1(new_n1027), .B2(G2090), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1024), .A2(KEYINPUT113), .A3(new_n789), .A4(new_n1026), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1113), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT55), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1099), .B1(KEYINPUT114), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(G303), .A2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1118), .A2(KEYINPUT114), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1121), .B(KEYINPUT115), .ZN(new_n1122));
  XOR2_X1   g697(.A(new_n1120), .B(new_n1122), .Z(new_n1123));
  NAND3_X1  g698(.A1(new_n1117), .A2(G8), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(G1976), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n576), .A2(new_n1125), .A3(new_n577), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT52), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1099), .B1(new_n1006), .B2(new_n983), .ZN(new_n1128));
  OR2_X1    g703(.A1(new_n574), .A2(new_n1125), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .A4(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1128), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(KEYINPUT52), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(G61), .B1(new_n551), .B2(new_n552), .ZN(new_n1134));
  AOI22_X1  g709(.A1(new_n1134), .A2(KEYINPUT79), .B1(G73), .B2(G543), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n534), .B1(new_n1135), .B2(new_n582), .ZN(new_n1136));
  INV_X1    g711(.A(new_n587), .ZN(new_n1137));
  OAI21_X1  g712(.A(G1981), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(G1981), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n586), .A2(new_n1139), .A3(new_n587), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT116), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1138), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(G305), .A2(KEYINPUT116), .A3(G1981), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT49), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(KEYINPUT117), .ZN(new_n1146));
  OR2_X1    g721(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1128), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1148), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1133), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1027), .A2(G2090), .ZN(new_n1151));
  AOI21_X1  g726(.A(G1971), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1152));
  OAI21_X1  g727(.A(G8), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1120), .B(new_n1122), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1124), .A2(new_n1150), .A3(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1111), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1050), .B1(new_n1038), .B2(G301), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1158), .B1(G301), .B2(new_n1159), .ZN(new_n1160));
  AND4_X1   g735(.A1(new_n1051), .A2(new_n1094), .A3(new_n1157), .A4(new_n1160), .ZN(new_n1161));
  XOR2_X1   g736(.A(new_n1140), .B(KEYINPUT118), .Z(new_n1162));
  NAND2_X1  g737(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1163));
  NOR2_X1   g738(.A1(G288), .A2(G1976), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1162), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1150), .ZN(new_n1166));
  OAI22_X1  g741(.A1(new_n1165), .A2(new_n1148), .B1(new_n1166), .B2(new_n1124), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT63), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1107), .A2(G8), .A3(new_n608), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1168), .B1(new_n1156), .B2(new_n1169), .ZN(new_n1170));
  NOR4_X1   g745(.A1(new_n1098), .A2(new_n1168), .A3(new_n1099), .A4(G286), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1117), .A2(G8), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(new_n1154), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1171), .A2(new_n1173), .A3(new_n1124), .A4(new_n1150), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1167), .B1(new_n1170), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1039), .A2(new_n1044), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1156), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT62), .ZN(new_n1178));
  OAI211_X1 g753(.A(new_n1176), .B(new_n1177), .C1(new_n1111), .C2(new_n1178), .ZN(new_n1179));
  AND2_X1   g754(.A1(new_n1111), .A2(new_n1178), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1175), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1005), .B1(new_n1161), .B2(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n992), .B(KEYINPUT46), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1183), .A2(new_n989), .A3(new_n986), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n1184), .B(KEYINPUT47), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n990), .A2(new_n1003), .A3(new_n594), .ZN(new_n1186));
  XOR2_X1   g761(.A(new_n1186), .B(KEYINPUT48), .Z(new_n1187));
  OAI21_X1  g762(.A(new_n1185), .B1(new_n1002), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n978), .A2(new_n984), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n994), .A2(new_n998), .A3(new_n1000), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n769), .A2(new_n771), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1189), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1188), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1182), .A2(new_n1193), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g769(.A1(new_n884), .A2(new_n887), .ZN(new_n1196));
  NOR2_X1   g770(.A1(G227), .A2(new_n459), .ZN(new_n1197));
  NAND2_X1  g771(.A1(new_n649), .A2(new_n1197), .ZN(new_n1198));
  XNOR2_X1  g772(.A(new_n1198), .B(KEYINPUT127), .ZN(new_n1199));
  NOR2_X1   g773(.A1(G229), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g774(.A1(new_n1196), .A2(new_n969), .A3(new_n1200), .ZN(G225));
  INV_X1    g775(.A(G225), .ZN(G308));
endmodule


