//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 0 0 1 1 1 0 1 0 0 1 0 0 1 0 0 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1324, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1390, new_n1391, new_n1392, new_n1393, new_n1394;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT0), .ZN(new_n206));
  OAI21_X1  g0006(.A(G50), .B1(G58), .B2(G68), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  AND2_X1   g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  NAND3_X1  g0009(.A1(new_n208), .A2(G20), .A3(new_n209), .ZN(new_n210));
  AND2_X1   g0010(.A1(KEYINPUT64), .A2(G77), .ZN(new_n211));
  NOR2_X1   g0011(.A1(KEYINPUT64), .A2(G77), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G244), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G58), .A2(G232), .ZN(new_n219));
  NAND4_X1  g0019(.A1(new_n216), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n203), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n206), .B(new_n210), .C1(KEYINPUT1), .C2(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n222), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XOR2_X1   g0023(.A(G226), .B(G232), .Z(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT66), .ZN(new_n225));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n227), .B(new_n228), .Z(new_n229));
  XOR2_X1   g0029(.A(G250), .B(G257), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT67), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n229), .B(new_n233), .Z(G358));
  XOR2_X1   g0034(.A(G87), .B(G97), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT68), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G351));
  XNOR2_X1  g0042(.A(KEYINPUT8), .B(G58), .ZN(new_n243));
  INV_X1    g0043(.A(new_n243), .ZN(new_n244));
  INV_X1    g0044(.A(G1), .ZN(new_n245));
  NAND3_X1  g0045(.A1(new_n245), .A2(G13), .A3(G20), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G20), .ZN(new_n249));
  OAI21_X1  g0049(.A(KEYINPUT72), .B1(new_n249), .B2(G1), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT72), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(new_n245), .A3(G20), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G1), .A2(G13), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g0056(.A(KEYINPUT71), .B1(new_n247), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NOR3_X1   g0058(.A1(new_n247), .A2(new_n256), .A3(KEYINPUT71), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n253), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n248), .B1(new_n260), .B2(new_n244), .ZN(new_n261));
  INV_X1    g0061(.A(new_n256), .ZN(new_n262));
  XNOR2_X1  g0062(.A(G58), .B(G68), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G20), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(KEYINPUT81), .A3(G159), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(KEYINPUT81), .B1(new_n265), .B2(G159), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n264), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT7), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT3), .B(G33), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n270), .B1(new_n271), .B2(G20), .ZN(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT3), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT3), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n249), .A2(KEYINPUT7), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n272), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n269), .B1(new_n281), .B2(G68), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n262), .B1(new_n282), .B2(KEYINPUT16), .ZN(new_n283));
  INV_X1    g0083(.A(new_n268), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n284), .A2(new_n266), .B1(G20), .B2(new_n263), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n275), .A2(G33), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n273), .A2(KEYINPUT3), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n249), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT82), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n289), .B1(new_n275), .B2(G33), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n273), .A2(KEYINPUT82), .A3(KEYINPUT3), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(new_n276), .A3(new_n291), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n270), .A2(new_n288), .B1(new_n292), .B2(new_n279), .ZN(new_n293));
  INV_X1    g0093(.A(G68), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n285), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT16), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n261), .B1(new_n283), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G169), .ZN(new_n299));
  OR2_X1    g0099(.A1(G223), .A2(G1698), .ZN(new_n300));
  INV_X1    g0100(.A(G226), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G1698), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n274), .A2(new_n300), .A3(new_n276), .A4(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(G33), .A2(G87), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n255), .B1(G33), .B2(G41), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G41), .ZN(new_n308));
  INV_X1    g0108(.A(G45), .ZN(new_n309));
  AOI21_X1  g0109(.A(G1), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(G33), .A2(G41), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n311), .A2(G1), .A3(G13), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n310), .A2(new_n312), .A3(G274), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n245), .B1(G41), .B2(G45), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n312), .A2(G232), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n299), .B1(new_n307), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n312), .B1(new_n303), .B2(new_n304), .ZN(new_n319));
  INV_X1    g0119(.A(G179), .ZN(new_n320));
  NOR3_X1   g0120(.A1(new_n319), .A2(new_n316), .A3(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(KEYINPUT83), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n307), .A2(new_n317), .A3(G179), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT83), .ZN(new_n324));
  OAI21_X1  g0124(.A(G169), .B1(new_n319), .B2(new_n316), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(KEYINPUT18), .B1(new_n298), .B2(new_n327), .ZN(new_n328));
  AND3_X1   g0128(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n324), .B1(new_n323), .B2(new_n325), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(KEYINPUT7), .B1(new_n277), .B2(new_n249), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n271), .A2(new_n278), .ZN(new_n333));
  OAI21_X1  g0133(.A(G68), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n334), .A2(KEYINPUT16), .A3(new_n285), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n292), .A2(new_n279), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n272), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n269), .B1(new_n337), .B2(G68), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n335), .B(new_n256), .C1(new_n338), .C2(KEYINPUT16), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n260), .A2(new_n244), .ZN(new_n340));
  INV_X1    g0140(.A(new_n248), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT18), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n331), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n328), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G200), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n347), .B1(new_n307), .B2(new_n317), .ZN(new_n348));
  INV_X1    g0148(.A(G190), .ZN(new_n349));
  NOR3_X1   g0149(.A1(new_n319), .A2(new_n316), .A3(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n339), .A2(new_n351), .A3(new_n342), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT17), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n339), .A2(new_n342), .A3(new_n351), .A4(KEYINPUT17), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n346), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n247), .A2(new_n294), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n358), .B(KEYINPUT12), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n265), .A2(G50), .B1(G20), .B2(new_n294), .ZN(new_n360));
  INV_X1    g0160(.A(G77), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n249), .A2(G33), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n363), .A2(KEYINPUT11), .A3(new_n256), .ZN(new_n364));
  AND3_X1   g0164(.A1(new_n246), .A2(new_n255), .A3(new_n254), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n365), .A2(G68), .A3(new_n253), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n359), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(KEYINPUT11), .B1(new_n363), .B2(new_n256), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n310), .A2(new_n312), .A3(KEYINPUT79), .A4(G274), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n312), .A2(G238), .A3(new_n314), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G274), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n374), .B1(new_n209), .B2(new_n311), .ZN(new_n375));
  AOI21_X1  g0175(.A(KEYINPUT79), .B1(new_n375), .B2(new_n310), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G1698), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n301), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G232), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(G1698), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n274), .A2(new_n379), .A3(new_n276), .A4(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G33), .A2(G97), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT78), .B1(new_n384), .B2(new_n306), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT78), .ZN(new_n386));
  AOI211_X1 g0186(.A(new_n386), .B(new_n312), .C1(new_n382), .C2(new_n383), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n377), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT13), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT13), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n377), .B(new_n390), .C1(new_n385), .C2(new_n387), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n389), .A2(G179), .A3(new_n391), .ZN(new_n392));
  OR2_X1    g0192(.A1(new_n299), .A2(KEYINPUT80), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(new_n389), .B2(new_n391), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT14), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n392), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AOI211_X1 g0196(.A(KEYINPUT14), .B(new_n393), .C1(new_n389), .C2(new_n391), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n370), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n389), .A2(new_n391), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n369), .B1(new_n399), .B2(new_n349), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n347), .B1(new_n389), .B2(new_n391), .ZN(new_n401));
  OR2_X1    g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n357), .A2(new_n398), .A3(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n277), .A2(new_n378), .ZN(new_n404));
  INV_X1    g0204(.A(new_n213), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n404), .A2(G223), .B1(new_n405), .B2(new_n277), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT69), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n378), .A2(G222), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n407), .B1(new_n277), .B2(new_n408), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n271), .A2(KEYINPUT69), .A3(G222), .A4(new_n378), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n312), .B1(new_n406), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n313), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n306), .A2(new_n310), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n414), .B1(G226), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n413), .A2(new_n320), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(G150), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n249), .A2(new_n273), .ZN(new_n419));
  OAI22_X1  g0219(.A1(new_n243), .A2(new_n362), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(G58), .A2(G68), .ZN(new_n421));
  INV_X1    g0221(.A(G50), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n249), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n256), .B1(new_n420), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT70), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n424), .A2(new_n425), .B1(new_n422), .B2(new_n247), .ZN(new_n426));
  OAI211_X1 g0226(.A(G50), .B(new_n253), .C1(new_n258), .C2(new_n259), .ZN(new_n427));
  OAI211_X1 g0227(.A(KEYINPUT70), .B(new_n256), .C1(new_n420), .C2(new_n423), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n416), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n299), .B1(new_n412), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n417), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(G200), .B1(new_n412), .B2(new_n430), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT76), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT10), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT75), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT9), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n429), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n439), .B1(new_n429), .B2(new_n440), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n413), .A2(G190), .A3(new_n416), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n426), .A2(KEYINPUT9), .A3(new_n427), .A4(new_n428), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n444), .A2(new_n434), .A3(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n438), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n442), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n429), .A2(new_n439), .A3(new_n440), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n446), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n450), .A2(new_n437), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n433), .B1(new_n447), .B2(new_n452), .ZN(new_n453));
  XNOR2_X1  g0253(.A(KEYINPUT15), .B(G87), .ZN(new_n454));
  OAI22_X1  g0254(.A1(new_n213), .A2(new_n249), .B1(new_n454), .B2(new_n362), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n243), .A2(new_n419), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n256), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n361), .B1(new_n250), .B2(new_n252), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n365), .A2(new_n458), .B1(new_n213), .B2(new_n247), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT73), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n457), .A2(new_n459), .A3(KEYINPUT73), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n414), .B1(G244), .B2(new_n415), .ZN(new_n465));
  NOR2_X1   g0265(.A1(G232), .A2(G1698), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n378), .A2(G238), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n271), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n468), .B(new_n306), .C1(G107), .C2(new_n271), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n299), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n464), .A2(KEYINPUT74), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n470), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n320), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(KEYINPUT74), .B1(new_n464), .B2(new_n471), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n464), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n470), .A2(new_n349), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n479), .B1(G200), .B2(new_n470), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n477), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n453), .A2(KEYINPUT77), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(KEYINPUT77), .B1(new_n453), .B2(new_n481), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n403), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n245), .A2(G45), .ZN(new_n485));
  NOR2_X1   g0285(.A1(KEYINPUT5), .A2(G41), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(KEYINPUT5), .A2(G41), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n485), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n375), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n214), .A2(G1698), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n491), .A2(new_n274), .A3(new_n276), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G33), .A2(G283), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n274), .A2(new_n276), .A3(G250), .A4(G1698), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n491), .A2(new_n274), .A3(new_n276), .A4(KEYINPUT4), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n494), .A2(new_n495), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n306), .ZN(new_n499));
  INV_X1    g0299(.A(G257), .ZN(new_n500));
  NOR3_X1   g0300(.A1(new_n489), .A2(new_n500), .A3(new_n306), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT86), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n349), .B1(new_n503), .B2(new_n347), .ZN(new_n504));
  AND4_X1   g0304(.A1(new_n490), .A2(new_n499), .A3(new_n502), .A4(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n503), .A2(G200), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n501), .B1(new_n498), .B2(new_n306), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n506), .B1(new_n507), .B2(new_n490), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n246), .A2(G97), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n245), .A2(G33), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n246), .A2(new_n511), .A3(new_n255), .A4(new_n254), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n510), .B1(new_n513), .B2(G97), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT85), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n419), .A2(new_n361), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT6), .ZN(new_n517));
  INV_X1    g0317(.A(G97), .ZN(new_n518));
  INV_X1    g0318(.A(G107), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(G97), .A2(G107), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n517), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n519), .A2(KEYINPUT6), .A3(G97), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n516), .B1(new_n524), .B2(G20), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n519), .B1(new_n336), .B2(new_n272), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT84), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR3_X1   g0328(.A1(new_n293), .A2(KEYINPUT84), .A3(new_n519), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n515), .B(new_n256), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(KEYINPUT84), .B1(new_n293), .B2(new_n519), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n337), .A2(new_n527), .A3(G107), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n532), .A2(new_n533), .A3(new_n525), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n515), .B1(new_n534), .B2(new_n256), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n509), .B(new_n514), .C1(new_n531), .C2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n514), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n256), .B1(new_n528), .B2(new_n529), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT85), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n537), .B1(new_n539), .B2(new_n530), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n507), .A2(new_n490), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n541), .A2(new_n320), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n299), .B1(new_n507), .B2(new_n490), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n536), .B1(new_n540), .B2(new_n544), .ZN(new_n545));
  OR2_X1    g0345(.A1(G238), .A2(G1698), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n214), .A2(G1698), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n274), .A2(new_n546), .A3(new_n276), .A4(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(G116), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n273), .A2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n312), .B1(new_n548), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n309), .A2(G1), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n312), .A2(G274), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(G250), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n555), .B1(new_n245), .B2(G45), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n312), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(G169), .B1(new_n552), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n375), .A2(new_n553), .B1(new_n312), .B2(new_n556), .ZN(new_n560));
  NOR2_X1   g0360(.A1(G238), .A2(G1698), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n561), .B1(new_n214), .B2(G1698), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n550), .B1(new_n562), .B2(new_n271), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n560), .B(G179), .C1(new_n563), .C2(new_n312), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT19), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n249), .B1(new_n383), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(G87), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n521), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n274), .A2(new_n276), .A3(new_n249), .A4(G68), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n566), .B1(new_n362), .B2(new_n518), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n256), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n454), .A2(new_n247), .ZN(new_n575));
  OR2_X1    g0375(.A1(new_n512), .A2(new_n454), .ZN(new_n576));
  AND4_X1   g0376(.A1(KEYINPUT87), .A2(new_n574), .A3(new_n575), .A4(new_n576), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n573), .A2(new_n256), .B1(new_n247), .B2(new_n454), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT87), .B1(new_n578), .B2(new_n576), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n565), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(G200), .B1(new_n552), .B2(new_n558), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT88), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n365), .A2(new_n582), .A3(G87), .A4(new_n511), .ZN(new_n583));
  OAI21_X1  g0383(.A(KEYINPUT88), .B1(new_n512), .B2(new_n568), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n581), .A2(new_n578), .A3(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n560), .B1(new_n563), .B2(new_n312), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n587), .A2(new_n349), .ZN(new_n588));
  OR2_X1    g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n580), .A2(new_n589), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n254), .A2(new_n255), .B1(G20), .B2(new_n549), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n495), .B(new_n249), .C1(G33), .C2(new_n518), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT20), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n591), .A2(KEYINPUT20), .A3(new_n592), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n247), .A2(new_n549), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n513), .A2(G116), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n488), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n553), .B1(new_n601), .B2(new_n486), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n602), .A2(G270), .A3(new_n312), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n378), .A2(G264), .ZN(new_n604));
  NOR2_X1   g0404(.A1(G257), .A2(G1698), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n606), .A2(new_n277), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n306), .B1(new_n271), .B2(G303), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n490), .B(new_n603), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n600), .A2(KEYINPUT21), .A3(G169), .A4(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT21), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n609), .A2(G169), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n598), .B1(new_n512), .B2(new_n549), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n613), .B1(new_n596), .B2(new_n595), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n611), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n609), .A2(new_n320), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n600), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n609), .A2(G200), .ZN(new_n618));
  INV_X1    g0418(.A(G303), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n312), .B1(new_n277), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(new_n277), .B2(new_n606), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n621), .A2(G190), .A3(new_n490), .A4(new_n603), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n618), .A2(new_n622), .A3(new_n614), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n610), .A2(new_n615), .A3(new_n617), .A4(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n590), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n274), .A2(new_n276), .A3(new_n249), .A4(G87), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(KEYINPUT22), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT22), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n271), .A2(new_n628), .A3(new_n249), .A4(G87), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT24), .ZN(new_n631));
  NAND2_X1  g0431(.A1(KEYINPUT23), .A2(G107), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n249), .A2(KEYINPUT23), .A3(G107), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n632), .B1(new_n633), .B2(KEYINPUT89), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT23), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n635), .A2(new_n519), .A3(G20), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT89), .ZN(new_n637));
  AOI21_X1  g0437(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n638));
  OAI22_X1  g0438(.A1(new_n636), .A2(new_n637), .B1(new_n638), .B2(G20), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n634), .A2(new_n639), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n630), .A2(new_n631), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n631), .B1(new_n630), .B2(new_n640), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n256), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT90), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OAI211_X1 g0445(.A(KEYINPUT90), .B(new_n256), .C1(new_n641), .C2(new_n642), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g0447(.A(KEYINPUT91), .B(KEYINPUT92), .Z(new_n648));
  OAI211_X1 g0448(.A(new_n519), .B(new_n247), .C1(new_n648), .C2(KEYINPUT25), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(KEYINPUT25), .ZN(new_n650));
  XNOR2_X1  g0450(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n513), .A2(G107), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n602), .A2(G264), .A3(new_n312), .ZN(new_n655));
  NOR2_X1   g0455(.A1(G250), .A2(G1698), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n656), .B1(new_n500), .B2(G1698), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n657), .A2(new_n271), .B1(G33), .B2(G294), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n490), .B(new_n655), .C1(new_n658), .C2(new_n312), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n659), .A2(new_n347), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(G190), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n647), .A2(new_n654), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n653), .B1(new_n645), .B2(new_n646), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n659), .A2(new_n299), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(G179), .B2(new_n659), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n625), .B(new_n664), .C1(new_n665), .C2(new_n667), .ZN(new_n668));
  NOR3_X1   g0468(.A1(new_n484), .A2(new_n545), .A3(new_n668), .ZN(G372));
  NAND2_X1  g0469(.A1(new_n402), .A2(new_n477), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n356), .B1(new_n670), .B2(new_n398), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT96), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n343), .B1(new_n318), .B2(new_n321), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(KEYINPUT18), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n343), .B(new_n344), .C1(new_n318), .C2(new_n321), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OR3_X1    g0476(.A1(new_n671), .A2(new_n672), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n447), .A2(new_n452), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n672), .B1(new_n671), .B2(new_n676), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n432), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n514), .B1(new_n531), .B2(new_n535), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n578), .A2(new_n576), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT87), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n578), .A2(KEYINPUT87), .A3(new_n576), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n559), .A2(new_n564), .A3(KEYINPUT93), .ZN(new_n689));
  AOI21_X1  g0489(.A(KEYINPUT93), .B1(new_n559), .B2(new_n564), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT94), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n588), .B1(new_n586), .B2(new_n692), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n581), .A2(new_n578), .A3(KEYINPUT94), .A4(new_n585), .ZN(new_n694));
  AOI22_X1  g0494(.A1(new_n688), .A2(new_n691), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n544), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n683), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT26), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(KEYINPUT95), .A3(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n540), .A2(new_n544), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n586), .A2(new_n588), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n701), .B1(new_n688), .B2(new_n565), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n700), .A2(KEYINPUT26), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(KEYINPUT95), .B1(new_n697), .B2(new_n698), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT93), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n565), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n559), .A2(new_n564), .A3(KEYINPUT93), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n708), .B(new_n709), .C1(new_n579), .C2(new_n577), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n683), .A2(new_n696), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n711), .A2(new_n536), .A3(new_n664), .A4(new_n695), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n610), .A2(new_n615), .A3(new_n617), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n665), .B2(new_n667), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n710), .B1(new_n712), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n706), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n682), .B1(new_n484), .B2(new_n718), .ZN(G369));
  NAND3_X1  g0519(.A1(new_n245), .A2(new_n249), .A3(G13), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n720), .A2(KEYINPUT27), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(KEYINPUT27), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n721), .A2(G213), .A3(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(G343), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(new_n614), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n713), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n728), .B1(new_n624), .B2(new_n727), .ZN(new_n729));
  XOR2_X1   g0529(.A(new_n729), .B(KEYINPUT97), .Z(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(G330), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n665), .A2(new_n667), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n664), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n665), .A2(new_n726), .ZN(new_n736));
  OAI22_X1  g0536(.A1(new_n735), .A2(new_n736), .B1(new_n734), .B2(new_n726), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n732), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n713), .A2(new_n726), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n734), .A2(new_n664), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n733), .A2(new_n726), .ZN(new_n742));
  AND2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n738), .A2(new_n743), .ZN(G399));
  NOR2_X1   g0544(.A1(new_n569), .A2(G116), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n204), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G41), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n746), .A2(new_n748), .A3(new_n245), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n749), .B1(new_n208), .B2(new_n748), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT98), .ZN(new_n751));
  XOR2_X1   g0551(.A(new_n751), .B(KEYINPUT28), .Z(new_n752));
  INV_X1    g0552(.A(KEYINPUT29), .ZN(new_n753));
  OAI211_X1 g0553(.A(new_n753), .B(new_n726), .C1(new_n706), .C2(new_n717), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n683), .A2(new_n695), .A3(new_n696), .A4(KEYINPUT26), .ZN(new_n756));
  NOR3_X1   g0556(.A1(new_n540), .A2(new_n544), .A3(new_n590), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n756), .B1(new_n757), .B2(KEYINPUT26), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT101), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n715), .A2(new_n759), .ZN(new_n760));
  OAI211_X1 g0560(.A(KEYINPUT101), .B(new_n714), .C1(new_n665), .C2(new_n667), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI211_X1 g0562(.A(new_n710), .B(new_n758), .C1(new_n762), .C2(new_n712), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n753), .B1(new_n763), .B2(new_n726), .ZN(new_n764));
  INV_X1    g0564(.A(G330), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n653), .B(new_n662), .C1(new_n645), .C2(new_n646), .ZN(new_n766));
  AND4_X1   g0566(.A1(new_n615), .A2(new_n610), .A3(new_n623), .A4(new_n617), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(new_n702), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n733), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n545), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n769), .A2(new_n770), .A3(new_n726), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT99), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(new_n552), .B2(new_n558), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n560), .B(KEYINPUT99), .C1(new_n563), .C2(new_n312), .ZN(new_n774));
  AND3_X1   g0574(.A1(new_n773), .A2(new_n774), .A3(new_n609), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n659), .A2(new_n320), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n775), .A2(new_n541), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(KEYINPUT100), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT100), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n775), .A2(new_n541), .A3(new_n776), .A4(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n659), .A2(new_n587), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n781), .A2(new_n616), .A3(new_n507), .ZN(new_n782));
  INV_X1    g0582(.A(KEYINPUT30), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n781), .A2(new_n616), .A3(KEYINPUT30), .A4(new_n507), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n778), .A2(new_n780), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(KEYINPUT31), .B1(new_n786), .B2(new_n725), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n784), .A2(new_n777), .A3(new_n785), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT31), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n726), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n787), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n765), .B1(new_n771), .B2(new_n791), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n755), .A2(new_n764), .A3(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n752), .B1(new_n793), .B2(G1), .ZN(G364));
  AND2_X1   g0594(.A1(new_n249), .A2(G13), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G45), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT102), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n797), .A2(new_n245), .A3(new_n748), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n271), .A2(G355), .A3(new_n204), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n241), .A2(new_n309), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n747), .A2(new_n271), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(G45), .B2(new_n207), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n800), .B1(G116), .B2(new_n204), .C1(new_n801), .C2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(G13), .A2(G33), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(G20), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n255), .B1(G20), .B2(new_n299), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n799), .B1(new_n804), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n808), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n349), .A2(new_n347), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n249), .A2(G179), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n277), .B1(new_n814), .B2(new_n619), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n249), .A2(new_n320), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NOR3_X1   g0617(.A1(new_n817), .A2(new_n347), .A3(G190), .ZN(new_n818));
  XNOR2_X1  g0618(.A(KEYINPUT33), .B(G317), .ZN(new_n819));
  NOR2_X1   g0619(.A1(G190), .A2(G200), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n813), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n818), .A2(new_n819), .B1(G329), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(G311), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n816), .A2(new_n820), .ZN(new_n825));
  INV_X1    g0625(.A(G322), .ZN(new_n826));
  NOR3_X1   g0626(.A1(new_n817), .A2(new_n349), .A3(G200), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n823), .B1(new_n824), .B2(new_n825), .C1(new_n826), .C2(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n813), .A2(new_n349), .A3(G200), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  OR2_X1    g0631(.A1(new_n831), .A2(KEYINPUT103), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(KEYINPUT103), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n815), .B(new_n829), .C1(G283), .C2(new_n835), .ZN(new_n836));
  NOR3_X1   g0636(.A1(new_n349), .A2(G179), .A3(G200), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n837), .A2(new_n249), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n812), .A2(new_n816), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n839), .A2(G294), .B1(new_n841), .B2(G326), .ZN(new_n842));
  XOR2_X1   g0642(.A(new_n842), .B(KEYINPUT104), .Z(new_n843));
  NOR2_X1   g0643(.A1(new_n838), .A2(new_n518), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n822), .A2(G159), .ZN(new_n845));
  INV_X1    g0645(.A(G58), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n271), .B1(new_n845), .B2(KEYINPUT32), .C1(new_n828), .C2(new_n846), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n844), .B(new_n847), .C1(KEYINPUT32), .C2(new_n845), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n834), .A2(new_n519), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n840), .A2(new_n422), .B1(new_n825), .B2(new_n213), .ZN(new_n850));
  INV_X1    g0650(.A(new_n818), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n851), .A2(new_n294), .B1(new_n814), .B2(new_n568), .ZN(new_n852));
  NOR3_X1   g0652(.A1(new_n849), .A2(new_n850), .A3(new_n852), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n836), .A2(new_n843), .B1(new_n848), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n807), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n810), .B1(new_n811), .B2(new_n854), .C1(new_n730), .C2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n731), .A2(new_n799), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n730), .A2(G330), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(G396));
  NOR2_X1   g0659(.A1(new_n718), .A2(new_n725), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n480), .A2(new_n478), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n464), .A2(new_n725), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n861), .B(new_n862), .C1(new_n475), .C2(new_n476), .ZN(new_n863));
  INV_X1    g0663(.A(new_n476), .ZN(new_n864));
  INV_X1    g0664(.A(new_n862), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n864), .A2(new_n474), .A3(new_n865), .A4(new_n472), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  OR3_X1    g0667(.A1(new_n860), .A2(KEYINPUT108), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(KEYINPUT108), .B1(new_n860), .B2(new_n867), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n481), .A2(new_n726), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n706), .B2(new_n717), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n771), .A2(new_n791), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(G330), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n798), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n870), .A2(new_n792), .A3(new_n873), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n811), .A2(new_n806), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n798), .B1(G77), .B2(new_n880), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n818), .A2(KEYINPUT105), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n818), .A2(KEYINPUT105), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(G283), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n814), .A2(new_n519), .ZN(new_n887));
  OAI22_X1  g0687(.A1(new_n840), .A2(new_n619), .B1(new_n825), .B2(new_n549), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n887), .B(new_n888), .C1(G294), .C2(new_n827), .ZN(new_n889));
  AOI211_X1 g0689(.A(new_n271), .B(new_n844), .C1(G311), .C2(new_n822), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n835), .A2(G87), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n886), .A2(new_n889), .A3(new_n890), .A4(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(G137), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n840), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(G159), .ZN(new_n895));
  OAI22_X1  g0695(.A1(new_n851), .A2(new_n418), .B1(new_n825), .B2(new_n895), .ZN(new_n896));
  AOI211_X1 g0696(.A(new_n894), .B(new_n896), .C1(G143), .C2(new_n827), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(KEYINPUT34), .ZN(new_n898));
  INV_X1    g0698(.A(G132), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n271), .B1(new_n821), .B2(new_n899), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT106), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n835), .A2(G68), .ZN(new_n903));
  INV_X1    g0703(.A(new_n814), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n839), .A2(G58), .B1(new_n904), .B2(G50), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n903), .B(new_n905), .C1(new_n897), .C2(KEYINPUT34), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n892), .B1(new_n902), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n881), .B1(new_n907), .B2(new_n808), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n867), .B2(new_n806), .ZN(new_n909));
  XOR2_X1   g0709(.A(new_n909), .B(KEYINPUT107), .Z(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n879), .A2(new_n911), .ZN(G384));
  NOR3_X1   g0712(.A1(new_n255), .A2(new_n249), .A3(new_n549), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n524), .B(KEYINPUT109), .Z(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT35), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n913), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n917), .B1(new_n916), .B2(new_n915), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n918), .B(KEYINPUT36), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n405), .B(new_n208), .C1(new_n846), .C2(new_n294), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n422), .A2(G68), .ZN(new_n921));
  AOI211_X1 g0721(.A(new_n245), .B(G13), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n764), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n484), .B1(new_n924), .B2(new_n754), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n925), .A2(new_n681), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n294), .B1(new_n272), .B2(new_n280), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n296), .B1(new_n927), .B2(new_n269), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n928), .A2(new_n335), .A3(new_n256), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n723), .B1(new_n929), .B2(new_n342), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n346), .B2(new_n356), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n331), .A2(new_n343), .ZN(new_n932));
  INV_X1    g0732(.A(new_n723), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n343), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT37), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n932), .A2(new_n934), .A3(new_n935), .A4(new_n352), .ZN(new_n936));
  AND3_X1   g0736(.A1(new_n339), .A2(new_n342), .A3(new_n351), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n929), .A2(new_n342), .B1(new_n325), .B2(new_n323), .ZN(new_n938));
  NOR3_X1   g0738(.A1(new_n937), .A2(new_n938), .A3(new_n930), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n936), .B1(new_n939), .B2(new_n935), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n931), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT38), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n931), .A2(new_n940), .A3(KEYINPUT38), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n370), .A2(new_n725), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n398), .A2(new_n402), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n946), .B1(new_n398), .B2(new_n402), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT95), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n586), .A2(new_n692), .ZN(new_n952));
  INV_X1    g0752(.A(new_n588), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n952), .A2(new_n953), .A3(new_n694), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n710), .A2(new_n954), .ZN(new_n955));
  NOR3_X1   g0755(.A1(new_n540), .A2(new_n955), .A3(new_n544), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n951), .B1(new_n956), .B2(KEYINPUT26), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n957), .A2(new_n703), .A3(new_n699), .ZN(new_n958));
  INV_X1    g0758(.A(new_n710), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n664), .A2(new_n695), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n545), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n959), .B1(new_n961), .B2(new_n715), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n871), .B1(new_n958), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n477), .A2(new_n726), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n945), .B(new_n950), .C1(new_n963), .C2(new_n965), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n394), .A2(new_n395), .ZN(new_n967));
  INV_X1    g0767(.A(new_n397), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n967), .A2(new_n968), .A3(new_n392), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n969), .A2(new_n370), .A3(new_n726), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n943), .A2(KEYINPUT39), .A3(new_n944), .ZN(new_n972));
  AND3_X1   g0772(.A1(new_n931), .A2(new_n940), .A3(KEYINPUT38), .ZN(new_n973));
  INV_X1    g0773(.A(new_n934), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n354), .A2(KEYINPUT110), .A3(new_n355), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n975), .A2(new_n674), .A3(new_n675), .ZN(new_n976));
  AOI21_X1  g0776(.A(KEYINPUT110), .B1(new_n354), .B2(new_n355), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n974), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n673), .A2(new_n934), .A3(new_n352), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(KEYINPUT37), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n936), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n973), .B1(new_n982), .B2(new_n942), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n971), .B(new_n972), .C1(new_n983), .C2(KEYINPUT39), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n676), .A2(new_n723), .ZN(new_n985));
  AND3_X1   g0785(.A1(new_n966), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n926), .B(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n786), .A2(KEYINPUT31), .A3(new_n725), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n989), .A2(new_n787), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n771), .A2(new_n990), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n863), .A2(new_n866), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n400), .A2(new_n401), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n370), .B(new_n725), .C1(new_n969), .C2(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n398), .A2(new_n402), .A3(new_n946), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n992), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(KEYINPUT38), .B1(new_n978), .B2(new_n981), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n991), .B(new_n996), .C1(new_n997), .C2(new_n973), .ZN(new_n998));
  NOR3_X1   g0798(.A1(new_n668), .A2(new_n545), .A3(new_n725), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n786), .A2(new_n725), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n789), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n988), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n867), .B1(new_n947), .B2(new_n948), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(KEYINPUT40), .B1(new_n943), .B2(new_n944), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n998), .A2(KEYINPUT40), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n484), .B2(new_n1003), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n484), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT40), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT110), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n356), .A2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1012), .A2(new_n674), .A3(new_n675), .A4(new_n975), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n1013), .A2(new_n974), .B1(new_n936), .B2(new_n980), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n944), .B1(new_n1014), .B2(KEYINPUT38), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1010), .B1(new_n1005), .B2(new_n1015), .ZN(new_n1016));
  AND3_X1   g0816(.A1(new_n1006), .A2(new_n991), .A3(new_n996), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1009), .B(new_n991), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1008), .A2(new_n1018), .A3(G330), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n987), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n245), .B2(new_n795), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n987), .A2(new_n1019), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n923), .B1(new_n1021), .B2(new_n1022), .ZN(G367));
  NAND2_X1  g0823(.A1(new_n700), .A2(new_n725), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT111), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT112), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n770), .B1(new_n540), .B2(new_n726), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1026), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n733), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n725), .B1(new_n1031), .B2(new_n711), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n741), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT42), .Z(new_n1034));
  NOR2_X1   g0834(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT43), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n726), .B1(new_n578), .B2(new_n585), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n955), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n959), .A2(new_n1037), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1035), .A2(new_n1036), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(new_n1036), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1040), .A2(KEYINPUT43), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1043), .B(new_n1044), .C1(new_n1032), .C2(new_n1034), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1042), .A2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1047), .A2(new_n738), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1042), .A2(new_n1048), .A3(new_n1045), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n748), .B(KEYINPUT41), .Z(new_n1052));
  NAND2_X1  g0852(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1053), .A2(new_n743), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1054), .A2(KEYINPUT44), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT44), .ZN(new_n1056));
  NOR3_X1   g0856(.A1(new_n1053), .A2(new_n1056), .A3(new_n743), .ZN(new_n1057));
  AND3_X1   g0857(.A1(new_n1053), .A2(KEYINPUT45), .A3(new_n743), .ZN(new_n1058));
  AOI21_X1  g0858(.A(KEYINPUT45), .B1(new_n1053), .B2(new_n743), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n1055), .A2(new_n1057), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1060), .A2(new_n732), .A3(new_n737), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n741), .B1(new_n737), .B2(new_n740), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(new_n731), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n738), .B1(new_n1058), .B2(new_n1059), .C1(new_n1055), .C2(new_n1057), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1061), .A2(new_n793), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1052), .B1(new_n1066), .B2(new_n793), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n797), .A2(new_n245), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1050), .B(new_n1051), .C1(new_n1067), .C2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n802), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n233), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n809), .B1(new_n204), .B2(new_n454), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n798), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n825), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n827), .A2(G150), .B1(G50), .B2(new_n1075), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1076), .B1(new_n893), .B2(new_n821), .C1(new_n884), .C2(new_n895), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n213), .A2(new_n830), .B1(new_n814), .B2(new_n846), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n277), .B(new_n1078), .C1(G143), .C2(new_n841), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n839), .A2(G68), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n904), .A2(G116), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT46), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n271), .B1(new_n1075), .B2(G283), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1083), .B(new_n1084), .C1(new_n519), .C2(new_n838), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n831), .A2(G97), .B1(new_n822), .B2(G317), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n827), .A2(G303), .B1(new_n841), .B2(G311), .ZN(new_n1087));
  INV_X1    g0887(.A(G294), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1086), .B(new_n1087), .C1(new_n884), .C2(new_n1088), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n1077), .A2(new_n1081), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT47), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1074), .B1(new_n1091), .B2(new_n808), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n1040), .B2(new_n855), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1070), .A2(new_n1093), .ZN(G387));
  OR2_X1    g0894(.A1(new_n737), .A2(new_n855), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n271), .A2(new_n204), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n1096), .A2(new_n745), .B1(G107), .B2(new_n204), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n229), .A2(G45), .ZN(new_n1098));
  AOI211_X1 g0898(.A(G45), .B(new_n746), .C1(G68), .C2(G77), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n243), .A2(G50), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT50), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1071), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1097), .B1(new_n1098), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n809), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n798), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n814), .A2(new_n213), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n271), .B1(new_n821), .B2(new_n418), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n1106), .B(new_n1107), .C1(new_n835), .C2(G97), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT113), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n838), .A2(new_n454), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n422), .A2(new_n828), .B1(new_n851), .B2(new_n243), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n840), .A2(new_n895), .B1(new_n825), .B2(new_n294), .ZN(new_n1112));
  NOR4_X1   g0912(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .A4(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT114), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n827), .A2(G317), .B1(new_n841), .B2(G322), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1115), .B1(new_n619), .B2(new_n825), .C1(new_n884), .C2(new_n824), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT48), .ZN(new_n1117));
  OR2_X1    g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n839), .A2(G283), .B1(new_n904), .B2(G294), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT49), .ZN(new_n1122));
  OR2_X1    g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n830), .A2(new_n549), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n271), .B(new_n1125), .C1(G326), .C2(new_n822), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1123), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1114), .A2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1105), .B1(new_n1128), .B2(new_n808), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n1064), .A2(new_n1069), .B1(new_n1095), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1064), .A2(new_n793), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n748), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1064), .A2(new_n793), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1130), .B1(new_n1132), .B2(new_n1133), .ZN(G393));
  AND2_X1   g0934(.A1(new_n238), .A2(new_n802), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n809), .B1(new_n518), .B2(new_n204), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n798), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n849), .B1(new_n885), .B2(G303), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n827), .A2(G311), .B1(new_n841), .B2(G317), .ZN(new_n1139));
  XOR2_X1   g0939(.A(new_n1139), .B(KEYINPUT52), .Z(new_n1140));
  OAI21_X1  g0940(.A(new_n277), .B1(new_n821), .B2(new_n826), .ZN(new_n1141));
  INV_X1    g0941(.A(G283), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n1142), .A2(new_n814), .B1(new_n825), .B2(new_n1088), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n1141), .B(new_n1143), .C1(G116), .C2(new_n839), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1138), .A2(new_n1140), .A3(new_n1144), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n827), .A2(G159), .B1(new_n841), .B2(G150), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT51), .ZN(new_n1147));
  INV_X1    g0947(.A(G143), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n814), .A2(new_n294), .B1(new_n821), .B2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n838), .A2(new_n361), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n271), .B1(new_n825), .B2(new_n243), .ZN(new_n1151));
  NOR3_X1   g0951(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n891), .B(new_n1152), .C1(new_n422), .C2(new_n884), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1145), .B1(new_n1147), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1137), .B1(new_n1154), .B2(new_n808), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1047), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1155), .B1(new_n1156), .B2(new_n855), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1061), .A2(new_n1065), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1157), .B1(new_n1158), .B2(new_n1068), .ZN(new_n1159));
  AND2_X1   g0959(.A1(new_n1066), .A2(new_n748), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1158), .A2(new_n1131), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1159), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(G390));
  OAI21_X1  g0963(.A(new_n950), .B1(new_n963), .B2(new_n965), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n970), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT39), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1015), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(new_n972), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1165), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT115), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n970), .B(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1015), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n763), .A2(new_n726), .A3(new_n867), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1174), .A2(new_n964), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1173), .B1(new_n1175), .B2(new_n949), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n792), .A2(new_n996), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1169), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n991), .A2(G330), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1179), .A2(new_n1004), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n1164), .A2(new_n970), .B1(new_n1167), .B2(new_n972), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1174), .A2(new_n964), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1172), .B1(new_n1182), .B2(new_n950), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1180), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1178), .A2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1185), .A2(new_n1068), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1168), .A2(new_n805), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n798), .B1(new_n244), .B2(new_n880), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n885), .A2(G107), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n825), .A2(new_n518), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n840), .A2(new_n1142), .B1(new_n821), .B2(new_n1088), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n1190), .B(new_n1191), .C1(G116), .C2(new_n827), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n271), .B(new_n1150), .C1(G87), .C2(new_n904), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1189), .A2(new_n903), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n277), .B1(new_n831), .B2(G50), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n885), .A2(G137), .B1(KEYINPUT118), .B2(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n814), .A2(new_n418), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT53), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1196), .B(new_n1198), .C1(KEYINPUT118), .C2(new_n1195), .ZN(new_n1199));
  XOR2_X1   g0999(.A(KEYINPUT54), .B(G143), .Z(new_n1200));
  AOI22_X1  g1000(.A1(new_n827), .A2(G132), .B1(new_n1075), .B2(new_n1200), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n841), .A2(G128), .B1(new_n822), .B2(G125), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1201), .B(new_n1202), .C1(new_n895), .C2(new_n838), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1194), .B1(new_n1199), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1188), .B1(new_n1204), .B2(new_n808), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1186), .B1(new_n1187), .B2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n950), .B1(new_n792), .B2(new_n867), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n1180), .A2(new_n1207), .B1(new_n963), .B2(new_n965), .ZN(new_n1208));
  OAI211_X1 g1008(.A(G330), .B(new_n867), .C1(new_n999), .C2(new_n1002), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n949), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n1177), .ZN(new_n1211));
  NOR3_X1   g1011(.A1(new_n1211), .A2(new_n1182), .A3(KEYINPUT116), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT116), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n949), .A2(new_n1209), .B1(new_n792), .B2(new_n996), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1213), .B1(new_n1175), .B2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1208), .B1(new_n1212), .B2(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n484), .A2(new_n1179), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(new_n925), .A2(new_n681), .A3(new_n1217), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1216), .A2(new_n1178), .A3(new_n1184), .A4(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1219), .A2(KEYINPUT117), .A3(new_n748), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n1185), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1220), .A2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(KEYINPUT117), .B1(new_n1219), .B2(new_n748), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1206), .B1(new_n1223), .B2(new_n1224), .ZN(G378));
  OAI21_X1  g1025(.A(new_n949), .B1(new_n876), .B2(new_n992), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1003), .A2(new_n765), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n996), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n1226), .A2(new_n1228), .B1(new_n873), .B2(new_n964), .ZN(new_n1229));
  OAI21_X1  g1029(.A(KEYINPUT116), .B1(new_n1211), .B2(new_n1182), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1175), .A2(new_n1214), .A3(new_n1213), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1229), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1218), .B1(new_n1185), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n429), .A2(new_n933), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n453), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1234), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n433), .B(new_n1236), .C1(new_n447), .C2(new_n452), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(new_n1235), .A2(new_n1237), .A3(new_n1239), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(new_n443), .A2(new_n438), .A3(new_n446), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n437), .B1(new_n450), .B2(new_n451), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n432), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1236), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n453), .A2(new_n1234), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1238), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1240), .A2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n1007), .B2(new_n765), .ZN(new_n1248));
  OR2_X1    g1048(.A1(new_n1240), .A2(new_n1246), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1249), .B(G330), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1248), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n986), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1248), .A2(new_n1250), .A3(new_n986), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1233), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT57), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n1219), .A2(new_n1218), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(KEYINPUT57), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1258), .A2(new_n1260), .A3(new_n748), .ZN(new_n1261));
  AND3_X1   g1061(.A1(new_n1248), .A2(new_n1250), .A3(new_n986), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n986), .B1(new_n1248), .B2(new_n1250), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1069), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1247), .A2(new_n805), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n798), .B1(G50), .B2(new_n880), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n846), .A2(new_n830), .B1(new_n825), .B2(new_n454), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n277), .A2(new_n308), .ZN(new_n1268));
  NOR3_X1   g1068(.A1(new_n1267), .A2(new_n1106), .A3(new_n1268), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n827), .A2(G107), .B1(G283), .B2(new_n822), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n818), .A2(G97), .B1(new_n841), .B2(G116), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1269), .A2(new_n1080), .A3(new_n1270), .A4(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT58), .ZN(new_n1273));
  AOI21_X1  g1073(.A(G50), .B1(new_n273), .B2(new_n308), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n1272), .A2(new_n1273), .B1(new_n1268), .B2(new_n1274), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n827), .A2(G128), .B1(new_n841), .B2(G125), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n893), .B2(new_n825), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(new_n818), .A2(G132), .B1(new_n904), .B2(new_n1200), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1278), .B1(new_n418), .B2(new_n838), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1277), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1281), .A2(KEYINPUT59), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n273), .B(new_n308), .C1(new_n830), .C2(new_n895), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1283), .B1(G124), .B2(new_n822), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT59), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1284), .B1(new_n1280), .B2(new_n1285), .ZN(new_n1286));
  OAI221_X1 g1086(.A(new_n1275), .B1(new_n1273), .B2(new_n1272), .C1(new_n1282), .C2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1266), .B1(new_n1287), .B2(new_n808), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1265), .A2(new_n1288), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1264), .A2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1261), .A2(new_n1290), .ZN(G375));
  OR3_X1    g1091(.A1(new_n925), .A2(new_n681), .A3(new_n1217), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1232), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1052), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1293), .A2(new_n1221), .A3(new_n1294), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n1295), .B(KEYINPUT119), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n798), .B1(G68), .B2(new_n880), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n885), .A2(new_n1200), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n839), .A2(G50), .ZN(new_n1299));
  OAI22_X1  g1099(.A1(new_n840), .A2(new_n899), .B1(new_n814), .B2(new_n895), .ZN(new_n1300));
  AOI211_X1 g1100(.A(new_n277), .B(new_n1300), .C1(G58), .C2(new_n831), .ZN(new_n1301));
  INV_X1    g1101(.A(G128), .ZN(new_n1302));
  OAI22_X1  g1102(.A1(new_n825), .A2(new_n418), .B1(new_n821), .B2(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1303), .B1(G137), .B2(new_n827), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1298), .A2(new_n1299), .A3(new_n1301), .A4(new_n1304), .ZN(new_n1305));
  AOI211_X1 g1105(.A(new_n271), .B(new_n1110), .C1(G97), .C2(new_n904), .ZN(new_n1306));
  AOI22_X1  g1106(.A1(new_n827), .A2(G283), .B1(G107), .B2(new_n1075), .ZN(new_n1307));
  AOI22_X1  g1107(.A1(new_n841), .A2(G294), .B1(new_n822), .B2(G303), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1306), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  OAI22_X1  g1109(.A1(new_n884), .A2(new_n549), .B1(new_n834), .B2(new_n361), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1305), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1297), .B1(new_n1311), .B2(new_n808), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1312), .B1(new_n950), .B2(new_n806), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1313), .B1(new_n1232), .B2(new_n1068), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1296), .A2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(G381));
  NOR3_X1   g1116(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1317));
  XNOR2_X1  g1117(.A(new_n1317), .B(KEYINPUT120), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1070), .A2(new_n1093), .A3(new_n1162), .ZN(new_n1319));
  NOR3_X1   g1119(.A1(new_n1318), .A2(G381), .A3(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(G378), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1320), .A2(new_n1321), .A3(new_n1290), .A4(new_n1261), .ZN(new_n1322));
  XNOR2_X1  g1122(.A(new_n1322), .B(KEYINPUT121), .ZN(G407));
  NAND2_X1  g1123(.A1(new_n1321), .A2(new_n724), .ZN(new_n1324));
  OAI211_X1 g1124(.A(G407), .B(G213), .C1(G375), .C2(new_n1324), .ZN(G409));
  INV_X1    g1125(.A(KEYINPUT125), .ZN(new_n1326));
  XOR2_X1   g1126(.A(G393), .B(G396), .Z(new_n1327));
  INV_X1    g1127(.A(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1162), .B1(new_n1070), .B2(new_n1093), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1329), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1328), .B1(new_n1330), .B2(new_n1319), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1319), .ZN(new_n1332));
  NOR3_X1   g1132(.A1(new_n1332), .A2(new_n1327), .A3(new_n1329), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1326), .B1(new_n1331), .B2(new_n1333), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1327), .B1(new_n1332), .B2(new_n1329), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1330), .A2(new_n1319), .A3(new_n1328), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1335), .A2(new_n1336), .A3(KEYINPUT125), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1334), .A2(new_n1337), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1261), .A2(G378), .A3(new_n1290), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1264), .A2(new_n1289), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1340), .B1(new_n1294), .B2(new_n1259), .ZN(new_n1341));
  OAI21_X1  g1141(.A(KEYINPUT122), .B1(G378), .B2(new_n1341), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1290), .B1(new_n1256), .B2(new_n1052), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1224), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1344), .A2(new_n1222), .A3(new_n1220), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT122), .ZN(new_n1346));
  NAND4_X1  g1146(.A1(new_n1343), .A2(new_n1345), .A3(new_n1346), .A4(new_n1206), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1339), .A2(new_n1342), .A3(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n724), .A2(G213), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1232), .A2(new_n1292), .A3(KEYINPUT60), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1350), .A2(new_n748), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1221), .A2(KEYINPUT60), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1351), .B1(new_n1293), .B2(new_n1352), .ZN(new_n1353));
  OAI211_X1 g1153(.A(new_n879), .B(new_n911), .C1(new_n1353), .C2(new_n1314), .ZN(new_n1354));
  INV_X1    g1154(.A(new_n1314), .ZN(new_n1355));
  AND2_X1   g1155(.A1(new_n1352), .A2(new_n1293), .ZN(new_n1356));
  OAI211_X1 g1156(.A(G384), .B(new_n1355), .C1(new_n1356), .C2(new_n1351), .ZN(new_n1357));
  AND2_X1   g1157(.A1(new_n1354), .A2(new_n1357), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1348), .A2(new_n1349), .A3(new_n1358), .ZN(new_n1359));
  XOR2_X1   g1159(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n1360));
  NAND2_X1  g1160(.A1(new_n1359), .A2(new_n1360), .ZN(new_n1361));
  AND3_X1   g1161(.A1(new_n1354), .A2(new_n1357), .A3(KEYINPUT62), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1348), .A2(new_n1349), .A3(new_n1362), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1363), .A2(KEYINPUT124), .ZN(new_n1364));
  INV_X1    g1164(.A(KEYINPUT124), .ZN(new_n1365));
  NAND4_X1  g1165(.A1(new_n1348), .A2(new_n1365), .A3(new_n1349), .A4(new_n1362), .ZN(new_n1366));
  NAND3_X1  g1166(.A1(new_n1361), .A2(new_n1364), .A3(new_n1366), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1368));
  NAND3_X1  g1168(.A1(new_n724), .A2(G213), .A3(G2897), .ZN(new_n1369));
  AND3_X1   g1169(.A1(new_n1354), .A2(new_n1357), .A3(new_n1369), .ZN(new_n1370));
  AOI21_X1  g1170(.A(new_n1369), .B1(new_n1354), .B2(new_n1357), .ZN(new_n1371));
  NOR2_X1   g1171(.A1(new_n1370), .A2(new_n1371), .ZN(new_n1372));
  AOI21_X1  g1172(.A(KEYINPUT61), .B1(new_n1368), .B2(new_n1372), .ZN(new_n1373));
  AOI21_X1  g1173(.A(new_n1338), .B1(new_n1367), .B2(new_n1373), .ZN(new_n1374));
  INV_X1    g1174(.A(KEYINPUT63), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1359), .A2(new_n1375), .ZN(new_n1376));
  NOR2_X1   g1176(.A1(new_n1331), .A2(new_n1333), .ZN(new_n1377));
  NAND4_X1  g1177(.A1(new_n1348), .A2(KEYINPUT63), .A3(new_n1349), .A4(new_n1358), .ZN(new_n1378));
  NAND4_X1  g1178(.A1(new_n1373), .A2(new_n1376), .A3(new_n1377), .A4(new_n1378), .ZN(new_n1379));
  INV_X1    g1179(.A(new_n1379), .ZN(new_n1380));
  OAI21_X1  g1180(.A(KEYINPUT126), .B1(new_n1374), .B2(new_n1380), .ZN(new_n1381));
  INV_X1    g1181(.A(KEYINPUT126), .ZN(new_n1382));
  NAND2_X1  g1182(.A1(new_n1368), .A2(new_n1372), .ZN(new_n1383));
  INV_X1    g1183(.A(KEYINPUT61), .ZN(new_n1384));
  NAND2_X1  g1184(.A1(new_n1383), .A2(new_n1384), .ZN(new_n1385));
  AOI22_X1  g1185(.A1(KEYINPUT124), .A2(new_n1363), .B1(new_n1359), .B2(new_n1360), .ZN(new_n1386));
  AOI21_X1  g1186(.A(new_n1385), .B1(new_n1386), .B2(new_n1366), .ZN(new_n1387));
  OAI211_X1 g1187(.A(new_n1382), .B(new_n1379), .C1(new_n1387), .C2(new_n1338), .ZN(new_n1388));
  NAND2_X1  g1188(.A1(new_n1381), .A2(new_n1388), .ZN(G405));
  NAND2_X1  g1189(.A1(G375), .A2(new_n1321), .ZN(new_n1390));
  NAND2_X1  g1190(.A1(new_n1390), .A2(new_n1339), .ZN(new_n1391));
  INV_X1    g1191(.A(KEYINPUT127), .ZN(new_n1392));
  NAND2_X1  g1192(.A1(new_n1358), .A2(new_n1392), .ZN(new_n1393));
  XNOR2_X1  g1193(.A(new_n1391), .B(new_n1393), .ZN(new_n1394));
  XNOR2_X1  g1194(.A(new_n1338), .B(new_n1394), .ZN(G402));
endmodule


