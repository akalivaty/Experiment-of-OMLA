//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 1 1 1 0 1 1 0 0 0 0 1 1 1 1 1 1 1 0 1 1 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n561, new_n562, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1272, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT66), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT67), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT68), .Z(G217));
  NOR4_X1   g026(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n455), .A2(G567), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT69), .Z(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(G2106), .B2(new_n453), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  OR2_X1    g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n461), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n464), .A2(G137), .A3(new_n461), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n461), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n467), .A2(new_n471), .ZN(G160));
  INV_X1    g047(.A(KEYINPUT70), .ZN(new_n473));
  AND2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n473), .B1(new_n476), .B2(G2105), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n464), .A2(KEYINPUT70), .A3(new_n461), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n477), .A2(new_n478), .A3(G136), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n461), .A2(G112), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n479), .B(new_n481), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT71), .ZN(G162));
  OAI211_X1 g060(.A(G126), .B(G2105), .C1(new_n474), .C2(new_n475), .ZN(new_n486));
  INV_X1    g061(.A(G114), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n461), .A2(G138), .ZN(new_n491));
  OAI21_X1  g066(.A(KEYINPUT4), .B1(new_n476), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(new_n491), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n464), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n490), .B1(new_n492), .B2(new_n495), .ZN(G164));
  NOR2_X1   g071(.A1(KEYINPUT5), .A2(G543), .ZN(new_n497));
  AND2_X1   g072(.A1(KEYINPUT5), .A2(G543), .ZN(new_n498));
  AND2_X1   g073(.A1(KEYINPUT6), .A2(G651), .ZN(new_n499));
  NOR2_X1   g074(.A1(KEYINPUT6), .A2(G651), .ZN(new_n500));
  OAI22_X1  g075(.A1(new_n497), .A2(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G88), .ZN(new_n502));
  OAI21_X1  g077(.A(G543), .B1(new_n499), .B2(new_n500), .ZN(new_n503));
  INV_X1    g078(.A(G50), .ZN(new_n504));
  OAI22_X1  g079(.A1(new_n501), .A2(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  OAI21_X1  g081(.A(G62), .B1(new_n498), .B2(new_n497), .ZN(new_n507));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT72), .B1(new_n505), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n507), .A2(new_n508), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G651), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n514));
  OR2_X1    g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OR2_X1    g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n517), .A2(new_n520), .A3(G88), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n522), .B1(new_n518), .B2(new_n519), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G50), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n513), .A2(new_n514), .A3(new_n521), .A4(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n511), .A2(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  INV_X1    g103(.A(G51), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n503), .A2(new_n529), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n498), .A2(new_n497), .ZN(new_n534));
  OAI21_X1  g109(.A(G89), .B1(new_n499), .B2(new_n500), .ZN(new_n535));
  NAND2_X1  g110(.A1(G63), .A2(G651), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n533), .A2(new_n537), .ZN(G168));
  INV_X1    g113(.A(G64), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n539), .B1(new_n515), .B2(new_n516), .ZN(new_n540));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g117(.A(G651), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  OAI211_X1 g118(.A(G52), .B(G543), .C1(new_n499), .C2(new_n500), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n517), .A2(new_n520), .A3(G90), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  XNOR2_X1  g122(.A(KEYINPUT74), .B(G81), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(G43), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n501), .A2(new_n549), .B1(new_n503), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G56), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n534), .B2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT73), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n506), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  OAI211_X1 g131(.A(KEYINPUT73), .B(new_n552), .C1(new_n534), .C2(new_n553), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n551), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n534), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n515), .A2(new_n516), .B1(new_n518), .B2(new_n519), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n566), .A2(G651), .B1(new_n567), .B2(G91), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n523), .A2(G53), .ZN(new_n569));
  AND2_X1   g144(.A1(new_n569), .A2(KEYINPUT9), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n569), .A2(KEYINPUT9), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n568), .B1(new_n570), .B2(new_n571), .ZN(G299));
  INV_X1    g147(.A(G168), .ZN(G286));
  OAI21_X1  g148(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n523), .A2(G49), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n517), .A2(new_n520), .A3(G87), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n574), .A2(new_n575), .A3(new_n576), .A4(KEYINPUT75), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G288));
  INV_X1    g157(.A(G86), .ZN(new_n583));
  INV_X1    g158(.A(G48), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n501), .A2(new_n583), .B1(new_n503), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g160(.A(G61), .B1(new_n498), .B2(new_n497), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n506), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g163(.A(KEYINPUT76), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  NOR3_X1   g165(.A1(new_n585), .A2(KEYINPUT76), .A3(new_n588), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n590), .A2(new_n591), .ZN(G305));
  AOI22_X1  g167(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n593), .A2(new_n506), .ZN(new_n594));
  INV_X1    g169(.A(G85), .ZN(new_n595));
  INV_X1    g170(.A(G47), .ZN(new_n596));
  OAI22_X1  g171(.A1(new_n501), .A2(new_n595), .B1(new_n503), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n567), .A2(KEYINPUT10), .A3(G92), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n602));
  INV_X1    g177(.A(G92), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n501), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n601), .A2(new_n604), .B1(G54), .B2(new_n523), .ZN(new_n605));
  NAND2_X1  g180(.A1(G79), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G66), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n534), .B2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT77), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI211_X1 g185(.A(KEYINPUT77), .B(new_n606), .C1(new_n534), .C2(new_n607), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n610), .A2(G651), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n605), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n600), .B1(new_n614), .B2(G868), .ZN(G284));
  OAI21_X1  g190(.A(new_n600), .B1(new_n614), .B2(G868), .ZN(G321));
  NAND2_X1  g191(.A1(G286), .A2(G868), .ZN(new_n617));
  INV_X1    g192(.A(G299), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G868), .ZN(G297));
  OAI21_X1  g194(.A(new_n617), .B1(new_n618), .B2(G868), .ZN(G280));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n614), .B1(new_n621), .B2(G860), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT78), .ZN(G148));
  NAND2_X1  g198(.A1(new_n614), .A2(new_n621), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G868), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n625), .A2(KEYINPUT79), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(KEYINPUT79), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n626), .B(new_n627), .C1(G868), .C2(new_n558), .ZN(G323));
  XNOR2_X1  g203(.A(KEYINPUT80), .B(KEYINPUT11), .ZN(new_n629));
  XNOR2_X1  g204(.A(G323), .B(new_n629), .ZN(G282));
  OR2_X1    g205(.A1(new_n461), .A2(G111), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n631), .A2(KEYINPUT81), .ZN(new_n632));
  OAI21_X1  g207(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n633), .B1(new_n631), .B2(KEYINPUT81), .ZN(new_n634));
  AOI22_X1  g209(.A1(new_n632), .A2(new_n634), .B1(new_n480), .B2(G123), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n477), .A2(new_n478), .A3(G135), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n637), .A2(G2096), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n464), .A2(new_n469), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT12), .Z(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT13), .Z(new_n641));
  INV_X1    g216(.A(G2100), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n638), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n637), .A2(G2096), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n643), .B(new_n644), .C1(new_n642), .C2(new_n641), .ZN(G156));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT84), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2427), .B(G2430), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  XOR2_X1   g226(.A(KEYINPUT83), .B(KEYINPUT14), .Z(new_n652));
  NAND3_X1  g227(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g233(.A1(new_n650), .A2(new_n651), .A3(new_n652), .A4(new_n656), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2451), .B(G2454), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n661), .B(new_n662), .Z(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n658), .A2(new_n663), .A3(new_n659), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n665), .A2(G14), .A3(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(G401));
  XOR2_X1   g243(.A(G2072), .B(G2078), .Z(new_n669));
  XNOR2_X1  g244(.A(G2084), .B(G2090), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT85), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n669), .B1(new_n674), .B2(KEYINPUT18), .ZN(new_n675));
  INV_X1    g250(.A(G2096), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n675), .A2(new_n676), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n672), .A2(new_n673), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n680), .A2(KEYINPUT17), .A3(new_n674), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT18), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n681), .A2(new_n682), .A3(new_n642), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n642), .B1(new_n681), .B2(new_n682), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n679), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n681), .A2(new_n682), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(G2100), .ZN(new_n688));
  NAND4_X1  g263(.A1(new_n688), .A2(new_n677), .A3(new_n678), .A4(new_n683), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(G227));
  XNOR2_X1  g266(.A(G1981), .B(G1986), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT86), .B(KEYINPUT19), .Z(new_n694));
  XNOR2_X1  g269(.A(G1971), .B(G1976), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1956), .B(G2474), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1961), .B(G1966), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n697), .A2(new_n698), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n696), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n700), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n702), .B1(new_n696), .B2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT87), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n699), .A2(new_n705), .ZN(new_n706));
  OR3_X1    g281(.A1(new_n697), .A2(new_n698), .A3(new_n705), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n696), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n708), .A2(KEYINPUT20), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n708), .A2(KEYINPUT20), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n704), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  XOR2_X1   g289(.A(G1991), .B(G1996), .Z(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n708), .B(KEYINPUT20), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n717), .A2(new_n704), .A3(new_n712), .ZN(new_n718));
  AND3_X1   g293(.A1(new_n714), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n716), .B1(new_n714), .B2(new_n718), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n693), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n711), .A2(new_n713), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n712), .B1(new_n717), .B2(new_n704), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n715), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n714), .A2(new_n716), .A3(new_n718), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n724), .A2(new_n692), .A3(new_n725), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n721), .A2(new_n726), .ZN(G229));
  NAND2_X1  g302(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT91), .Z(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G29), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G25), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n477), .A2(new_n478), .A3(G131), .ZN(new_n733));
  OAI21_X1  g308(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n734));
  INV_X1    g309(.A(G107), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(G2105), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G119), .B2(new_n480), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n733), .A2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n732), .B1(new_n739), .B2(new_n731), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT35), .B(G1991), .Z(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G16), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G24), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n598), .B2(new_n743), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT88), .B(G1986), .Z(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n742), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(G6), .A2(G16), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G305), .B2(new_n743), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT32), .B(G1981), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(new_n752), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n754), .B(new_n750), .C1(G305), .C2(new_n743), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n743), .B1(new_n510), .B2(new_n525), .ZN(new_n756));
  NOR2_X1   g331(.A1(G16), .A2(G22), .ZN(new_n757));
  OR3_X1    g332(.A1(new_n756), .A2(G1971), .A3(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(G1971), .B1(new_n756), .B2(new_n757), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n753), .A2(new_n755), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n577), .A2(KEYINPUT89), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n577), .A2(KEYINPUT89), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n743), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n743), .A2(G23), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT33), .B(G1976), .ZN(new_n767));
  OR3_X1    g342(.A1(new_n764), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(new_n764), .B2(new_n766), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n760), .A2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT34), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n760), .A2(KEYINPUT34), .A3(new_n770), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n748), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n730), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(new_n776), .ZN(new_n778));
  AND3_X1   g353(.A1(new_n760), .A2(KEYINPUT34), .A3(new_n770), .ZN(new_n779));
  AOI21_X1  g354(.A(KEYINPUT34), .B1(new_n760), .B2(new_n770), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n778), .B(new_n729), .C1(new_n781), .C2(new_n748), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n777), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n731), .A2(G32), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n480), .A2(G129), .ZN(new_n785));
  NAND3_X1  g360(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT26), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n469), .A2(G105), .ZN(new_n789));
  AND3_X1   g364(.A1(new_n785), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n477), .A2(new_n478), .A3(G141), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n784), .B1(new_n793), .B2(new_n731), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT27), .B(G1996), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n794), .A2(new_n796), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n743), .A2(G21), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G168), .B2(new_n743), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n800), .A2(G1966), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT24), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n731), .B1(new_n802), .B2(G34), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(new_n802), .B2(G34), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G160), .B2(G29), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n805), .A2(G2084), .ZN(new_n806));
  NOR4_X1   g381(.A1(new_n797), .A2(new_n798), .A3(new_n801), .A4(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(G4), .A2(G16), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT92), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n613), .B2(new_n743), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G1348), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n731), .A2(G33), .ZN(new_n812));
  INV_X1    g387(.A(G127), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n476), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(G115), .A2(G2104), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(G2105), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(G103), .A2(G2104), .ZN(new_n818));
  OAI21_X1  g393(.A(KEYINPUT93), .B1(new_n818), .B2(G2105), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT93), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n820), .A2(new_n461), .A3(G103), .A4(G2104), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(KEYINPUT25), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT25), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n819), .A2(new_n821), .A3(new_n824), .ZN(new_n825));
  AOI22_X1  g400(.A1(new_n817), .A2(KEYINPUT94), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n477), .A2(new_n478), .A3(G139), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n464), .A2(G127), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n461), .B1(new_n828), .B2(new_n815), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT94), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n826), .A2(new_n827), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n812), .B1(new_n832), .B2(G29), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(G2072), .ZN(new_n834));
  AND3_X1   g409(.A1(new_n807), .A2(new_n811), .A3(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(G5), .A2(G16), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT96), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(G301), .B2(new_n743), .ZN(new_n838));
  INV_X1    g413(.A(G1961), .ZN(new_n839));
  AOI22_X1  g414(.A1(G1966), .A2(new_n800), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n805), .A2(G2084), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n840), .B(new_n841), .C1(new_n839), .C2(new_n838), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT98), .ZN(new_n843));
  NAND2_X1  g418(.A1(G164), .A2(G29), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(G27), .B2(G29), .ZN(new_n845));
  XNOR2_X1  g420(.A(KEYINPUT97), .B(G2078), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n842), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n847), .A2(new_n843), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n743), .A2(G20), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT23), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(new_n618), .B2(new_n743), .ZN(new_n852));
  INV_X1    g427(.A(G1956), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  AND3_X1   g429(.A1(new_n848), .A2(new_n849), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n731), .A2(G35), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n856), .B1(G162), .B2(new_n731), .ZN(new_n857));
  XOR2_X1   g432(.A(KEYINPUT29), .B(G2090), .Z(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(KEYINPUT30), .B(G28), .ZN(new_n860));
  OR2_X1    g435(.A1(KEYINPUT31), .A2(G11), .ZN(new_n861));
  NAND2_X1  g436(.A1(KEYINPUT31), .A2(G11), .ZN(new_n862));
  AOI22_X1  g437(.A1(new_n860), .A2(new_n731), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(new_n637), .B2(new_n731), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(KEYINPUT95), .Z(new_n865));
  NAND2_X1  g440(.A1(new_n743), .A2(G19), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n866), .B1(new_n558), .B2(new_n743), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(G1341), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n731), .A2(G26), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(KEYINPUT28), .Z(new_n870));
  NAND3_X1  g445(.A1(new_n477), .A2(new_n478), .A3(G140), .ZN(new_n871));
  OAI21_X1  g446(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n872));
  INV_X1    g447(.A(G116), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n872), .B1(new_n873), .B2(G2105), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n874), .B1(G128), .B2(new_n480), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n870), .B1(new_n876), .B2(G29), .ZN(new_n877));
  INV_X1    g452(.A(G2067), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  NOR3_X1   g454(.A1(new_n865), .A2(new_n868), .A3(new_n879), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n835), .A2(new_n855), .A3(new_n859), .A4(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(KEYINPUT99), .B1(new_n783), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT99), .ZN(new_n884));
  AOI211_X1 g459(.A(new_n884), .B(new_n881), .C1(new_n777), .C2(new_n782), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n883), .A2(new_n885), .ZN(G311));
  NAND2_X1  g461(.A1(new_n783), .A2(new_n882), .ZN(G150));
  NAND2_X1  g462(.A1(new_n614), .A2(G559), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT38), .ZN(new_n889));
  INV_X1    g464(.A(G67), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n890), .B1(new_n515), .B2(new_n516), .ZN(new_n891));
  NAND2_X1  g466(.A1(G80), .A2(G543), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(G651), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n517), .A2(new_n520), .A3(G93), .ZN(new_n895));
  INV_X1    g470(.A(G55), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(KEYINPUT100), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT100), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(G55), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n523), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n894), .A2(new_n895), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n553), .B1(new_n515), .B2(new_n516), .ZN(new_n902));
  INV_X1    g477(.A(new_n552), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n555), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(G651), .A3(new_n557), .ZN(new_n905));
  INV_X1    g480(.A(new_n551), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n901), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(G93), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n897), .A2(new_n899), .ZN(new_n909));
  OAI22_X1  g484(.A1(new_n501), .A2(new_n908), .B1(new_n503), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(G67), .B1(new_n498), .B2(new_n497), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n506), .B1(new_n911), .B2(new_n892), .ZN(new_n912));
  OAI21_X1  g487(.A(KEYINPUT101), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT101), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n894), .A2(new_n900), .A3(new_n914), .A4(new_n895), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  OAI211_X1 g491(.A(KEYINPUT102), .B(new_n907), .C1(new_n916), .C2(new_n558), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n905), .A2(new_n906), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT102), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n918), .A2(new_n919), .A3(new_n913), .A4(new_n915), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n889), .B(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT39), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(KEYINPUT103), .ZN(new_n925));
  AOI21_X1  g500(.A(G860), .B1(new_n922), .B2(new_n923), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n916), .A2(G860), .ZN(new_n928));
  XOR2_X1   g503(.A(new_n928), .B(KEYINPUT37), .Z(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(G145));
  OR2_X1    g505(.A1(new_n637), .A2(G160), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n637), .A2(G160), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(G162), .B(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n492), .A2(new_n495), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n486), .A2(new_n489), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n831), .A2(new_n827), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n823), .A2(new_n825), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(new_n829), .B2(new_n830), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n937), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n826), .A2(G164), .A3(new_n827), .A4(new_n831), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT105), .B1(new_n733), .B2(new_n737), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n640), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n733), .A2(KEYINPUT105), .A3(new_n737), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n947), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n640), .B1(new_n949), .B2(new_n944), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n943), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n792), .A2(new_n876), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n477), .A2(new_n478), .A3(G142), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n480), .A2(G130), .ZN(new_n955));
  OAI21_X1  g530(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n956), .A2(KEYINPUT104), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(KEYINPUT104), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n958), .B1(G118), .B2(new_n461), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n954), .B(new_n955), .C1(new_n957), .C2(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n790), .A2(new_n791), .A3(new_n871), .A4(new_n875), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n953), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n960), .B1(new_n953), .B2(new_n961), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n941), .A2(new_n942), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n965), .A2(new_n950), .A3(new_n948), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n952), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n964), .B1(new_n952), .B2(new_n966), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n934), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n952), .A2(new_n966), .ZN(new_n971));
  OR2_X1    g546(.A1(new_n962), .A2(new_n963), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n934), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n973), .A2(new_n974), .A3(new_n967), .ZN(new_n975));
  INV_X1    g550(.A(G37), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n970), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n977), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g553(.A(new_n921), .B(new_n624), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n613), .A2(G299), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT41), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n569), .B(KEYINPUT9), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n982), .A2(new_n605), .A3(new_n568), .A4(new_n612), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n980), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT106), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT106), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n980), .A2(new_n986), .A3(new_n983), .A4(new_n981), .ZN(new_n987));
  XNOR2_X1  g562(.A(KEYINPUT107), .B(KEYINPUT41), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n983), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n982), .A2(new_n568), .B1(new_n605), .B2(new_n612), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n989), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n985), .A2(new_n987), .A3(new_n992), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n979), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n979), .B1(new_n991), .B2(new_n990), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  XOR2_X1   g571(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT108), .ZN(new_n999));
  NAND2_X1  g574(.A1(G290), .A2(new_n999), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n594), .A2(new_n999), .A3(new_n597), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n1000), .B(new_n1002), .C1(new_n590), .C2(new_n591), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n598), .A2(KEYINPUT108), .ZN(new_n1004));
  OAI21_X1  g579(.A(G305), .B1(new_n1004), .B2(new_n1001), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n763), .ZN(new_n1007));
  OAI21_X1  g582(.A(G303), .B1(new_n1007), .B2(new_n761), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n763), .B(new_n762), .C1(new_n511), .C2(new_n526), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1003), .A2(new_n1008), .A3(new_n1009), .A4(new_n1005), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n997), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n994), .A2(new_n1015), .A3(new_n995), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n998), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1014), .B1(new_n998), .B2(new_n1016), .ZN(new_n1018));
  OAI21_X1  g593(.A(G868), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n916), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1019), .B1(G868), .B2(new_n1020), .ZN(G295));
  OAI21_X1  g596(.A(new_n1019), .B1(G868), .B2(new_n1020), .ZN(G331));
  INV_X1    g597(.A(G90), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n544), .B1(new_n501), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(G64), .B1(new_n498), .B2(new_n497), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n506), .B1(new_n1025), .B2(new_n541), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT110), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT110), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n543), .A2(new_n1028), .A3(new_n544), .A4(new_n545), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n1027), .A2(G168), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(G168), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1032), .A2(new_n917), .A3(new_n920), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT111), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT111), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1032), .A2(new_n917), .A3(new_n1035), .A4(new_n920), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1032), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n921), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n993), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n990), .A2(new_n991), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1039), .A2(new_n1042), .A3(new_n1033), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1013), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1032), .B1(new_n917), .B2(new_n920), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1045), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n985), .A2(new_n987), .A3(new_n992), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1013), .B(new_n1043), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n976), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT43), .B1(new_n1044), .B2(new_n1049), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n1045), .A2(new_n991), .A3(new_n990), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n1051), .A2(new_n1037), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1039), .A2(new_n1033), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT41), .B1(new_n980), .B2(new_n983), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1054), .B1(new_n1042), .B2(new_n989), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1014), .B1(new_n1052), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT43), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1057), .A2(new_n1058), .A3(new_n976), .A4(new_n1048), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1050), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT44), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AOI22_X1  g637(.A1(new_n1051), .A2(new_n1037), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1048), .B(new_n976), .C1(new_n1013), .C2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1061), .B1(new_n1064), .B2(KEYINPUT43), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT112), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1043), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(new_n1014), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1068), .A2(new_n1058), .A3(new_n976), .A4(new_n1048), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1065), .A2(new_n1066), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1066), .B1(new_n1065), .B2(new_n1069), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1062), .B1(new_n1070), .B2(new_n1071), .ZN(G397));
  INV_X1    g647(.A(G1384), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n937), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G40), .ZN(new_n1075));
  NOR3_X1   g650(.A1(new_n467), .A2(new_n471), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT45), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1074), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  XOR2_X1   g653(.A(new_n1078), .B(KEYINPUT113), .Z(new_n1079));
  AND2_X1   g654(.A1(new_n792), .A2(G1996), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n876), .A2(G2067), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n871), .A2(new_n878), .A3(new_n875), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  OR2_X1    g658(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1078), .A2(G1996), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1079), .A2(new_n1084), .B1(new_n793), .B2(new_n1085), .ZN(new_n1086));
  XOR2_X1   g661(.A(new_n738), .B(new_n741), .Z(new_n1087));
  NAND2_X1  g662(.A1(new_n1079), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1078), .ZN(new_n1090));
  XOR2_X1   g665(.A(new_n598), .B(G1986), .Z(new_n1091));
  AOI21_X1  g666(.A(new_n1089), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G1966), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT115), .B1(G164), .B2(G1384), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT115), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n937), .A2(new_n1095), .A3(new_n1073), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT45), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n937), .A2(KEYINPUT45), .A3(new_n1073), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(new_n1076), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1093), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT116), .B(KEYINPUT50), .Z(new_n1101));
  NAND3_X1  g676(.A1(new_n1094), .A2(new_n1096), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(G125), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n476), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n466), .ZN(new_n1105));
  OAI21_X1  g680(.A(G2105), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1106), .A2(G40), .A3(new_n470), .A4(new_n468), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1107), .B1(new_n1074), .B2(KEYINPUT50), .ZN(new_n1108));
  INV_X1    g683(.A(G2084), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1102), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1100), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(G8), .ZN(new_n1112));
  NOR2_X1   g687(.A1(G168), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT51), .B1(new_n1113), .B2(KEYINPUT121), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1111), .A2(G8), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1113), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1112), .B1(new_n1100), .B2(new_n1110), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1115), .ZN(new_n1120));
  NOR3_X1   g695(.A1(new_n1119), .A2(new_n1113), .A3(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1114), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT62), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n510), .A2(new_n525), .A3(G8), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1124), .B(KEYINPUT55), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1107), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n937), .A2(KEYINPUT114), .A3(KEYINPUT45), .A4(new_n1073), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT114), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1098), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1126), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(G1971), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(G2090), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1102), .A2(new_n1108), .A3(new_n1133), .ZN(new_n1134));
  AOI211_X1 g709(.A(new_n1112), .B(new_n1125), .C1(new_n1132), .C2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(G1976), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n579), .A2(new_n1136), .A3(new_n580), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT52), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1137), .A2(KEYINPUT117), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(KEYINPUT117), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n762), .A2(G1976), .A3(new_n763), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1094), .A2(new_n1096), .A3(new_n1076), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1142), .A2(new_n1143), .A3(G8), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT49), .ZN(new_n1146));
  OAI21_X1  g721(.A(G1981), .B1(new_n585), .B2(new_n588), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  NOR3_X1   g723(.A1(new_n585), .A2(G1981), .A3(new_n588), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1146), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(KEYINPUT118), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT118), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1152), .B(new_n1146), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1149), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1155), .A2(KEYINPUT49), .A3(new_n1147), .ZN(new_n1156));
  AND3_X1   g731(.A1(new_n1143), .A2(G8), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1142), .A2(new_n1143), .A3(G8), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(KEYINPUT52), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1145), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1135), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(G2078), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1126), .A2(new_n1129), .A3(new_n1163), .A4(new_n1127), .ZN(new_n1164));
  XOR2_X1   g739(.A(KEYINPUT123), .B(KEYINPUT53), .Z(new_n1165));
  NAND2_X1  g740(.A1(new_n1102), .A2(new_n1108), .ZN(new_n1166));
  AOI22_X1  g741(.A1(new_n1164), .A2(new_n1165), .B1(new_n1166), .B2(new_n839), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(new_n1077), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n1163), .A2(KEYINPUT53), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1099), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(G301), .B1(new_n1167), .B2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1101), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1076), .B1(new_n1074), .B2(KEYINPUT50), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  AOI22_X1  g751(.A1(new_n1176), .A2(new_n1133), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1125), .B1(new_n1177), .B2(new_n1112), .ZN(new_n1178));
  AND3_X1   g753(.A1(new_n1162), .A2(new_n1173), .A3(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT62), .ZN(new_n1180));
  OAI211_X1 g755(.A(new_n1180), .B(new_n1114), .C1(new_n1118), .C2(new_n1121), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1123), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n581), .A2(new_n1136), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1183), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1184));
  OAI211_X1 g759(.A(G8), .B(new_n1143), .C1(new_n1184), .C2(new_n1149), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1125), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1132), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1134), .ZN(new_n1188));
  OAI211_X1 g763(.A(G8), .B(new_n1186), .C1(new_n1187), .C2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1185), .B1(new_n1189), .B2(new_n1161), .ZN(new_n1190));
  AND3_X1   g765(.A1(new_n1145), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1191));
  AOI211_X1 g766(.A(new_n1112), .B(G286), .C1(new_n1100), .C2(new_n1110), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1191), .A2(new_n1178), .A3(new_n1189), .A4(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT63), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g770(.A(G8), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1196), .A2(new_n1125), .ZN(new_n1197));
  NAND4_X1  g772(.A1(new_n1162), .A2(KEYINPUT63), .A3(new_n1192), .A4(new_n1197), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1190), .B1(new_n1195), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1182), .A2(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g775(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n1201));
  XNOR2_X1  g776(.A(G299), .B(new_n1201), .ZN(new_n1202));
  INV_X1    g777(.A(new_n1202), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n853), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1204));
  XNOR2_X1  g779(.A(KEYINPUT56), .B(G2072), .ZN(new_n1205));
  NAND4_X1  g780(.A1(new_n1126), .A2(new_n1129), .A3(new_n1127), .A4(new_n1205), .ZN(new_n1206));
  AND3_X1   g781(.A1(new_n1203), .A2(new_n1204), .A3(new_n1206), .ZN(new_n1207));
  AOI21_X1  g782(.A(G1348), .B1(new_n1102), .B2(new_n1108), .ZN(new_n1208));
  NOR2_X1   g783(.A1(new_n1143), .A2(G2067), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n614), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1211), .A2(new_n1202), .ZN(new_n1212));
  AOI21_X1  g787(.A(new_n1207), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g788(.A(KEYINPUT61), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1203), .B1(new_n1204), .B2(new_n1206), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n1214), .B1(new_n1207), .B2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g791(.A1(new_n1203), .A2(new_n1204), .A3(new_n1206), .ZN(new_n1217));
  NAND3_X1  g792(.A1(new_n1212), .A2(KEYINPUT61), .A3(new_n1217), .ZN(new_n1218));
  INV_X1    g793(.A(KEYINPUT60), .ZN(new_n1219));
  OR3_X1    g794(.A1(new_n1208), .A2(new_n1209), .A3(new_n1219), .ZN(new_n1220));
  OAI21_X1  g795(.A(new_n1219), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1221));
  NAND3_X1  g796(.A1(new_n1220), .A2(new_n614), .A3(new_n1221), .ZN(new_n1222));
  AND3_X1   g797(.A1(new_n1216), .A2(new_n1218), .A3(new_n1222), .ZN(new_n1223));
  NOR2_X1   g798(.A1(new_n1220), .A2(new_n614), .ZN(new_n1224));
  XOR2_X1   g799(.A(KEYINPUT120), .B(G1996), .Z(new_n1225));
  INV_X1    g800(.A(new_n1143), .ZN(new_n1226));
  XNOR2_X1  g801(.A(KEYINPUT58), .B(G1341), .ZN(new_n1227));
  OAI22_X1  g802(.A1(new_n1130), .A2(new_n1225), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  AND3_X1   g803(.A1(new_n1228), .A2(KEYINPUT59), .A3(new_n558), .ZN(new_n1229));
  AOI21_X1  g804(.A(KEYINPUT59), .B1(new_n1228), .B2(new_n558), .ZN(new_n1230));
  NOR3_X1   g805(.A1(new_n1224), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  AOI21_X1  g806(.A(new_n1213), .B1(new_n1223), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g807(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1233));
  NAND2_X1  g808(.A1(new_n1166), .A2(new_n839), .ZN(new_n1234));
  NAND4_X1  g809(.A1(new_n1126), .A2(new_n1129), .A3(new_n1127), .A4(new_n1170), .ZN(new_n1235));
  NAND3_X1  g810(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1236));
  NAND2_X1  g811(.A1(new_n1236), .A2(G171), .ZN(new_n1237));
  NAND2_X1  g812(.A1(new_n1237), .A2(KEYINPUT124), .ZN(new_n1238));
  NAND4_X1  g813(.A1(new_n1233), .A2(new_n1234), .A3(new_n1172), .A4(G301), .ZN(new_n1239));
  AND2_X1   g814(.A1(new_n1239), .A2(KEYINPUT54), .ZN(new_n1240));
  INV_X1    g815(.A(KEYINPUT124), .ZN(new_n1241));
  NAND3_X1  g816(.A1(new_n1236), .A2(new_n1241), .A3(G171), .ZN(new_n1242));
  NAND3_X1  g817(.A1(new_n1238), .A2(new_n1240), .A3(new_n1242), .ZN(new_n1243));
  INV_X1    g818(.A(new_n1175), .ZN(new_n1244));
  INV_X1    g819(.A(new_n1168), .ZN(new_n1245));
  OAI211_X1 g820(.A(new_n1244), .B(new_n1133), .C1(new_n1245), .C2(new_n1101), .ZN(new_n1246));
  NAND2_X1  g821(.A1(new_n1246), .A2(new_n1132), .ZN(new_n1247));
  AOI21_X1  g822(.A(new_n1186), .B1(new_n1247), .B2(G8), .ZN(new_n1248));
  NOR3_X1   g823(.A1(new_n1248), .A2(new_n1135), .A3(new_n1161), .ZN(new_n1249));
  XOR2_X1   g824(.A(KEYINPUT122), .B(KEYINPUT54), .Z(new_n1250));
  NOR2_X1   g825(.A1(new_n1236), .A2(G171), .ZN(new_n1251));
  OAI21_X1  g826(.A(new_n1250), .B1(new_n1251), .B2(new_n1173), .ZN(new_n1252));
  NAND4_X1  g827(.A1(new_n1243), .A2(new_n1122), .A3(new_n1249), .A4(new_n1252), .ZN(new_n1253));
  NOR2_X1   g828(.A1(new_n1232), .A2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g829(.A(new_n1092), .B1(new_n1200), .B2(new_n1254), .ZN(new_n1255));
  OAI21_X1  g830(.A(new_n1079), .B1(new_n792), .B2(new_n1083), .ZN(new_n1256));
  INV_X1    g831(.A(KEYINPUT46), .ZN(new_n1257));
  INV_X1    g832(.A(new_n1085), .ZN(new_n1258));
  OAI21_X1  g833(.A(new_n1256), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g834(.A1(new_n1258), .A2(new_n1257), .ZN(new_n1260));
  XNOR2_X1  g835(.A(new_n1260), .B(KEYINPUT126), .ZN(new_n1261));
  NOR2_X1   g836(.A1(new_n1259), .A2(new_n1261), .ZN(new_n1262));
  XNOR2_X1  g837(.A(new_n1262), .B(KEYINPUT47), .ZN(new_n1263));
  NAND2_X1  g838(.A1(new_n739), .A2(new_n741), .ZN(new_n1264));
  XNOR2_X1  g839(.A(new_n1264), .B(KEYINPUT125), .ZN(new_n1265));
  NAND2_X1  g840(.A1(new_n1086), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g841(.A1(new_n1266), .A2(new_n1082), .ZN(new_n1267));
  AND2_X1   g842(.A1(new_n1267), .A2(new_n1079), .ZN(new_n1268));
  NOR3_X1   g843(.A1(new_n1078), .A2(G1986), .A3(G290), .ZN(new_n1269));
  XOR2_X1   g844(.A(new_n1269), .B(KEYINPUT48), .Z(new_n1270));
  AND3_X1   g845(.A1(new_n1270), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1271));
  NOR3_X1   g846(.A1(new_n1263), .A2(new_n1268), .A3(new_n1271), .ZN(new_n1272));
  NAND2_X1  g847(.A1(new_n1255), .A2(new_n1272), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g848(.A(KEYINPUT127), .ZN(new_n1275));
  NAND3_X1  g849(.A1(new_n690), .A2(new_n667), .A3(G319), .ZN(new_n1276));
  AOI21_X1  g850(.A(new_n1276), .B1(new_n721), .B2(new_n726), .ZN(new_n1277));
  NAND2_X1  g851(.A1(new_n977), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g852(.A(new_n1278), .ZN(new_n1279));
  AOI21_X1  g853(.A(new_n1275), .B1(new_n1060), .B2(new_n1279), .ZN(new_n1280));
  AOI211_X1 g854(.A(KEYINPUT127), .B(new_n1278), .C1(new_n1050), .C2(new_n1059), .ZN(new_n1281));
  NOR2_X1   g855(.A1(new_n1280), .A2(new_n1281), .ZN(G308));
  NAND2_X1  g856(.A1(new_n1060), .A2(new_n1279), .ZN(G225));
endmodule


