//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 0 1 1 1 0 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 0 1 1 1 1 0 0 0 1 0 0 0 0 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961;
  XNOR2_X1  g000(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XNOR2_X1  g002(.A(G127gat), .B(G155gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(G211gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G231gat), .ZN(new_n207));
  INV_X1    g006(.A(G233gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G64gat), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n210), .A2(G57gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(G57gat), .ZN(new_n212));
  INV_X1    g011(.A(G71gat), .ZN(new_n213));
  INV_X1    g012(.A(G78gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT9), .ZN(new_n215));
  NAND2_X1  g014(.A1(G71gat), .A2(G78gat), .ZN(new_n216));
  AOI22_X1  g015(.A1(new_n211), .A2(new_n212), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT9), .ZN(new_n218));
  AOI22_X1  g017(.A1(new_n211), .A2(new_n212), .B1(new_n218), .B2(new_n216), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT96), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT95), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n222), .A2(new_n213), .A3(new_n214), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT95), .B1(G71gat), .B2(G78gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n221), .B1(new_n225), .B2(new_n216), .ZN(new_n226));
  AND2_X1   g025(.A1(G71gat), .A2(G78gat), .ZN(new_n227));
  AOI211_X1 g026(.A(KEYINPUT96), .B(new_n227), .C1(new_n223), .C2(new_n224), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n220), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT97), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI211_X1 g030(.A(KEYINPUT97), .B(new_n220), .C1(new_n226), .C2(new_n228), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n217), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n233), .A2(KEYINPUT21), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(KEYINPUT21), .ZN(new_n235));
  INV_X1    g034(.A(G183gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(G15gat), .B(G22gat), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT16), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n237), .B1(new_n238), .B2(G1gat), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n239), .B1(G1gat), .B2(new_n237), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n240), .B(G8gat), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n235), .A2(new_n236), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n236), .B1(new_n235), .B2(new_n242), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n234), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n245), .ZN(new_n247));
  INV_X1    g046(.A(new_n234), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n247), .A2(new_n243), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n209), .B1(new_n246), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n246), .A2(new_n249), .A3(new_n209), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n206), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n252), .ZN(new_n254));
  NOR3_X1   g053(.A1(new_n254), .A2(new_n250), .A3(new_n205), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n203), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n251), .A2(new_n206), .A3(new_n252), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n205), .B1(new_n254), .B2(new_n250), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n257), .A2(new_n258), .A3(new_n202), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT100), .ZN(new_n261));
  XNOR2_X1  g060(.A(G43gat), .B(G50gat), .ZN(new_n262));
  OR2_X1    g061(.A1(new_n262), .A2(KEYINPUT91), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(KEYINPUT91), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(KEYINPUT15), .A3(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT92), .ZN(new_n266));
  INV_X1    g065(.A(G29gat), .ZN(new_n267));
  INV_X1    g066(.A(G36gat), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT92), .B1(G29gat), .B2(G36gat), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(KEYINPUT14), .A3(new_n270), .ZN(new_n271));
  OAI221_X1 g070(.A(new_n271), .B1(KEYINPUT14), .B2(new_n270), .C1(new_n267), .C2(new_n268), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n265), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(KEYINPUT93), .B(KEYINPUT15), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n262), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT91), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n262), .B(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n275), .B1(new_n277), .B2(KEYINPUT15), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n273), .B1(new_n278), .B2(new_n272), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  XOR2_X1   g079(.A(G99gat), .B(G106gat), .Z(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(G85gat), .ZN(new_n283));
  INV_X1    g082(.A(G92gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G85gat), .A2(G92gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n286), .B(KEYINPUT7), .ZN(new_n287));
  INV_X1    g086(.A(G99gat), .ZN(new_n288));
  INV_X1    g087(.A(G106gat), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT8), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n282), .A2(new_n285), .A3(new_n287), .A4(new_n290), .ZN(new_n291));
  AND2_X1   g090(.A1(new_n286), .A2(KEYINPUT7), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n286), .A2(KEYINPUT7), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n285), .B(new_n290), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(new_n281), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  AND2_X1   g096(.A1(G232gat), .A2(G233gat), .ZN(new_n298));
  AOI22_X1  g097(.A1(new_n280), .A2(new_n297), .B1(KEYINPUT41), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n275), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n272), .B1(new_n265), .B2(new_n300), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n265), .A2(new_n272), .ZN(new_n302));
  OAI21_X1  g101(.A(KEYINPUT17), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT17), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n304), .B(new_n273), .C1(new_n278), .C2(new_n272), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n303), .A2(new_n296), .A3(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(G190gat), .B(G218gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n307), .B(KEYINPUT101), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT102), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n299), .A2(new_n306), .A3(new_n310), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n309), .A2(KEYINPUT102), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n261), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n312), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n314), .B1(new_n299), .B2(new_n306), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n298), .A2(KEYINPUT41), .ZN(new_n316));
  XNOR2_X1  g115(.A(G134gat), .B(G162gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n316), .B(new_n317), .ZN(new_n318));
  XOR2_X1   g117(.A(KEYINPUT98), .B(KEYINPUT99), .Z(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  OR3_X1    g120(.A1(new_n313), .A2(new_n315), .A3(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n321), .B1(new_n313), .B2(new_n315), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  AND2_X1   g124(.A1(G226gat), .A2(G233gat), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT65), .ZN(new_n327));
  NAND2_X1  g126(.A1(G169gat), .A2(G176gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT64), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT64), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n330), .A2(G169gat), .A3(G176gat), .ZN(new_n331));
  AND2_X1   g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(G169gat), .ZN(new_n333));
  INV_X1    g132(.A(G176gat), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n333), .A2(new_n334), .A3(KEYINPUT23), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT23), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n336), .B1(G169gat), .B2(G176gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n327), .B1(new_n332), .B2(new_n338), .ZN(new_n339));
  NOR2_X1   g138(.A1(G183gat), .A2(G190gat), .ZN(new_n340));
  INV_X1    g139(.A(G190gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n236), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n340), .B1(new_n342), .B2(KEYINPUT24), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n343), .B1(KEYINPUT24), .B2(new_n342), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n331), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n345), .A2(KEYINPUT65), .A3(new_n337), .A4(new_n335), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n339), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT25), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n236), .A2(KEYINPUT67), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT67), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(G183gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n352), .A2(new_n341), .B1(KEYINPUT24), .B2(new_n342), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT66), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n354), .B(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n348), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n332), .A2(new_n338), .ZN(new_n358));
  AOI22_X1  g157(.A1(new_n347), .A2(new_n348), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT67), .B(G183gat), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT27), .ZN(new_n361));
  OAI21_X1  g160(.A(KEYINPUT68), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT68), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n352), .A2(new_n363), .A3(KEYINPUT27), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT28), .B1(new_n361), .B2(G183gat), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n362), .A2(new_n364), .A3(new_n341), .A4(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n342), .ZN(new_n367));
  XOR2_X1   g166(.A(KEYINPUT27), .B(G183gat), .Z(new_n368));
  OAI21_X1  g167(.A(KEYINPUT28), .B1(new_n368), .B2(G190gat), .ZN(new_n369));
  OR4_X1    g168(.A1(KEYINPUT69), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n333), .A2(new_n334), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT69), .B1(new_n371), .B2(KEYINPUT26), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(KEYINPUT26), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n370), .A2(new_n372), .A3(new_n345), .A4(new_n373), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n366), .A2(new_n367), .A3(new_n369), .A4(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n326), .B1(new_n359), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n347), .A2(new_n348), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n357), .A2(new_n358), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT29), .B1(new_n380), .B2(new_n375), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n377), .B1(new_n381), .B2(new_n326), .ZN(new_n382));
  XNOR2_X1  g181(.A(G197gat), .B(G204gat), .ZN(new_n383));
  INV_X1    g182(.A(G211gat), .ZN(new_n384));
  INV_X1    g183(.A(G218gat), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n383), .B1(KEYINPUT22), .B2(new_n386), .ZN(new_n387));
  XOR2_X1   g186(.A(G211gat), .B(G218gat), .Z(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n387), .B(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n382), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT74), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n387), .B(new_n388), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n377), .B(new_n393), .C1(new_n381), .C2(new_n326), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n391), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  OR2_X1    g194(.A1(new_n394), .A2(new_n392), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(G8gat), .B(G36gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(G64gat), .B(G92gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n397), .A2(KEYINPUT30), .A3(new_n401), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT75), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n400), .B1(new_n395), .B2(new_n396), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT75), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT30), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n402), .B1(new_n404), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT35), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT76), .ZN(new_n410));
  INV_X1    g209(.A(G141gat), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n411), .A2(G148gat), .ZN(new_n412));
  INV_X1    g211(.A(G148gat), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n413), .A2(G141gat), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n410), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(G155gat), .A2(G162gat), .ZN(new_n416));
  INV_X1    g215(.A(G155gat), .ZN(new_n417));
  INV_X1    g216(.A(G162gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n416), .B1(new_n419), .B2(KEYINPUT2), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n413), .A2(G141gat), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n411), .A2(G148gat), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(new_n422), .A3(KEYINPUT76), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n415), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G141gat), .B(G148gat), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n416), .B(new_n419), .C1(new_n425), .C2(KEYINPUT2), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT77), .B(KEYINPUT3), .ZN(new_n427));
  AND3_X1   g226(.A1(new_n424), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  OR2_X1    g227(.A1(G127gat), .A2(G134gat), .ZN(new_n429));
  NAND2_X1  g228(.A1(G127gat), .A2(G134gat), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT1), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(G113gat), .ZN(new_n432));
  OR2_X1    g231(.A1(KEYINPUT70), .A2(G120gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(KEYINPUT70), .A2(G120gat), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(G120gat), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n436), .A2(G113gat), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n431), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  XNOR2_X1  g237(.A(G113gat), .B(G120gat), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n429), .B(new_n430), .C1(new_n439), .C2(KEYINPUT1), .ZN(new_n440));
  AND2_X1   g239(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT3), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n442), .B1(new_n424), .B2(new_n426), .ZN(new_n443));
  NOR3_X1   g242(.A1(new_n428), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n446));
  NAND2_X1  g245(.A1(G225gat), .A2(G233gat), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n441), .A2(KEYINPUT4), .A3(new_n424), .A4(new_n426), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n438), .A2(new_n440), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n424), .A2(new_n426), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT78), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n424), .A2(KEYINPUT78), .A3(new_n426), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n451), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n450), .B1(new_n456), .B2(KEYINPUT4), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT80), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n424), .A2(KEYINPUT78), .A3(new_n426), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT78), .B1(new_n424), .B2(new_n426), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n441), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT4), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT80), .B1(new_n464), .B2(new_n450), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n445), .B(new_n449), .C1(new_n459), .C2(new_n465), .ZN(new_n466));
  OAI22_X1  g265(.A1(new_n444), .A2(new_n463), .B1(new_n452), .B2(new_n451), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n456), .A2(KEYINPUT4), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n467), .A2(new_n447), .A3(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n441), .B(new_n452), .ZN(new_n470));
  OR2_X1    g269(.A1(new_n470), .A2(new_n447), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n469), .A2(new_n471), .A3(new_n446), .ZN(new_n472));
  XNOR2_X1  g271(.A(G1gat), .B(G29gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n473), .B(G85gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(KEYINPUT0), .B(G57gat), .ZN(new_n475));
  XOR2_X1   g274(.A(new_n474), .B(new_n475), .Z(new_n476));
  NAND3_X1  g275(.A1(new_n466), .A2(new_n472), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT81), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n466), .A2(new_n472), .ZN(new_n480));
  INV_X1    g279(.A(new_n476), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT6), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n466), .A2(new_n472), .A3(KEYINPUT81), .A4(new_n476), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n479), .A2(new_n482), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n480), .A2(KEYINPUT6), .A3(new_n481), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OR2_X1    g286(.A1(new_n405), .A2(KEYINPUT30), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n408), .A2(new_n409), .A3(new_n487), .A4(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(G228gat), .A2(G233gat), .ZN(new_n490));
  INV_X1    g289(.A(new_n428), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT29), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT86), .ZN(new_n494));
  OR3_X1    g293(.A1(new_n428), .A2(KEYINPUT86), .A3(KEYINPUT29), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n490), .B1(new_n496), .B2(new_n390), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n442), .B1(new_n390), .B2(KEYINPUT29), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(new_n452), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT85), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT85), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n498), .A2(new_n501), .A3(new_n452), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n497), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(KEYINPUT87), .B(G22gat), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n490), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n493), .A2(new_n390), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n427), .B1(new_n390), .B2(KEYINPUT29), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n460), .A2(new_n461), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n507), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT84), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n512), .A2(KEYINPUT84), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n504), .B(new_n506), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G78gat), .B(G106gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(KEYINPUT31), .B(G50gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(G22gat), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT84), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n508), .A2(new_n511), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n521), .B1(new_n522), .B2(new_n507), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n523), .A2(new_n513), .B1(new_n497), .B2(new_n503), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n516), .B(new_n519), .C1(new_n520), .C2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  XOR2_X1   g325(.A(new_n519), .B(KEYINPUT83), .Z(new_n527));
  OAI21_X1  g326(.A(new_n504), .B1(new_n514), .B2(new_n515), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(new_n505), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n527), .B1(new_n529), .B2(new_n516), .ZN(new_n530));
  OR2_X1    g329(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(G227gat), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n532), .A2(new_n208), .ZN(new_n533));
  NOR3_X1   g332(.A1(new_n359), .A2(new_n376), .A3(new_n451), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n441), .B1(new_n380), .B2(new_n375), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT33), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n536), .A2(KEYINPUT71), .A3(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT71), .ZN(new_n539));
  INV_X1    g338(.A(new_n533), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n451), .B1(new_n359), .B2(new_n376), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n380), .A2(new_n441), .A3(new_n375), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n539), .B1(new_n543), .B2(KEYINPUT33), .ZN(new_n544));
  XOR2_X1   g343(.A(G15gat), .B(G43gat), .Z(new_n545));
  XNOR2_X1  g344(.A(G71gat), .B(G99gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n536), .A2(KEYINPUT32), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n538), .A2(new_n544), .A3(new_n547), .A4(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(KEYINPUT33), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n536), .A2(KEYINPUT32), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n541), .A2(new_n542), .A3(new_n540), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT34), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n554), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n549), .A2(new_n556), .A3(new_n551), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n555), .A2(KEYINPUT73), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT73), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n552), .A2(new_n559), .A3(new_n554), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n531), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(KEYINPUT90), .B1(new_n489), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n402), .ZN(new_n564));
  AND4_X1   g363(.A1(new_n406), .A2(new_n397), .A3(KEYINPUT30), .A4(new_n401), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n406), .B1(new_n405), .B2(KEYINPUT30), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n488), .B(new_n564), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  AND2_X1   g366(.A1(new_n485), .A2(new_n486), .ZN(new_n568));
  NOR3_X1   g367(.A1(new_n567), .A2(new_n568), .A3(KEYINPUT35), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT90), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n526), .A2(new_n530), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n571), .B1(new_n560), .B2(new_n558), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n569), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n555), .A2(new_n557), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n531), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT82), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n576), .B1(new_n567), .B2(new_n568), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n408), .A2(KEYINPUT82), .A3(new_n487), .A4(new_n488), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n575), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI211_X1 g378(.A(new_n563), .B(new_n573), .C1(new_n579), .C2(new_n409), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT36), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n558), .A2(new_n581), .A3(new_n560), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n555), .A2(KEYINPUT36), .A3(new_n557), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(KEYINPUT72), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT72), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n577), .A2(new_n578), .A3(new_n571), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n470), .A2(new_n447), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n457), .A2(new_n458), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n464), .A2(KEYINPUT80), .A3(new_n450), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n444), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  OAI211_X1 g392(.A(KEYINPUT39), .B(new_n590), .C1(new_n593), .C2(new_n447), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n445), .B1(new_n459), .B2(new_n465), .ZN(new_n595));
  XNOR2_X1  g394(.A(KEYINPUT88), .B(KEYINPUT39), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n595), .A2(new_n448), .A3(new_n596), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n594), .A2(new_n597), .A3(KEYINPUT40), .A4(new_n476), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(new_n482), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n594), .A2(new_n476), .A3(new_n597), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT40), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n567), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n391), .A2(new_n394), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n401), .B1(new_n604), .B2(KEYINPUT37), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT38), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT37), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT89), .B1(new_n397), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT89), .ZN(new_n609));
  AOI211_X1 g408(.A(new_n609), .B(KEYINPUT37), .C1(new_n395), .C2(new_n396), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n605), .B(new_n606), .C1(new_n608), .C2(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n401), .B1(new_n397), .B2(KEYINPUT38), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n568), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  OR2_X1    g412(.A1(new_n608), .A2(new_n610), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n395), .A2(KEYINPUT37), .A3(new_n396), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n606), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n531), .B(new_n603), .C1(new_n613), .C2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n588), .A2(new_n589), .A3(new_n617), .ZN(new_n618));
  AOI211_X1 g417(.A(new_n260), .B(new_n325), .C1(new_n580), .C2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G230gat), .A2(G233gat), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n217), .ZN(new_n622));
  INV_X1    g421(.A(new_n224), .ZN(new_n623));
  NOR3_X1   g422(.A1(KEYINPUT95), .A2(G71gat), .A3(G78gat), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n216), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT96), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n225), .A2(new_n221), .A3(new_n216), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(KEYINPUT97), .B1(new_n628), .B2(new_n220), .ZN(new_n629));
  AOI211_X1 g428(.A(new_n230), .B(new_n219), .C1(new_n626), .C2(new_n627), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n622), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(new_n296), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n233), .A2(new_n297), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT103), .B(KEYINPUT10), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  AOI211_X1 g434(.A(new_n217), .B(new_n296), .C1(new_n231), .C2(new_n232), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(KEYINPUT10), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n621), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n620), .B1(new_n632), .B2(new_n633), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G120gat), .B(G148gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(G176gat), .B(G204gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n638), .A2(new_n639), .A3(new_n643), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n303), .A2(new_n242), .A3(new_n305), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n280), .A2(new_n241), .ZN(new_n650));
  NAND2_X1  g449(.A1(G229gat), .A2(G233gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT94), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n649), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT18), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n242), .A2(new_n279), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n650), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n652), .B(KEYINPUT13), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n649), .A2(new_n650), .A3(KEYINPUT18), .A4(new_n652), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n655), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(G113gat), .B(G141gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(G197gat), .ZN(new_n664));
  XOR2_X1   g463(.A(KEYINPUT11), .B(G169gat), .Z(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT12), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n655), .A2(new_n667), .A3(new_n660), .A4(new_n661), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n648), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n619), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n568), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(G1gat), .ZN(G1324gat));
  NAND3_X1  g476(.A1(new_n619), .A2(new_n673), .A3(new_n567), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT42), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT16), .B(G8gat), .ZN(new_n680));
  OR3_X1    g479(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n678), .B(KEYINPUT104), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n679), .B1(new_n682), .B2(G8gat), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n682), .A2(new_n680), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n681), .B1(new_n683), .B2(new_n684), .ZN(G1325gat));
  INV_X1    g484(.A(new_n588), .ZN(new_n686));
  AND3_X1   g485(.A1(new_n675), .A2(G15gat), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(G15gat), .B1(new_n675), .B2(new_n561), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(G1326gat));
  NOR2_X1   g488(.A1(new_n674), .A2(new_n531), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT43), .B(G22gat), .Z(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1327gat));
  AOI21_X1  g491(.A(new_n324), .B1(new_n580), .B2(new_n618), .ZN(new_n693));
  AND3_X1   g492(.A1(new_n693), .A2(new_n673), .A3(new_n260), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n694), .A2(new_n267), .A3(new_n568), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT45), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n613), .A2(new_n616), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n603), .A2(new_n531), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n586), .B1(new_n582), .B2(new_n583), .ZN(new_n700));
  INV_X1    g499(.A(new_n587), .ZN(new_n701));
  OAI22_X1  g500(.A1(new_n698), .A2(new_n699), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n589), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n697), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n588), .A2(KEYINPUT107), .A3(new_n589), .A4(new_n617), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n704), .A2(new_n580), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(KEYINPUT44), .B1(new_n706), .B2(new_n325), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  AOI211_X1 g507(.A(new_n708), .B(new_n324), .C1(new_n580), .C2(new_n618), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n256), .A2(new_n259), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n647), .B(KEYINPUT105), .Z(new_n712));
  NOR3_X1   g511(.A1(new_n711), .A2(new_n672), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT106), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n710), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(G29gat), .B1(new_n715), .B2(new_n487), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n696), .A2(new_n716), .ZN(G1328gat));
  INV_X1    g516(.A(new_n567), .ZN(new_n718));
  OAI21_X1  g517(.A(G36gat), .B1(new_n715), .B2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n694), .A2(new_n268), .A3(new_n567), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT46), .ZN(new_n721));
  OR2_X1    g520(.A1(new_n720), .A2(KEYINPUT46), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n719), .A2(new_n721), .A3(new_n722), .ZN(G1329gat));
  AOI21_X1  g522(.A(G43gat), .B1(new_n558), .B2(new_n560), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n694), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n706), .A2(new_n325), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n708), .ZN(new_n727));
  INV_X1    g526(.A(new_n709), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n727), .A2(new_n728), .A3(new_n686), .A4(new_n714), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n725), .B1(new_n729), .B2(G43gat), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g530(.A1(new_n710), .A2(G50gat), .A3(new_n571), .A4(new_n714), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n694), .A2(new_n571), .ZN(new_n733));
  INV_X1    g532(.A(G50gat), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n732), .A2(KEYINPUT48), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(KEYINPUT48), .B1(new_n732), .B2(new_n735), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(G1331gat));
  NAND4_X1  g537(.A1(new_n711), .A2(new_n672), .A3(new_n324), .A4(new_n712), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT108), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n706), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n741), .A2(new_n487), .ZN(new_n742));
  XNOR2_X1  g541(.A(KEYINPUT109), .B(G57gat), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(G1332gat));
  INV_X1    g543(.A(new_n741), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n718), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n746), .B(KEYINPUT110), .Z(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT111), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT111), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n745), .A2(new_n750), .A3(new_n747), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(G1333gat));
  OAI21_X1  g553(.A(G71gat), .B1(new_n741), .B2(new_n588), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n561), .A2(new_n213), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n755), .B1(new_n741), .B2(new_n756), .ZN(new_n757));
  XOR2_X1   g556(.A(new_n757), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g557(.A1(new_n741), .A2(new_n531), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(new_n214), .ZN(G1335gat));
  NOR2_X1   g559(.A1(new_n711), .A2(new_n671), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(new_n648), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n707), .A2(new_n709), .A3(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(G85gat), .B1(new_n764), .B2(new_n487), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n706), .A2(new_n325), .A3(new_n761), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n706), .A2(KEYINPUT51), .A3(new_n325), .A4(new_n761), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n770), .A2(new_n283), .A3(new_n568), .A4(new_n648), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n765), .A2(new_n771), .ZN(G1336gat));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n773));
  NOR4_X1   g572(.A1(new_n707), .A2(new_n718), .A3(new_n709), .A4(new_n762), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n773), .B1(new_n774), .B2(new_n284), .ZN(new_n775));
  INV_X1    g574(.A(new_n712), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n718), .A2(G92gat), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  AOI211_X1 g577(.A(new_n776), .B(new_n778), .C1(new_n768), .C2(new_n769), .ZN(new_n779));
  OAI21_X1  g578(.A(KEYINPUT52), .B1(new_n775), .B2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n762), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n710), .A2(new_n567), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(G92gat), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n770), .A2(new_n712), .A3(new_n777), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n783), .A2(new_n784), .A3(new_n773), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n780), .A2(new_n786), .ZN(G1337gat));
  OAI21_X1  g586(.A(G99gat), .B1(new_n764), .B2(new_n588), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n770), .A2(new_n288), .A3(new_n648), .A4(new_n561), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(G1338gat));
  NAND2_X1  g589(.A1(new_n763), .A2(new_n571), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(G106gat), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n770), .A2(new_n289), .A3(new_n571), .A4(new_n712), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n289), .B1(new_n763), .B2(new_n571), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n571), .A2(new_n289), .ZN(new_n797));
  AOI211_X1 g596(.A(new_n776), .B(new_n797), .C1(new_n768), .C2(new_n769), .ZN(new_n798));
  OAI21_X1  g597(.A(KEYINPUT53), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n795), .A2(new_n799), .ZN(G1339gat));
  NOR2_X1   g599(.A1(new_n567), .A2(new_n487), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n635), .A2(new_n621), .A3(new_n637), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(KEYINPUT54), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n805), .A2(new_n638), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n233), .A2(new_n297), .ZN(new_n808));
  INV_X1    g607(.A(new_n634), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n808), .A2(new_n636), .A3(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n637), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n807), .B(new_n620), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n643), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n803), .B1(new_n806), .B2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n646), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n620), .B1(new_n810), .B2(new_n811), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n816), .A2(KEYINPUT54), .A3(new_n804), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n644), .B1(new_n638), .B2(new_n807), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n817), .A2(new_n818), .A3(KEYINPUT55), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n814), .A2(new_n815), .A3(new_n671), .A4(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n657), .A2(new_n659), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n652), .B1(new_n649), .B2(new_n650), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n666), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n670), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n824), .B1(new_n645), .B2(new_n646), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n820), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n324), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT113), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n814), .A2(new_n815), .A3(new_n824), .A4(new_n819), .ZN(new_n829));
  OR2_X1    g628(.A1(new_n829), .A2(new_n324), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n827), .A2(new_n828), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n325), .B1(new_n820), .B2(new_n825), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n829), .A2(new_n324), .ZN(new_n833));
  OAI21_X1  g632(.A(KEYINPUT113), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n831), .A2(new_n260), .A3(new_n834), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n711), .A2(new_n647), .A3(new_n672), .A4(new_n324), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n802), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n572), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(KEYINPUT114), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(G113gat), .B1(new_n840), .B2(new_n672), .ZN(new_n841));
  INV_X1    g640(.A(new_n575), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n837), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n843), .A2(new_n432), .A3(new_n671), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n841), .A2(new_n844), .ZN(G1340gat));
  OAI21_X1  g644(.A(G120gat), .B1(new_n840), .B2(new_n776), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n647), .B1(new_n433), .B2(new_n434), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(G1341gat));
  AOI21_X1  g648(.A(G127gat), .B1(new_n843), .B2(new_n711), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n711), .A2(G127gat), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n850), .B1(new_n839), .B2(new_n851), .ZN(G1342gat));
  OAI21_X1  g651(.A(G134gat), .B1(new_n840), .B2(new_n324), .ZN(new_n853));
  INV_X1    g652(.A(G134gat), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n843), .A2(new_n854), .A3(new_n325), .ZN(new_n855));
  XOR2_X1   g654(.A(KEYINPUT115), .B(KEYINPUT56), .Z(new_n856));
  XNOR2_X1  g655(.A(new_n855), .B(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n853), .A2(new_n857), .ZN(G1343gat));
  NOR4_X1   g657(.A1(new_n260), .A2(new_n648), .A3(new_n671), .A4(new_n325), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n646), .B1(new_n669), .B2(new_n670), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n817), .A2(new_n818), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n861), .A2(KEYINPUT116), .A3(new_n803), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n861), .A2(KEYINPUT116), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n860), .B(new_n862), .C1(new_n863), .C2(new_n803), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT117), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n864), .A2(new_n865), .A3(new_n825), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n324), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n865), .B1(new_n864), .B2(new_n825), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n830), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n859), .B1(new_n869), .B2(new_n260), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT57), .B1(new_n870), .B2(new_n531), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n531), .B1(new_n835), .B2(new_n836), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT57), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n686), .A2(new_n802), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n871), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(G141gat), .B1(new_n876), .B2(new_n672), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n875), .A2(new_n872), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n671), .A2(new_n411), .ZN(new_n879));
  XOR2_X1   g678(.A(new_n879), .B(KEYINPUT118), .Z(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(KEYINPUT58), .ZN(G1344gat));
  NAND3_X1  g682(.A1(new_n878), .A2(new_n413), .A3(new_n648), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT59), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n885), .B(G148gat), .C1(new_n876), .C2(new_n647), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n886), .B(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n873), .B1(new_n870), .B2(new_n531), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n872), .A2(KEYINPUT57), .ZN(new_n892));
  OAI211_X1 g691(.A(KEYINPUT120), .B(new_n873), .C1(new_n870), .C2(new_n531), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n648), .A3(new_n875), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n885), .B1(new_n895), .B2(G148gat), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n884), .B1(new_n888), .B2(new_n896), .ZN(G1345gat));
  AOI21_X1  g696(.A(G155gat), .B1(new_n878), .B2(new_n711), .ZN(new_n898));
  INV_X1    g697(.A(new_n876), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n260), .A2(new_n417), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(G1346gat));
  AOI21_X1  g700(.A(G162gat), .B1(new_n878), .B2(new_n325), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n324), .A2(new_n418), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(new_n899), .B2(new_n903), .ZN(G1347gat));
  NAND2_X1  g703(.A1(new_n835), .A2(new_n836), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n561), .A2(new_n567), .A3(new_n487), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT122), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n905), .A2(new_n531), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(G169gat), .B1(new_n908), .B2(new_n672), .ZN(new_n909));
  XOR2_X1   g708(.A(new_n909), .B(KEYINPUT123), .Z(new_n910));
  AOI21_X1  g709(.A(KEYINPUT121), .B1(new_n905), .B2(new_n487), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n912));
  AOI211_X1 g711(.A(new_n912), .B(new_n568), .C1(new_n835), .C2(new_n836), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n567), .B(new_n842), .C1(new_n911), .C2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n915), .A2(new_n333), .A3(new_n671), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n910), .A2(new_n916), .ZN(G1348gat));
  NOR3_X1   g716(.A1(new_n908), .A2(new_n334), .A3(new_n776), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n915), .A2(new_n648), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(new_n334), .ZN(G1349gat));
  OAI21_X1  g719(.A(new_n360), .B1(new_n908), .B2(new_n260), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT124), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n914), .A2(new_n260), .ZN(new_n923));
  INV_X1    g722(.A(new_n368), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NOR4_X1   g724(.A1(new_n914), .A2(KEYINPUT124), .A3(new_n368), .A4(new_n260), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n921), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(KEYINPUT60), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT60), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n929), .B(new_n921), .C1(new_n925), .C2(new_n926), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(G1350gat));
  NAND3_X1  g730(.A1(new_n915), .A2(new_n341), .A3(new_n325), .ZN(new_n932));
  OAI21_X1  g731(.A(G190gat), .B1(new_n908), .B2(new_n324), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT61), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(G1351gat));
  NOR3_X1   g734(.A1(new_n686), .A2(new_n568), .A3(new_n718), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n894), .A2(new_n671), .A3(new_n936), .ZN(new_n937));
  XOR2_X1   g736(.A(KEYINPUT125), .B(G197gat), .Z(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n911), .A2(new_n913), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n588), .A2(new_n571), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n940), .A2(new_n718), .A3(new_n941), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n672), .A2(new_n938), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n939), .A2(new_n944), .ZN(G1352gat));
  INV_X1    g744(.A(G204gat), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n942), .A2(new_n946), .A3(new_n648), .ZN(new_n947));
  OR2_X1    g746(.A1(new_n947), .A2(KEYINPUT62), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(KEYINPUT62), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n894), .A2(new_n712), .A3(new_n936), .ZN(new_n950));
  OAI211_X1 g749(.A(new_n948), .B(new_n949), .C1(new_n946), .C2(new_n950), .ZN(G1353gat));
  NAND3_X1  g750(.A1(new_n894), .A2(new_n711), .A3(new_n936), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(G211gat), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n953), .A2(KEYINPUT126), .A3(KEYINPUT63), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n942), .A2(new_n384), .A3(new_n711), .ZN(new_n955));
  NAND2_X1  g754(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n956));
  OR2_X1    g755(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n952), .A2(G211gat), .A3(new_n956), .A4(new_n957), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n954), .A2(new_n955), .A3(new_n958), .ZN(G1354gat));
  NAND3_X1  g758(.A1(new_n942), .A2(new_n385), .A3(new_n325), .ZN(new_n960));
  AND3_X1   g759(.A1(new_n894), .A2(new_n325), .A3(new_n936), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n960), .B1(new_n961), .B2(new_n385), .ZN(G1355gat));
endmodule


