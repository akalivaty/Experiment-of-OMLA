//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 0 1 1 1 0 1 0 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n784, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009;
  INV_X1    g000(.A(KEYINPUT30), .ZN(new_n202));
  INV_X1    g001(.A(G226gat), .ZN(new_n203));
  INV_X1    g002(.A(G233gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  AND2_X1   g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT24), .ZN(new_n208));
  AOI22_X1  g007(.A1(new_n207), .A2(new_n208), .B1(G169gat), .B2(G176gat), .ZN(new_n209));
  OR2_X1    g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n210), .A2(KEYINPUT24), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT23), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n213), .B1(G169gat), .B2(G176gat), .ZN(new_n214));
  AND3_X1   g013(.A1(new_n209), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT65), .ZN(new_n216));
  INV_X1    g015(.A(G169gat), .ZN(new_n217));
  INV_X1    g016(.A(G176gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(KEYINPUT23), .A3(new_n220), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n221), .A2(KEYINPUT25), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n215), .A2(new_n222), .A3(KEYINPUT66), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n209), .A2(new_n212), .A3(new_n214), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n221), .A2(KEYINPUT25), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT23), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n215), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n231));
  AOI22_X1  g030(.A1(new_n223), .A2(new_n227), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT68), .ZN(new_n234));
  OR3_X1    g033(.A1(new_n233), .A2(new_n228), .A3(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n234), .B1(new_n233), .B2(new_n228), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n220), .ZN(new_n237));
  OAI211_X1 g036(.A(new_n235), .B(new_n236), .C1(new_n237), .C2(KEYINPUT26), .ZN(new_n238));
  XNOR2_X1  g037(.A(KEYINPUT27), .B(G183gat), .ZN(new_n239));
  INV_X1    g038(.A(G190gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT28), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT67), .ZN(new_n243));
  OR2_X1    g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n207), .B1(new_n241), .B2(new_n243), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n238), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n232), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n206), .B1(new_n248), .B2(KEYINPUT29), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n205), .B1(new_n232), .B2(new_n247), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(KEYINPUT75), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT75), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n252), .B(new_n205), .C1(new_n232), .C2(new_n247), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n249), .A2(new_n251), .A3(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G211gat), .B(G218gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT74), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT72), .B(KEYINPUT22), .ZN(new_n258));
  INV_X1    g057(.A(G211gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT73), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT73), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(G211gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n258), .B1(G218gat), .B2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G197gat), .B(G204gat), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n265), .B1(new_n255), .B2(KEYINPUT74), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n257), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  AND2_X1   g066(.A1(KEYINPUT72), .A2(KEYINPUT22), .ZN(new_n268));
  NOR2_X1   g067(.A1(KEYINPUT72), .A2(KEYINPUT22), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(KEYINPUT73), .B(G211gat), .ZN(new_n271));
  INV_X1    g070(.A(G218gat), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT74), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n259), .A2(G218gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n272), .A2(G211gat), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n273), .A2(new_n256), .A3(new_n277), .A4(new_n265), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n267), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n254), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT76), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n223), .A2(new_n227), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n230), .A2(new_n231), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT29), .B1(new_n284), .B2(new_n246), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n281), .B1(new_n285), .B2(new_n205), .ZN(new_n286));
  INV_X1    g085(.A(new_n279), .ZN(new_n287));
  OAI211_X1 g086(.A(KEYINPUT76), .B(new_n206), .C1(new_n248), .C2(KEYINPUT29), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n286), .A2(new_n287), .A3(new_n288), .A4(new_n250), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n280), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G8gat), .B(G36gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(G64gat), .B(G92gat), .ZN(new_n292));
  XOR2_X1   g091(.A(new_n291), .B(new_n292), .Z(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n202), .B1(new_n290), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n295), .B1(new_n294), .B2(new_n290), .ZN(new_n296));
  INV_X1    g095(.A(new_n290), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n297), .A2(new_n202), .A3(new_n293), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(G225gat), .A2(G233gat), .ZN(new_n300));
  INV_X1    g099(.A(G120gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT69), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT69), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G120gat), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n302), .A2(new_n304), .A3(G113gat), .ZN(new_n305));
  INV_X1    g104(.A(G113gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G120gat), .ZN(new_n307));
  AND3_X1   g106(.A1(new_n305), .A2(KEYINPUT70), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT70), .B1(new_n305), .B2(new_n307), .ZN(new_n309));
  XNOR2_X1  g108(.A(G127gat), .B(G134gat), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT1), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NOR3_X1   g111(.A1(new_n308), .A2(new_n309), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n301), .A2(G113gat), .ZN(new_n314));
  AOI21_X1  g113(.A(KEYINPUT1), .B1(new_n307), .B2(new_n314), .ZN(new_n315));
  OR2_X1    g114(.A1(new_n315), .A2(new_n310), .ZN(new_n316));
  NAND2_X1  g115(.A1(G155gat), .A2(G162gat), .ZN(new_n317));
  INV_X1    g116(.A(G155gat), .ZN(new_n318));
  INV_X1    g117(.A(G162gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G141gat), .B(G148gat), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n317), .B(new_n320), .C1(new_n321), .C2(KEYINPUT2), .ZN(new_n322));
  INV_X1    g121(.A(G141gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G148gat), .ZN(new_n324));
  INV_X1    g123(.A(G148gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G141gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n320), .A2(new_n317), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n317), .A2(KEYINPUT2), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n316), .A2(new_n322), .A3(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n313), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n332), .A2(KEYINPUT4), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT77), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n334), .B1(new_n313), .B2(new_n331), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n305), .A2(new_n307), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT70), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n305), .A2(KEYINPUT70), .A3(new_n307), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n338), .A2(new_n311), .A3(new_n339), .A4(new_n310), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n322), .A2(new_n330), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n340), .A2(KEYINPUT77), .A3(new_n342), .A4(new_n316), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n335), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n333), .B1(new_n344), .B2(KEYINPUT4), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n340), .A2(new_n316), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT3), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n322), .A2(new_n347), .A3(new_n330), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n341), .A2(KEYINPUT3), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n346), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n300), .B1(new_n345), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT39), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  XOR2_X1   g152(.A(KEYINPUT79), .B(KEYINPUT0), .Z(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(KEYINPUT80), .ZN(new_n355));
  XNOR2_X1  g154(.A(G1gat), .B(G29gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n355), .B(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G57gat), .B(G85gat), .ZN(new_n358));
  XOR2_X1   g157(.A(new_n357), .B(new_n358), .Z(new_n359));
  NOR2_X1   g158(.A1(new_n315), .A2(new_n310), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n341), .B1(new_n313), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n335), .A2(new_n361), .A3(new_n343), .ZN(new_n362));
  INV_X1    g161(.A(new_n300), .ZN(new_n363));
  OAI21_X1  g162(.A(KEYINPUT39), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n353), .B(new_n359), .C1(new_n351), .C2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT40), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT84), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT84), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n365), .A2(new_n369), .A3(new_n366), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n365), .A2(new_n366), .ZN(new_n372));
  AND2_X1   g171(.A1(new_n350), .A2(new_n300), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n332), .A2(KEYINPUT4), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n373), .B(new_n374), .C1(new_n344), .C2(KEYINPUT4), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT78), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n362), .A2(new_n363), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n376), .B1(new_n377), .B2(KEYINPUT5), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT5), .ZN(new_n379));
  AOI211_X1 g178(.A(KEYINPUT78), .B(new_n379), .C1(new_n362), .C2(new_n363), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n375), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n345), .A2(new_n379), .A3(new_n373), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n359), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n372), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n299), .A2(new_n371), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT29), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n267), .A2(new_n386), .A3(new_n278), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n347), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(new_n341), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n348), .A2(new_n386), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT82), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n348), .A2(KEYINPUT82), .A3(new_n386), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(new_n279), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G228gat), .A2(G233gat), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n389), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(G78gat), .B(G106gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(KEYINPUT31), .B(G50gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT83), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n342), .B1(new_n387), .B2(new_n347), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n267), .A2(new_n278), .B1(new_n348), .B2(new_n386), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n395), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n397), .A2(new_n401), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(G22gat), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n400), .A2(KEYINPUT83), .ZN(new_n407));
  INV_X1    g206(.A(G22gat), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n397), .A2(new_n404), .A3(new_n408), .A4(new_n401), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n406), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n407), .B1(new_n406), .B2(new_n409), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(KEYINPUT85), .B(KEYINPUT38), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT37), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n294), .B1(new_n297), .B2(new_n414), .ZN(new_n415));
  OR2_X1    g214(.A1(new_n415), .A2(KEYINPUT87), .ZN(new_n416));
  XOR2_X1   g215(.A(KEYINPUT86), .B(KEYINPUT37), .Z(new_n417));
  NOR2_X1   g216(.A1(new_n290), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n418), .B1(new_n415), .B2(KEYINPUT87), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n413), .B1(new_n416), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n418), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n294), .A2(new_n413), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n414), .B1(new_n254), .B2(new_n287), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n286), .A2(new_n279), .A3(new_n288), .A4(new_n250), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AOI22_X1  g224(.A1(new_n421), .A2(new_n425), .B1(new_n293), .B2(new_n297), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n383), .A2(KEYINPUT6), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n381), .A2(new_n382), .ZN(new_n428));
  INV_X1    g227(.A(new_n359), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT6), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n381), .A2(new_n359), .A3(new_n382), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n426), .A2(new_n427), .A3(new_n433), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n385), .B(new_n412), .C1(new_n420), .C2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT34), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n284), .A2(new_n346), .A3(new_n246), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n313), .A2(new_n360), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n438), .B1(new_n232), .B2(new_n247), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(G227gat), .A2(G233gat), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n436), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n440), .A2(new_n436), .A3(new_n441), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n442), .B1(KEYINPUT71), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n441), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n437), .A2(new_n439), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT32), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT33), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XOR2_X1   g248(.A(G15gat), .B(G43gat), .Z(new_n450));
  XNOR2_X1  g249(.A(G71gat), .B(G99gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n447), .A2(new_n449), .A3(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n452), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n446), .B(KEYINPUT32), .C1(new_n448), .C2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT71), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n440), .A2(new_n456), .A3(new_n436), .A4(new_n441), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n444), .A2(new_n453), .A3(new_n455), .A4(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n453), .A2(new_n455), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n443), .A2(KEYINPUT71), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n440), .A2(new_n441), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT34), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(new_n457), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  AND3_X1   g263(.A1(new_n458), .A2(new_n464), .A3(KEYINPUT36), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT36), .B1(new_n458), .B2(new_n464), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT81), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n431), .B(new_n432), .C1(new_n383), .C2(new_n468), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n383), .A2(new_n468), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n427), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n296), .A2(new_n298), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n412), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n467), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n435), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n458), .A2(new_n464), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n471), .A2(new_n472), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT35), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT88), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT35), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n412), .A2(new_n482), .A3(new_n458), .A4(new_n464), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n483), .B1(new_n427), .B2(new_n433), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n481), .B1(new_n484), .B2(new_n472), .ZN(new_n485));
  INV_X1    g284(.A(new_n483), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n433), .A2(new_n427), .ZN(new_n487));
  AND4_X1   g286(.A1(new_n481), .A2(new_n486), .A3(new_n487), .A4(new_n472), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n480), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n476), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(G71gat), .ZN(new_n491));
  INV_X1    g290(.A(G78gat), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g292(.A1(G71gat), .A2(G78gat), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n493), .B1(KEYINPUT9), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(G57gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(G64gat), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  OR2_X1    g297(.A1(KEYINPUT95), .A2(G64gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(KEYINPUT95), .A2(G64gat), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n496), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT96), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n498), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(KEYINPUT95), .B(G64gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(G57gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT96), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n495), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  XOR2_X1   g306(.A(G57gat), .B(G64gat), .Z(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT9), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n493), .A2(new_n494), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n513), .A2(KEYINPUT21), .ZN(new_n514));
  XNOR2_X1  g313(.A(G127gat), .B(G155gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n514), .B(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT94), .ZN(new_n517));
  INV_X1    g316(.A(G8gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n408), .A2(G15gat), .ZN(new_n519));
  INV_X1    g318(.A(G15gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(G22gat), .ZN(new_n521));
  AND3_X1   g320(.A1(new_n519), .A2(new_n521), .A3(KEYINPUT93), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT93), .B1(new_n519), .B2(new_n521), .ZN(new_n523));
  INV_X1    g322(.A(G1gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT16), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NOR3_X1   g325(.A1(new_n522), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT93), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n520), .A2(G22gat), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n408), .A2(G15gat), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n519), .A2(new_n521), .A3(KEYINPUT93), .ZN(new_n532));
  AOI21_X1  g331(.A(G1gat), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n517), .B(new_n518), .C1(new_n527), .C2(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n524), .B1(new_n522), .B2(new_n523), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n531), .A2(new_n532), .A3(new_n525), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n517), .A2(new_n518), .ZN(new_n537));
  NAND2_X1  g336(.A1(KEYINPUT94), .A2(G8gat), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n535), .A2(new_n536), .A3(new_n537), .A4(new_n538), .ZN(new_n539));
  AOI22_X1  g338(.A1(new_n513), .A2(KEYINPUT21), .B1(new_n534), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n516), .B(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G231gat), .A2(G233gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(KEYINPUT97), .ZN(new_n543));
  XOR2_X1   g342(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G183gat), .B(G211gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n541), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n541), .A2(new_n547), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(G43gat), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT15), .B1(new_n551), .B2(G50gat), .ZN(new_n552));
  INV_X1    g351(.A(G50gat), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n553), .A2(G43gat), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(G29gat), .A2(G36gat), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT89), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(KEYINPUT89), .A2(G29gat), .A3(G36gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT91), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n562), .B1(new_n551), .B2(G50gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n551), .A2(G50gat), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n553), .A2(KEYINPUT91), .A3(G43gat), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT90), .B(KEYINPUT15), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(G29gat), .ZN(new_n569));
  INV_X1    g368(.A(G36gat), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n569), .A2(new_n570), .A3(KEYINPUT14), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT14), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n572), .B1(G29gat), .B2(G36gat), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n571), .A2(new_n573), .A3(KEYINPUT92), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n571), .A2(new_n573), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT92), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n561), .A2(new_n568), .A3(new_n574), .A4(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT17), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n555), .B1(new_n575), .B2(new_n560), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n579), .B1(new_n578), .B2(new_n580), .ZN(new_n583));
  NAND2_X1  g382(.A1(G85gat), .A2(G92gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(KEYINPUT7), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT7), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n586), .A2(G85gat), .A3(G92gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT99), .ZN(new_n589));
  INV_X1    g388(.A(G92gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(G85gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(KEYINPUT99), .A2(G92gat), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G99gat), .A2(G106gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT8), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n588), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n595), .ZN(new_n598));
  NOR2_X1   g397(.A1(G99gat), .A2(G106gat), .ZN(new_n599));
  OAI21_X1  g398(.A(KEYINPUT100), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(G99gat), .ZN(new_n601));
  INV_X1    g400(.A(G106gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT100), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n603), .A2(new_n604), .A3(new_n595), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n597), .A2(new_n606), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n597), .A2(new_n606), .ZN(new_n608));
  OAI22_X1  g407(.A1(new_n582), .A2(new_n583), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n607), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n578), .A2(new_n580), .ZN(new_n611));
  AND2_X1   g410(.A1(G232gat), .A2(G233gat), .ZN(new_n612));
  AOI22_X1  g411(.A1(new_n610), .A2(new_n611), .B1(KEYINPUT41), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT101), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n613), .A2(new_n614), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n609), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n612), .A2(KEYINPUT41), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT98), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n619), .ZN(new_n621));
  OAI211_X1 g420(.A(new_n609), .B(new_n621), .C1(new_n615), .C2(new_n616), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(G190gat), .B(G218gat), .Z(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT102), .ZN(new_n625));
  XNOR2_X1  g424(.A(G134gat), .B(G162gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n620), .A2(new_n622), .A3(new_n627), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OAI22_X1  g430(.A1(new_n507), .A2(new_n512), .B1(new_n608), .B2(new_n607), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT10), .ZN(new_n633));
  INV_X1    g432(.A(new_n495), .ZN(new_n634));
  AND2_X1   g433(.A1(KEYINPUT95), .A2(G64gat), .ZN(new_n635));
  NOR2_X1   g434(.A1(KEYINPUT95), .A2(G64gat), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n502), .B(G57gat), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n497), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n502), .B1(new_n504), .B2(G57gat), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n634), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n595), .A2(KEYINPUT8), .ZN(new_n641));
  AND2_X1   g440(.A1(KEYINPUT99), .A2(G92gat), .ZN(new_n642));
  NOR2_X1   g441(.A1(KEYINPUT99), .A2(G92gat), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n641), .B1(new_n644), .B2(new_n592), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n645), .A2(new_n600), .A3(new_n605), .A4(new_n588), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n597), .A2(new_n606), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n640), .A2(new_n646), .A3(new_n511), .A4(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n632), .A2(new_n633), .A3(new_n648), .ZN(new_n649));
  AND4_X1   g448(.A1(new_n640), .A2(new_n646), .A3(new_n511), .A4(new_n647), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(KEYINPUT10), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(G230gat), .A2(G233gat), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G120gat), .B(G148gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(G176gat), .B(G204gat), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n655), .B(new_n656), .Z(new_n657));
  AND2_X1   g456(.A1(new_n632), .A2(new_n648), .ZN(new_n658));
  OAI211_X1 g457(.A(new_n654), .B(new_n657), .C1(new_n658), .C2(new_n653), .ZN(new_n659));
  INV_X1    g458(.A(new_n657), .ZN(new_n660));
  INV_X1    g459(.A(new_n653), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n661), .B1(new_n649), .B2(new_n651), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n653), .B1(new_n632), .B2(new_n648), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n660), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n659), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n550), .A2(new_n631), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(G113gat), .B(G141gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(G197gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT11), .B(G169gat), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n669), .B(new_n670), .Z(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT12), .ZN(new_n672));
  NAND2_X1  g471(.A1(G229gat), .A2(G233gat), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n673), .B(KEYINPUT13), .Z(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n534), .A2(new_n539), .ZN(new_n676));
  INV_X1    g475(.A(new_n611), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n534), .A2(new_n611), .A3(new_n539), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n675), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n676), .B1(new_n582), .B2(new_n583), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n681), .A2(new_n673), .A3(new_n679), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT18), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n680), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n681), .A2(KEYINPUT18), .A3(new_n673), .A4(new_n679), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n672), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n684), .A2(new_n672), .A3(new_n685), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n667), .A2(new_n690), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n490), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n471), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(G1gat), .ZN(G1324gat));
  INV_X1    g494(.A(new_n692), .ZN(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT16), .B(G8gat), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n696), .A2(new_n472), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n518), .B1(new_n692), .B2(new_n299), .ZN(new_n699));
  OAI21_X1  g498(.A(KEYINPUT42), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n700), .B1(KEYINPUT42), .B2(new_n698), .ZN(G1325gat));
  INV_X1    g500(.A(new_n467), .ZN(new_n702));
  OAI21_X1  g501(.A(G15gat), .B1(new_n696), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n477), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n692), .A2(new_n520), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(G1326gat));
  NAND2_X1  g505(.A1(new_n692), .A2(new_n474), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT103), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT43), .B(G22gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1327gat));
  AOI21_X1  g509(.A(new_n631), .B1(new_n476), .B2(new_n489), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n550), .A2(new_n690), .A3(new_n665), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n713), .A2(G29gat), .A3(new_n471), .ZN(new_n714));
  XOR2_X1   g513(.A(new_n714), .B(KEYINPUT45), .Z(new_n715));
  NAND2_X1  g514(.A1(new_n489), .A2(KEYINPUT104), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n486), .A2(new_n472), .A3(new_n487), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(KEYINPUT88), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n484), .A2(new_n481), .A3(new_n472), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT104), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n720), .A2(new_n721), .A3(new_n480), .ZN(new_n722));
  AOI22_X1  g521(.A1(new_n716), .A2(new_n722), .B1(new_n435), .B2(new_n475), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n631), .A2(KEYINPUT44), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n726));
  OAI22_X1  g525(.A1(new_n723), .A2(new_n725), .B1(new_n711), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(new_n712), .ZN(new_n728));
  OAI21_X1  g527(.A(G29gat), .B1(new_n728), .B2(new_n471), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n715), .A2(new_n729), .ZN(G1328gat));
  NOR3_X1   g529(.A1(new_n713), .A2(G36gat), .A3(new_n472), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT46), .ZN(new_n732));
  OAI21_X1  g531(.A(G36gat), .B1(new_n728), .B2(new_n472), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(G1329gat));
  OAI21_X1  g533(.A(new_n551), .B1(new_n713), .B2(new_n477), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n467), .A2(G43gat), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n735), .B1(new_n728), .B2(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g537(.A1(new_n716), .A2(new_n722), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n725), .B1(new_n739), .B2(new_n476), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n711), .A2(new_n726), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n474), .B(new_n712), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT105), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n727), .A2(KEYINPUT105), .A3(new_n474), .A4(new_n712), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n744), .A2(G50gat), .A3(new_n745), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n711), .A2(new_n553), .A3(new_n474), .A4(new_n712), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(KEYINPUT48), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n742), .A2(G50gat), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n747), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT48), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n750), .A2(new_n754), .A3(KEYINPUT106), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT106), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n553), .B1(new_n742), .B2(new_n743), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n748), .B1(new_n757), .B2(new_n745), .ZN(new_n758));
  AOI21_X1  g557(.A(KEYINPUT48), .B1(new_n751), .B2(new_n747), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n756), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n755), .A2(new_n760), .ZN(G1331gat));
  NOR2_X1   g560(.A1(new_n489), .A2(KEYINPUT104), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n721), .B1(new_n720), .B2(new_n480), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n476), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(new_n550), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n629), .A2(new_n630), .ZN(new_n766));
  NOR4_X1   g565(.A1(new_n765), .A2(new_n689), .A3(new_n766), .A4(new_n666), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n768), .A2(new_n471), .ZN(new_n769));
  XOR2_X1   g568(.A(KEYINPUT107), .B(G57gat), .Z(new_n770));
  XNOR2_X1  g569(.A(new_n769), .B(new_n770), .ZN(G1332gat));
  NOR2_X1   g570(.A1(new_n768), .A2(new_n472), .ZN(new_n772));
  NOR2_X1   g571(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n773));
  AND2_X1   g572(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n772), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n775), .B1(new_n772), .B2(new_n773), .ZN(G1333gat));
  INV_X1    g575(.A(KEYINPUT108), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n768), .A2(new_n777), .A3(new_n477), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n768), .B2(new_n477), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n491), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n467), .A2(G71gat), .ZN(new_n781));
  OAI22_X1  g580(.A1(new_n778), .A2(new_n780), .B1(new_n768), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g582(.A1(new_n768), .A2(new_n412), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(new_n492), .ZN(G1335gat));
  AND2_X1   g584(.A1(KEYINPUT109), .A2(KEYINPUT51), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n765), .A2(new_n690), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(new_n631), .ZN(new_n789));
  AND3_X1   g588(.A1(new_n764), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n787), .B1(new_n764), .B2(new_n789), .ZN(new_n791));
  OAI22_X1  g590(.A1(new_n790), .A2(new_n791), .B1(KEYINPUT109), .B2(KEYINPUT51), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n665), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n693), .A2(new_n592), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n740), .A2(new_n741), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n788), .A2(new_n666), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n795), .A2(new_n471), .A3(new_n797), .ZN(new_n798));
  OAI22_X1  g597(.A1(new_n793), .A2(new_n794), .B1(new_n592), .B2(new_n798), .ZN(G1336gat));
  NAND4_X1  g598(.A1(new_n792), .A2(new_n590), .A3(new_n299), .A4(new_n665), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n727), .A2(new_n299), .A3(new_n796), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n801), .B1(new_n643), .B2(new_n642), .ZN(new_n802));
  XNOR2_X1  g601(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n800), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n803), .B1(new_n800), .B2(new_n802), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n804), .A2(new_n805), .ZN(G1337gat));
  INV_X1    g605(.A(KEYINPUT111), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n477), .A2(G99gat), .ZN(new_n808));
  AND3_X1   g607(.A1(new_n792), .A2(new_n665), .A3(new_n808), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n795), .A2(new_n702), .A3(new_n797), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n810), .A2(new_n601), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n807), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(new_n808), .ZN(new_n813));
  OAI221_X1 g612(.A(KEYINPUT111), .B1(new_n601), .B2(new_n810), .C1(new_n793), .C2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(G1338gat));
  NOR2_X1   g614(.A1(new_n412), .A2(G106gat), .ZN(new_n816));
  AND3_X1   g615(.A1(new_n792), .A2(new_n665), .A3(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n795), .A2(new_n412), .A3(new_n797), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n818), .A2(new_n602), .ZN(new_n819));
  OAI21_X1  g618(.A(KEYINPUT53), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n821));
  INV_X1    g620(.A(new_n816), .ZN(new_n822));
  OAI221_X1 g621(.A(new_n821), .B1(new_n602), .B2(new_n818), .C1(new_n793), .C2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n820), .A2(new_n823), .ZN(G1339gat));
  NOR2_X1   g623(.A1(new_n667), .A2(new_n689), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n652), .A2(new_n827), .A3(new_n653), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n632), .A2(new_n633), .A3(new_n648), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n661), .B1(new_n648), .B2(new_n633), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT54), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n828), .B(new_n660), .C1(new_n831), .C2(new_n662), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT55), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n662), .A2(new_n663), .A3(new_n660), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n653), .B1(new_n650), .B2(KEYINPUT10), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n827), .B1(new_n836), .B2(new_n649), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n833), .B1(new_n654), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n657), .B1(new_n662), .B2(new_n827), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n835), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n629), .A2(new_n630), .A3(new_n834), .A4(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n678), .A2(new_n679), .A3(new_n675), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n673), .B1(new_n681), .B2(new_n679), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n671), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT112), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n673), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n611), .A2(KEYINPUT17), .ZN(new_n849));
  AOI22_X1  g648(.A1(new_n849), .A2(new_n581), .B1(new_n534), .B2(new_n539), .ZN(new_n850));
  INV_X1    g649(.A(new_n679), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n848), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n842), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n853), .A2(KEYINPUT112), .A3(new_n671), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n847), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n688), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n682), .A2(new_n683), .ZN(new_n858));
  INV_X1    g657(.A(new_n680), .ZN(new_n859));
  AND4_X1   g658(.A1(new_n672), .A2(new_n858), .A3(new_n685), .A4(new_n859), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n840), .B(new_n834), .C1(new_n860), .C2(new_n686), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT112), .B1(new_n853), .B2(new_n671), .ZN(new_n862));
  INV_X1    g661(.A(new_n671), .ZN(new_n863));
  AOI211_X1 g662(.A(new_n846), .B(new_n863), .C1(new_n852), .C2(new_n842), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n688), .B(new_n665), .C1(new_n862), .C2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT113), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n766), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n861), .A2(KEYINPUT113), .A3(new_n865), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n857), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n826), .B1(new_n870), .B2(new_n550), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n871), .A2(new_n478), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n693), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT114), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n873), .B(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n472), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT115), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n876), .B(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n878), .A2(new_n306), .A3(new_n689), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n872), .A2(new_n693), .A3(new_n472), .ZN(new_n880));
  OAI21_X1  g679(.A(G113gat), .B1(new_n880), .B2(new_n690), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(new_n881), .ZN(G1340gat));
  NAND4_X1  g681(.A1(new_n878), .A2(new_n302), .A3(new_n304), .A4(new_n665), .ZN(new_n883));
  OAI21_X1  g682(.A(G120gat), .B1(new_n880), .B2(new_n666), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(G1341gat));
  OAI21_X1  g684(.A(G127gat), .B1(new_n880), .B2(new_n765), .ZN(new_n886));
  OR2_X1    g685(.A1(new_n765), .A2(G127gat), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n886), .B1(new_n876), .B2(new_n887), .ZN(G1342gat));
  INV_X1    g687(.A(G134gat), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n299), .A2(new_n631), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n875), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n891), .A2(KEYINPUT56), .ZN(new_n892));
  INV_X1    g691(.A(new_n890), .ZN(new_n893));
  OAI21_X1  g692(.A(G134gat), .B1(new_n873), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n891), .A2(KEYINPUT56), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n892), .A2(new_n894), .A3(new_n895), .ZN(G1343gat));
  NOR3_X1   g695(.A1(new_n299), .A2(new_n467), .A3(new_n471), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n871), .A2(new_n897), .A3(new_n474), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n898), .A2(G141gat), .A3(new_n690), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n899), .A2(KEYINPUT58), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT118), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n865), .A2(new_n901), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n855), .A2(KEYINPUT118), .A3(new_n688), .A4(new_n665), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n902), .A2(new_n861), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n631), .ZN(new_n905));
  INV_X1    g704(.A(new_n857), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n550), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI211_X1 g706(.A(KEYINPUT57), .B(new_n474), .C1(new_n907), .C2(new_n825), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT119), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n857), .B1(new_n904), .B2(new_n631), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n826), .B1(new_n911), .B2(new_n550), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n912), .A2(KEYINPUT119), .A3(KEYINPUT57), .A4(new_n474), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT117), .ZN(new_n915));
  XNOR2_X1  g714(.A(KEYINPUT116), .B(KEYINPUT57), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  AOI211_X1 g716(.A(new_n915), .B(new_n917), .C1(new_n871), .C2(new_n474), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n866), .A2(new_n867), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n631), .A3(new_n869), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n550), .B1(new_n920), .B2(new_n906), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n474), .B1(new_n921), .B2(new_n825), .ZN(new_n922));
  AOI21_X1  g721(.A(KEYINPUT117), .B1(new_n922), .B2(new_n916), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n914), .A2(new_n918), .A3(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(new_n897), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n924), .A2(new_n690), .A3(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n900), .B1(new_n926), .B2(new_n323), .ZN(new_n927));
  OAI21_X1  g726(.A(KEYINPUT120), .B1(new_n924), .B2(new_n925), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT120), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n922), .A2(new_n916), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(new_n915), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n922), .A2(KEYINPUT117), .A3(new_n916), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n929), .B(new_n897), .C1(new_n933), .C2(new_n914), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n928), .A2(new_n689), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n899), .B1(new_n935), .B2(G141gat), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT58), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n927), .B1(new_n936), .B2(new_n937), .ZN(G1344gat));
  AND2_X1   g737(.A1(new_n912), .A2(new_n474), .ZN(new_n939));
  OAI22_X1  g738(.A1(new_n939), .A2(KEYINPUT57), .B1(new_n922), .B2(new_n916), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n940), .A2(new_n665), .A3(new_n897), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n941), .A2(KEYINPUT122), .ZN(new_n942));
  OAI21_X1  g741(.A(G148gat), .B1(new_n941), .B2(KEYINPUT122), .ZN(new_n943));
  OAI21_X1  g742(.A(KEYINPUT59), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n928), .A2(new_n665), .A3(new_n934), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT121), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n325), .A2(KEYINPUT59), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n946), .B1(new_n945), .B2(new_n947), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n944), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(new_n898), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n951), .A2(new_n325), .A3(new_n665), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(G1345gat));
  OAI21_X1  g752(.A(new_n318), .B1(new_n898), .B2(new_n765), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n928), .A2(new_n934), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n550), .A2(G155gat), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT123), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n957), .B(new_n958), .ZN(G1346gat));
  OAI21_X1  g758(.A(G162gat), .B1(new_n955), .B2(new_n631), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n951), .A2(new_n319), .A3(new_n766), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(G1347gat));
  NOR2_X1   g761(.A1(new_n693), .A2(new_n472), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n872), .A2(new_n963), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n964), .A2(new_n217), .A3(new_n690), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n871), .A2(new_n471), .ZN(new_n966));
  NOR3_X1   g765(.A1(new_n472), .A2(new_n474), .A3(new_n477), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(new_n689), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n965), .B1(new_n217), .B2(new_n970), .ZN(G1348gat));
  OAI21_X1  g770(.A(G176gat), .B1(new_n964), .B2(new_n666), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n665), .A2(new_n218), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n972), .B1(new_n968), .B2(new_n973), .ZN(G1349gat));
  OAI21_X1  g773(.A(G183gat), .B1(new_n964), .B2(new_n765), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n550), .A2(new_n239), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n975), .B1(new_n968), .B2(new_n976), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT60), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n978), .A2(KEYINPUT124), .ZN(new_n979));
  XNOR2_X1  g778(.A(new_n977), .B(new_n979), .ZN(G1350gat));
  NAND3_X1  g779(.A1(new_n969), .A2(new_n240), .A3(new_n766), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n872), .A2(new_n766), .A3(new_n963), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT61), .ZN(new_n983));
  AND3_X1   g782(.A1(new_n982), .A2(new_n983), .A3(G190gat), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n983), .B1(new_n982), .B2(G190gat), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n981), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  XOR2_X1   g785(.A(new_n986), .B(KEYINPUT125), .Z(G1351gat));
  NOR3_X1   g786(.A1(new_n467), .A2(new_n412), .A3(new_n472), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n966), .A2(new_n988), .ZN(new_n989));
  NOR3_X1   g788(.A1(new_n989), .A2(G197gat), .A3(new_n690), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n963), .A2(new_n702), .ZN(new_n991));
  XNOR2_X1  g790(.A(new_n991), .B(KEYINPUT126), .ZN(new_n992));
  AND2_X1   g791(.A1(new_n940), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n993), .A2(new_n689), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n990), .B1(new_n994), .B2(G197gat), .ZN(new_n995));
  XOR2_X1   g794(.A(new_n995), .B(KEYINPUT127), .Z(G1352gat));
  NOR3_X1   g795(.A1(new_n989), .A2(G204gat), .A3(new_n666), .ZN(new_n997));
  XNOR2_X1  g796(.A(new_n997), .B(KEYINPUT62), .ZN(new_n998));
  AND2_X1   g797(.A1(new_n993), .A2(new_n665), .ZN(new_n999));
  INV_X1    g798(.A(G204gat), .ZN(new_n1000));
  OAI21_X1  g799(.A(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(G1353gat));
  NOR2_X1   g800(.A1(new_n991), .A2(new_n765), .ZN(new_n1002));
  AOI21_X1  g801(.A(new_n259), .B1(new_n940), .B2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g802(.A(new_n1003), .B(KEYINPUT63), .ZN(new_n1004));
  INV_X1    g803(.A(new_n989), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n1005), .A2(new_n271), .A3(new_n550), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1004), .A2(new_n1006), .ZN(G1354gat));
  NAND3_X1  g806(.A1(new_n1005), .A2(new_n272), .A3(new_n766), .ZN(new_n1008));
  AND2_X1   g807(.A1(new_n993), .A2(new_n766), .ZN(new_n1009));
  OAI21_X1  g808(.A(new_n1008), .B1(new_n1009), .B2(new_n272), .ZN(G1355gat));
endmodule


