//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 1 0 0 1 0 0 1 0 1 0 1 1 1 1 1 0 1 0 0 1 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 0 1 0 0 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n563, new_n564, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n620, new_n622, new_n623, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1206, new_n1208;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT66), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT67), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT68), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT69), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G567), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  INV_X1    g031(.A(new_n451), .ZN(new_n457));
  AOI21_X1  g032(.A(new_n456), .B1(new_n457), .B2(G2106), .ZN(G319));
  OR2_X1    g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G137), .ZN(new_n462));
  NAND2_X1  g037(.A1(G101), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(G2105), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(G125), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT70), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n469), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n464), .B1(new_n472), .B2(new_n473), .ZN(G160));
  NOR2_X1   g049(.A1(new_n465), .A2(new_n466), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n475), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n476), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n478), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  INV_X1    g059(.A(KEYINPUT71), .ZN(new_n485));
  AND2_X1   g060(.A1(G126), .A2(G2105), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n461), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n486), .B1(new_n465), .B2(new_n466), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(KEYINPUT71), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n461), .A2(G138), .A3(new_n476), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G114), .C2(new_n476), .ZN(new_n495));
  AND2_X1   g070(.A1(KEYINPUT4), .A2(G138), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n476), .B(new_n496), .C1(new_n465), .C2(new_n466), .ZN(new_n497));
  AND2_X1   g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n490), .A2(new_n493), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  OR2_X1    g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n503), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  OR2_X1    g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT72), .B1(new_n507), .B2(G651), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(new_n505), .A3(KEYINPUT6), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(G50), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT73), .B(KEYINPUT6), .ZN(new_n514));
  AOI21_X1  g089(.A(KEYINPUT74), .B1(new_n514), .B2(G651), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT73), .A2(KEYINPUT6), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT73), .A2(KEYINPUT6), .ZN(new_n517));
  OAI211_X1 g092(.A(KEYINPUT74), .B(G651), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  OAI211_X1 g094(.A(new_n511), .B(new_n513), .C1(new_n515), .C2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n508), .A2(new_n510), .B1(new_n501), .B2(new_n502), .ZN(new_n521));
  OAI211_X1 g096(.A(G88), .B(new_n521), .C1(new_n515), .C2(new_n519), .ZN(new_n522));
  AND3_X1   g097(.A1(new_n520), .A2(new_n522), .A3(KEYINPUT75), .ZN(new_n523));
  AOI21_X1  g098(.A(KEYINPUT75), .B1(new_n520), .B2(new_n522), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n506), .B1(new_n523), .B2(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  AND2_X1   g101(.A1(new_n508), .A2(new_n510), .ZN(new_n527));
  OAI21_X1  g102(.A(G651), .B1(new_n516), .B2(new_n517), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT74), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n527), .B1(new_n530), .B2(new_n518), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n531), .A2(G543), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G51), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n503), .A2(G63), .A3(G651), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n530), .A2(new_n518), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(new_n521), .ZN(new_n539));
  INV_X1    g114(.A(G89), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(KEYINPUT76), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n541), .A2(KEYINPUT76), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n535), .A2(new_n542), .A3(new_n543), .ZN(G286));
  INV_X1    g119(.A(G286), .ZN(G168));
  NAND2_X1  g120(.A1(new_n532), .A2(G52), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n503), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(new_n505), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n511), .A2(new_n503), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n549), .B1(new_n530), .B2(new_n518), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G90), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n546), .A2(new_n548), .A3(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  NAND2_X1  g128(.A1(new_n532), .A2(G43), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n503), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n555), .A2(new_n505), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n556), .B1(new_n550), .B2(G81), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT77), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  NAND4_X1  g140(.A1(new_n538), .A2(G53), .A3(G543), .A4(new_n511), .ZN(new_n566));
  OR3_X1    g141(.A1(new_n566), .A2(KEYINPUT79), .A3(KEYINPUT9), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(KEYINPUT9), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT78), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT79), .B1(new_n566), .B2(KEYINPUT9), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT78), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n566), .A2(new_n571), .A3(KEYINPUT9), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n567), .A2(new_n569), .A3(new_n570), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(new_n503), .ZN(new_n575));
  INV_X1    g150(.A(G65), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT80), .ZN(new_n578));
  OR2_X1    g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n505), .B1(new_n577), .B2(new_n578), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n579), .A2(new_n580), .B1(G91), .B2(new_n550), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n573), .A2(new_n581), .ZN(G299));
  INV_X1    g157(.A(G74), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n505), .B1(new_n575), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n584), .B1(new_n550), .B2(G87), .ZN(new_n585));
  AND2_X1   g160(.A1(G49), .A2(G543), .ZN(new_n586));
  AND4_X1   g161(.A1(KEYINPUT81), .A2(new_n538), .A3(new_n511), .A4(new_n586), .ZN(new_n587));
  AOI21_X1  g162(.A(KEYINPUT81), .B1(new_n531), .B2(new_n586), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n585), .B1(new_n587), .B2(new_n588), .ZN(G288));
  NAND4_X1  g164(.A1(new_n538), .A2(G48), .A3(G543), .A4(new_n511), .ZN(new_n590));
  AND2_X1   g165(.A1(G73), .A2(G543), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n591), .B(KEYINPUT82), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n503), .A2(G61), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n505), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n538), .A2(G86), .A3(new_n521), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n590), .A2(new_n595), .A3(new_n596), .ZN(G305));
  NAND2_X1  g172(.A1(new_n532), .A2(G47), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n503), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n599), .A2(new_n505), .ZN(new_n600));
  XNOR2_X1  g175(.A(KEYINPUT83), .B(G85), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n600), .B1(new_n550), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n598), .A2(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n550), .A2(G92), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n605), .B(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(G79), .A2(G543), .ZN(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(KEYINPUT84), .Z(new_n609));
  INV_X1    g184(.A(G66), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(new_n575), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n532), .A2(G54), .B1(G651), .B2(new_n611), .ZN(new_n612));
  AND2_X1   g187(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n604), .B1(new_n613), .B2(G868), .ZN(G284));
  OAI21_X1  g189(.A(new_n604), .B1(new_n613), .B2(G868), .ZN(G321));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  INV_X1    g191(.A(G299), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(G297));
  XNOR2_X1  g193(.A(G297), .B(KEYINPUT85), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n613), .B1(new_n620), .B2(G860), .ZN(G148));
  INV_X1    g196(.A(G868), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n558), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n607), .A2(new_n612), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n624), .A2(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n623), .B1(new_n625), .B2(new_n622), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n479), .A2(G2104), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G2100), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT87), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n479), .A2(G135), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT88), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n477), .A2(G123), .ZN(new_n636));
  NOR2_X1   g211(.A1(G99), .A2(G2105), .ZN(new_n637));
  OAI21_X1  g212(.A(G2104), .B1(new_n476), .B2(G111), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n635), .B(new_n636), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(G2096), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n633), .B(new_n641), .C1(G2100), .C2(new_n631), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT89), .ZN(G156));
  XOR2_X1   g218(.A(G2451), .B(G2454), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2427), .B(G2438), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2430), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT15), .B(G2435), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(new_n654), .A3(KEYINPUT14), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n649), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n649), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(new_n658), .A3(G14), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(G401));
  XOR2_X1   g235(.A(G2072), .B(G2078), .Z(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT17), .Z(new_n662));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  XNOR2_X1  g238(.A(G2067), .B(G2678), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  INV_X1    g241(.A(new_n663), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(new_n661), .ZN(new_n668));
  OAI211_X1 g243(.A(new_n665), .B(new_n666), .C1(new_n664), .C2(new_n668), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n666), .A2(new_n661), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT18), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(new_n640), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n673), .A2(G2100), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(G2100), .ZN(new_n675));
  AND2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(G227));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n680), .A2(KEYINPUT90), .ZN(new_n681));
  XOR2_X1   g256(.A(G1971), .B(G1976), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(KEYINPUT90), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n681), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT20), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n678), .A2(new_n679), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(new_n680), .ZN(new_n688));
  MUX2_X1   g263(.A(new_n688), .B(new_n687), .S(new_n683), .Z(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1991), .B(G1996), .ZN(new_n695));
  INV_X1    g270(.A(G1981), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n694), .B(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(G229));
  INV_X1    g274(.A(G29), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(KEYINPUT24), .B2(G34), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(KEYINPUT24), .B2(G34), .ZN(new_n702));
  INV_X1    g277(.A(G160), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(G29), .ZN(new_n704));
  INV_X1    g279(.A(G2084), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT99), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n700), .A2(G33), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n476), .A2(G103), .A3(G2104), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT25), .ZN(new_n710));
  AOI22_X1  g285(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n711), .A2(new_n476), .ZN(new_n712));
  AOI211_X1 g287(.A(new_n710), .B(new_n712), .C1(G139), .C2(new_n479), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n708), .B1(new_n713), .B2(new_n700), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(G2072), .Z(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT27), .B(G1996), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT101), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n700), .A2(G32), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n479), .A2(G141), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT100), .ZN(new_n720));
  AND3_X1   g295(.A1(new_n476), .A2(G105), .A3(G2104), .ZN(new_n721));
  NAND3_X1  g296(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT26), .ZN(new_n723));
  AOI211_X1 g298(.A(new_n721), .B(new_n723), .C1(G129), .C2(new_n477), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n718), .B1(new_n725), .B2(G29), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n707), .B(new_n715), .C1(new_n717), .C2(new_n727), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT102), .Z(new_n729));
  XOR2_X1   g304(.A(KEYINPUT105), .B(KEYINPUT23), .Z(new_n730));
  INV_X1    g305(.A(G16), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G20), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n730), .B(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(new_n617), .B2(new_n731), .ZN(new_n734));
  INV_X1    g309(.A(G1956), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n731), .A2(G4), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n613), .B2(new_n731), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G1348), .ZN(new_n739));
  NOR2_X1   g314(.A1(G162), .A2(new_n700), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n700), .B2(G35), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT29), .B(G2090), .Z(new_n742));
  NOR2_X1   g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n639), .A2(new_n700), .ZN(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n743), .B1(KEYINPUT104), .B2(new_n745), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n745), .A2(KEYINPUT104), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n700), .A2(G27), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G164), .B2(new_n700), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n749), .A2(G2078), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT30), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n751), .A2(G28), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n700), .B1(new_n751), .B2(G28), .ZN(new_n753));
  AND2_X1   g328(.A1(KEYINPUT31), .A2(G11), .ZN(new_n754));
  NOR2_X1   g329(.A1(KEYINPUT31), .A2(G11), .ZN(new_n755));
  OAI22_X1  g330(.A1(new_n752), .A2(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n741), .B2(new_n742), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n746), .A2(new_n747), .A3(new_n750), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n731), .A2(G19), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n559), .B2(new_n731), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G1341), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n704), .A2(new_n705), .ZN(new_n762));
  NOR4_X1   g337(.A1(new_n739), .A2(new_n758), .A3(new_n761), .A4(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(G171), .A2(new_n731), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G5), .B2(new_n731), .ZN(new_n765));
  INV_X1    g340(.A(G1961), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT97), .B(KEYINPUT28), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT98), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n700), .A2(G26), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n770), .B(new_n771), .Z(new_n772));
  OR2_X1    g347(.A1(G104), .A2(G2105), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n773), .B(G2104), .C1(G116), .C2(new_n476), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT96), .ZN(new_n775));
  AOI22_X1  g350(.A1(G128), .A2(new_n477), .B1(new_n479), .B2(G140), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n772), .B1(G29), .B2(new_n777), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G2067), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n727), .A2(new_n717), .B1(G2078), .B2(new_n749), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n767), .A2(new_n768), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n731), .A2(G21), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G168), .B2(new_n731), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT103), .B(G1966), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  AND2_X1   g360(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n783), .A2(new_n785), .ZN(new_n787));
  NOR3_X1   g362(.A1(new_n781), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n729), .A2(new_n736), .A3(new_n763), .A4(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT36), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n790), .A2(KEYINPUT94), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n700), .A2(G25), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n477), .A2(G119), .ZN(new_n793));
  OR2_X1    g368(.A1(G95), .A2(G2105), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n794), .B(G2104), .C1(G107), .C2(new_n476), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G131), .B2(new_n479), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n792), .B1(new_n797), .B2(new_n700), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT35), .B(G1991), .Z(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT91), .Z(new_n800));
  XNOR2_X1  g375(.A(new_n798), .B(new_n800), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n731), .A2(G24), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G290), .B2(G16), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n803), .A2(G1986), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(G1986), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n801), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT33), .B(G1976), .Z(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT92), .ZN(new_n809));
  NAND2_X1  g384(.A1(G288), .A2(G16), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n731), .A2(G23), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(new_n811), .ZN(new_n813));
  AOI211_X1 g388(.A(KEYINPUT92), .B(new_n813), .C1(G288), .C2(G16), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n808), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  OAI211_X1 g390(.A(G16), .B(new_n506), .C1(new_n523), .C2(new_n524), .ZN(new_n816));
  OR2_X1    g391(.A1(G16), .A2(G22), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n816), .A2(G1971), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n538), .A2(new_n511), .A3(new_n586), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT81), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n531), .A2(KEYINPUT81), .A3(new_n586), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n731), .B1(new_n823), .B2(new_n585), .ZN(new_n824));
  OAI21_X1  g399(.A(KEYINPUT92), .B1(new_n824), .B2(new_n813), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n810), .A2(new_n809), .A3(new_n811), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n825), .A2(new_n807), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n816), .A2(new_n817), .ZN(new_n828));
  INV_X1    g403(.A(G1971), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT32), .B(G1981), .Z(new_n830));
  AOI21_X1  g405(.A(new_n594), .B1(new_n550), .B2(G86), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n731), .B1(new_n831), .B2(new_n590), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n731), .A2(G6), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n830), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n833), .B1(G305), .B2(G16), .ZN(new_n835));
  INV_X1    g410(.A(new_n830), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n828), .A2(new_n829), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n815), .A2(new_n818), .A3(new_n827), .A4(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n806), .B1(new_n839), .B2(KEYINPUT34), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(KEYINPUT93), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT93), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n842), .B(new_n806), .C1(new_n839), .C2(KEYINPUT34), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n839), .A2(KEYINPUT34), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n841), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT95), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT94), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n847), .A2(KEYINPUT36), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n845), .A2(new_n846), .A3(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n846), .B1(new_n845), .B2(new_n849), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n791), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n843), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n828), .A2(new_n829), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n834), .A2(new_n837), .ZN(new_n856));
  AND3_X1   g431(.A1(new_n855), .A2(new_n818), .A3(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT34), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n857), .A2(new_n858), .A3(new_n827), .A4(new_n815), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n842), .B1(new_n859), .B2(new_n806), .ZN(new_n860));
  INV_X1    g435(.A(new_n844), .ZN(new_n861));
  NOR3_X1   g436(.A1(new_n854), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(KEYINPUT95), .B1(new_n862), .B2(new_n848), .ZN(new_n863));
  INV_X1    g438(.A(new_n791), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n863), .A2(new_n864), .A3(new_n850), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n789), .B1(new_n853), .B2(new_n865), .ZN(G311));
  INV_X1    g441(.A(new_n789), .ZN(new_n867));
  NOR3_X1   g442(.A1(new_n851), .A2(new_n852), .A3(new_n791), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n864), .B1(new_n863), .B2(new_n850), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(G150));
  NAND2_X1  g445(.A1(new_n532), .A2(G55), .ZN(new_n871));
  AOI22_X1  g446(.A1(new_n503), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n872), .A2(new_n505), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n873), .B1(new_n550), .B2(G93), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(G860), .ZN(new_n876));
  XOR2_X1   g451(.A(KEYINPUT108), .B(KEYINPUT37), .Z(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n624), .A2(new_n620), .ZN(new_n879));
  XNOR2_X1  g454(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n879), .B(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT107), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n882), .B1(new_n871), .B2(new_n874), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n871), .A2(new_n882), .A3(new_n874), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(new_n559), .A3(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n559), .B1(new_n884), .B2(new_n885), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n881), .B(new_n889), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n890), .A2(KEYINPUT39), .ZN(new_n891));
  INV_X1    g466(.A(G860), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n892), .B1(new_n890), .B2(KEYINPUT39), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n878), .B1(new_n891), .B2(new_n893), .ZN(G145));
  XNOR2_X1  g469(.A(new_n639), .B(new_n483), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(G160), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n479), .A2(G142), .ZN(new_n898));
  NOR2_X1   g473(.A1(G106), .A2(G2105), .ZN(new_n899));
  OAI21_X1  g474(.A(G2104), .B1(new_n476), .B2(G118), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n477), .A2(KEYINPUT110), .A3(G130), .ZN(new_n901));
  AOI21_X1  g476(.A(KEYINPUT110), .B1(new_n477), .B2(G130), .ZN(new_n902));
  OAI221_X1 g477(.A(new_n898), .B1(new_n899), .B2(new_n900), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(new_n797), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n903), .A2(new_n797), .ZN(new_n906));
  NOR3_X1   g481(.A1(new_n905), .A2(new_n906), .A3(new_n630), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n630), .B1(new_n905), .B2(new_n906), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n908), .A2(KEYINPUT111), .A3(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n777), .B(new_n499), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n911), .A2(new_n725), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n911), .A2(new_n725), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n713), .A2(KEYINPUT109), .ZN(new_n914));
  OR3_X1    g489(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n914), .B1(new_n912), .B2(new_n913), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT111), .ZN(new_n917));
  INV_X1    g492(.A(new_n630), .ZN(new_n918));
  INV_X1    g493(.A(new_n906), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n918), .B1(new_n919), .B2(new_n904), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n917), .B1(new_n920), .B2(new_n907), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n910), .A2(new_n915), .A3(new_n916), .A4(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  AOI22_X1  g498(.A1(new_n910), .A2(new_n921), .B1(new_n915), .B2(new_n916), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n897), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(G37), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n915), .A2(new_n916), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n920), .A2(new_n907), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n922), .B(new_n896), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n925), .A2(new_n926), .A3(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT112), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n925), .A2(KEYINPUT112), .A3(new_n929), .A4(new_n926), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n934), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g510(.A1(new_n613), .A2(new_n620), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n889), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n625), .B1(new_n887), .B2(new_n888), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n617), .A2(new_n624), .ZN(new_n940));
  NAND2_X1  g515(.A1(G299), .A2(new_n613), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n940), .A2(KEYINPUT41), .A3(new_n941), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT41), .B1(new_n940), .B2(new_n941), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n943), .B1(new_n946), .B2(new_n939), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT113), .ZN(new_n948));
  XOR2_X1   g523(.A(G303), .B(G288), .Z(new_n949));
  XNOR2_X1  g524(.A(G290), .B(G305), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n949), .B(new_n950), .ZN(new_n951));
  XOR2_X1   g526(.A(new_n951), .B(KEYINPUT42), .Z(new_n952));
  AND2_X1   g527(.A1(new_n948), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT113), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n943), .B(new_n954), .C1(new_n939), .C2(new_n946), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n952), .B1(new_n948), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(G868), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n875), .A2(new_n622), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(G295));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n958), .ZN(G331));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT43), .ZN(new_n962));
  NAND2_X1  g537(.A1(G286), .A2(G171), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n535), .A2(new_n542), .A3(G301), .A4(new_n543), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n965), .B1(new_n887), .B2(new_n888), .ZN(new_n966));
  INV_X1    g541(.A(new_n885), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n558), .B1(new_n967), .B2(new_n883), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n963), .A2(new_n886), .A3(new_n968), .A4(new_n964), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n970), .B1(new_n945), .B2(new_n944), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n966), .A2(new_n942), .A3(new_n969), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(G37), .B1(new_n973), .B2(new_n951), .ZN(new_n974));
  INV_X1    g549(.A(new_n951), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n971), .A2(new_n975), .A3(new_n972), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n962), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT41), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n942), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n940), .A2(KEYINPUT41), .A3(new_n941), .ZN(new_n980));
  AOI22_X1  g555(.A1(new_n979), .A2(new_n980), .B1(new_n966), .B2(new_n969), .ZN(new_n981));
  INV_X1    g556(.A(new_n972), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n951), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  AND4_X1   g558(.A1(new_n962), .A2(new_n983), .A3(new_n926), .A4(new_n976), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n961), .B1(new_n977), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n974), .A2(new_n962), .A3(new_n976), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n983), .A2(new_n926), .A3(new_n976), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT43), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n986), .A2(new_n988), .A3(KEYINPUT44), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n985), .A2(new_n989), .ZN(G397));
  INV_X1    g565(.A(G1384), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n499), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n464), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT70), .B1(new_n469), .B2(G2105), .ZN(new_n996));
  AOI211_X1 g571(.A(new_n471), .B(new_n476), .C1(new_n467), .C2(new_n468), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n995), .B(G40), .C1(new_n996), .C2(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n994), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G1996), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n725), .B(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G2067), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n777), .B(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n797), .A2(new_n799), .ZN(new_n1004));
  OR2_X1    g579(.A1(new_n797), .A2(new_n799), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1001), .A2(new_n1003), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(G290), .A2(G1986), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n598), .A2(new_n691), .A3(new_n602), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n999), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT119), .ZN(new_n1011));
  NAND2_X1  g586(.A1(G303), .A2(G8), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G8), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n499), .A2(KEYINPUT114), .A3(new_n991), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT114), .B1(new_n499), .B2(new_n991), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT50), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G2090), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n495), .A2(new_n497), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1020), .B1(new_n492), .B2(new_n491), .ZN(new_n1021));
  AOI21_X1  g596(.A(G1384), .B1(new_n1021), .B2(new_n490), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n998), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1018), .A2(new_n1019), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n998), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n499), .A2(KEYINPUT45), .A3(new_n991), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n994), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n829), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1015), .B1(new_n1025), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1011), .B1(new_n1014), .B2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g606(.A(new_n1012), .B(KEYINPUT55), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1025), .A2(new_n1029), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(G8), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1032), .A2(new_n1034), .A3(KEYINPUT119), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1031), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n992), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n499), .A2(KEYINPUT114), .A3(new_n991), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1038), .A2(new_n1026), .A3(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n823), .A2(G1976), .A3(new_n585), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(G8), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT52), .ZN(new_n1043));
  XNOR2_X1  g618(.A(KEYINPUT116), .B(G1976), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT52), .B1(G288), .B2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1045), .A2(new_n1040), .A3(G8), .A4(new_n1041), .ZN(new_n1046));
  AND2_X1   g621(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(G305), .A2(G1981), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n831), .A2(new_n696), .A3(new_n590), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1048), .A2(new_n1049), .A3(KEYINPUT49), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1015), .B1(new_n1051), .B2(new_n1026), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT117), .B(KEYINPUT49), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1053), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1054), .A2(KEYINPUT118), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n1056));
  AOI211_X1 g631(.A(new_n1056), .B(new_n1053), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1050), .B(new_n1052), .C1(new_n1055), .C2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1047), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(KEYINPUT115), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n992), .A2(new_n1062), .A3(KEYINPUT50), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n998), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1038), .A2(new_n1023), .A3(new_n1039), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1029), .B1(new_n1066), .B2(G2090), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1067), .A2(new_n1014), .A3(G8), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1036), .A2(new_n1060), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT126), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1036), .A2(new_n1060), .A3(KEYINPUT126), .A4(new_n1068), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1018), .A2(new_n1024), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1028), .ZN(new_n1075));
  XNOR2_X1  g650(.A(KEYINPUT56), .B(G2072), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n735), .A2(new_n1074), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  XNOR2_X1  g652(.A(KEYINPUT121), .B(KEYINPUT57), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n573), .A2(new_n581), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1078), .B1(new_n573), .B2(new_n581), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1077), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1077), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT122), .B1(new_n1051), .B2(new_n1026), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT122), .ZN(new_n1084));
  NOR4_X1   g659(.A1(new_n1016), .A2(new_n1017), .A3(new_n998), .A4(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1002), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G1348), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1062), .B1(new_n992), .B2(KEYINPUT50), .ZN(new_n1088));
  AOI211_X1 g663(.A(KEYINPUT115), .B(new_n1023), .C1(new_n499), .C2(new_n991), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1026), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1065), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1087), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n624), .B1(new_n1086), .B2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1081), .B1(new_n1082), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT60), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1040), .A2(new_n1084), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1051), .A2(KEYINPUT122), .A3(new_n1026), .ZN(new_n1097));
  AOI21_X1  g672(.A(G2067), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(G1348), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1095), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1086), .A2(new_n1092), .A3(KEYINPUT60), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1100), .A2(new_n1101), .A3(new_n613), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1081), .A2(KEYINPUT61), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT61), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1077), .B(new_n1104), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1086), .A2(new_n1092), .A3(KEYINPUT60), .A4(new_n624), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1102), .A2(new_n1103), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT123), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT59), .ZN(new_n1109));
  XOR2_X1   g684(.A(KEYINPUT58), .B(G1341), .Z(new_n1110));
  NAND3_X1  g685(.A1(new_n1096), .A2(new_n1097), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1075), .A2(new_n1000), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n558), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1108), .A2(KEYINPUT59), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1109), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1114), .ZN(new_n1116));
  AOI211_X1 g691(.A(new_n558), .B(new_n1116), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1094), .B1(new_n1107), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1066), .A2(new_n766), .ZN(new_n1120));
  AOI21_X1  g695(.A(KEYINPUT45), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(G2078), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1123), .A2(KEYINPUT53), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT53), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1126), .B1(new_n1028), .B2(G2078), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1120), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  AND2_X1   g703(.A1(G301), .A2(KEYINPUT54), .ZN(new_n1129));
  NOR2_X1   g704(.A1(G301), .A2(KEYINPUT54), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1128), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1132));
  NAND2_X1  g707(.A1(KEYINPUT53), .A2(G40), .ZN(new_n1133));
  OR2_X1    g708(.A1(new_n1124), .A2(KEYINPUT125), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1124), .A2(KEYINPUT125), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1133), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n995), .A2(new_n470), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n994), .A2(new_n1027), .A3(new_n1137), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1120), .A2(new_n1127), .A3(new_n1132), .A4(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1131), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT51), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1015), .B1(KEYINPUT124), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1143), .A2(new_n705), .A3(new_n1065), .A4(new_n1026), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n784), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  OAI221_X1 g721(.A(new_n1142), .B1(KEYINPUT124), .B2(new_n1141), .C1(new_n1146), .C2(G286), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1142), .B1(new_n1146), .B2(G286), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1141), .A2(KEYINPUT124), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1015), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1150));
  AOI22_X1  g725(.A1(new_n1148), .A2(new_n1149), .B1(G286), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1140), .B1(new_n1147), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1119), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1151), .A2(new_n1147), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(KEYINPUT62), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT62), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1151), .A2(new_n1156), .A3(new_n1147), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1128), .A2(G171), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1155), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1073), .B1(new_n1153), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT63), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1150), .A2(new_n1161), .A3(G168), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1162), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n1014), .A2(new_n1030), .A3(new_n1011), .ZN(new_n1164));
  AOI21_X1  g739(.A(KEYINPUT119), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1163), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1059), .B1(new_n1166), .B2(new_n1068), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1047), .A2(new_n1058), .A3(G168), .A4(new_n1150), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1014), .B1(new_n1067), .B2(G8), .ZN(new_n1169));
  OAI21_X1  g744(.A(KEYINPUT63), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  OR2_X1    g745(.A1(G288), .A2(G1976), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1058), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(new_n1049), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(new_n1052), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1170), .A2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(KEYINPUT120), .B1(new_n1167), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1162), .B1(new_n1031), .B2(new_n1035), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1068), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1060), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT120), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1180), .A2(new_n1181), .A3(new_n1175), .A4(new_n1170), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1177), .A2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1010), .B1(new_n1160), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT46), .ZN(new_n1185));
  INV_X1    g760(.A(new_n999), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1185), .B1(new_n1186), .B2(G1996), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1003), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n999), .B1(new_n1188), .B2(new_n725), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n999), .A2(KEYINPUT46), .A3(new_n1000), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1187), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  XOR2_X1   g766(.A(new_n1191), .B(KEYINPUT47), .Z(new_n1192));
  NAND2_X1  g767(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1004), .B1(new_n1193), .B2(new_n999), .ZN(new_n1194));
  INV_X1    g769(.A(new_n777), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1194), .B1(new_n1002), .B2(new_n1195), .ZN(new_n1196));
  AND2_X1   g771(.A1(new_n1196), .A2(KEYINPUT127), .ZN(new_n1197));
  NOR2_X1   g772(.A1(new_n1196), .A2(KEYINPUT127), .ZN(new_n1198));
  NOR3_X1   g773(.A1(new_n1197), .A2(new_n1198), .A3(new_n1186), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1006), .A2(new_n999), .ZN(new_n1200));
  NOR2_X1   g775(.A1(new_n1186), .A2(new_n1008), .ZN(new_n1201));
  XOR2_X1   g776(.A(new_n1201), .B(KEYINPUT48), .Z(new_n1202));
  AOI211_X1 g777(.A(new_n1192), .B(new_n1199), .C1(new_n1200), .C2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1184), .A2(new_n1203), .ZN(G329));
  assign    G231 = 1'b0;
  NAND4_X1  g779(.A1(new_n698), .A2(G319), .A3(new_n659), .A4(new_n676), .ZN(new_n1206));
  AOI221_X4 g780(.A(new_n1206), .B1(new_n932), .B2(new_n933), .C1(new_n988), .C2(new_n986), .ZN(G308));
  AOI21_X1  g781(.A(new_n1206), .B1(new_n932), .B2(new_n933), .ZN(new_n1208));
  OAI21_X1  g782(.A(new_n1208), .B1(new_n977), .B2(new_n984), .ZN(G225));
endmodule


