//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 1 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032;
  XOR2_X1   g000(.A(KEYINPUT9), .B(G234), .Z(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT78), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G221), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n191), .B(KEYINPUT79), .ZN(new_n192));
  INV_X1    g006(.A(G104), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT3), .B1(new_n193), .B2(G107), .ZN(new_n194));
  AOI21_X1  g008(.A(G101), .B1(new_n193), .B2(G107), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT3), .ZN(new_n196));
  INV_X1    g010(.A(G107), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n197), .A3(G104), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n194), .A2(new_n195), .A3(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT81), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT81), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n194), .A2(new_n195), .A3(new_n198), .A4(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n193), .A2(G107), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n194), .A2(new_n198), .A3(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G101), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT80), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n205), .A2(KEYINPUT80), .A3(G101), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n203), .A2(new_n208), .A3(KEYINPUT4), .A4(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT64), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(KEYINPUT64), .A2(G146), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(G143), .A3(new_n215), .ZN(new_n216));
  AND2_X1   g030(.A1(KEYINPUT0), .A2(G128), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n213), .A2(G143), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  AND3_X1   g033(.A1(new_n216), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT0), .B(G128), .ZN(new_n221));
  INV_X1    g035(.A(G143), .ZN(new_n222));
  AND2_X1   g036(.A1(KEYINPUT64), .A2(G146), .ZN(new_n223));
  NOR2_X1   g037(.A1(KEYINPUT64), .A2(G146), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n222), .A2(G146), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n221), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n211), .B1(new_n220), .B2(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(KEYINPUT0), .A2(G128), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n217), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(G143), .B1(new_n214), .B2(new_n215), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n231), .B1(new_n232), .B2(new_n226), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n216), .A2(new_n217), .A3(new_n219), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n233), .A2(KEYINPUT66), .A3(new_n234), .ZN(new_n235));
  XOR2_X1   g049(.A(KEYINPUT82), .B(KEYINPUT4), .Z(new_n236));
  NAND3_X1  g050(.A1(new_n205), .A2(G101), .A3(new_n236), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n210), .A2(new_n229), .A3(new_n235), .A4(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G137), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(KEYINPUT11), .A3(G134), .ZN(new_n240));
  INV_X1    g054(.A(G134), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G137), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT65), .ZN(new_n244));
  INV_X1    g058(.A(G131), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT11), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n246), .B1(new_n241), .B2(G137), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n243), .A2(new_n244), .A3(new_n245), .A4(new_n247), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n247), .A2(new_n240), .A3(new_n245), .A4(new_n242), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT65), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n243), .A2(new_n247), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n248), .A2(new_n250), .B1(new_n251), .B2(G131), .ZN(new_n252));
  INV_X1    g066(.A(G101), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n197), .A2(G104), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n253), .B1(new_n254), .B2(new_n204), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n255), .B1(new_n200), .B2(new_n202), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT1), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n216), .A2(new_n257), .A3(G128), .A4(new_n219), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n223), .A2(new_n224), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n218), .B1(new_n259), .B2(G143), .ZN(new_n260));
  INV_X1    g074(.A(G128), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n261), .B1(new_n227), .B2(KEYINPUT1), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n258), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n256), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT10), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n261), .B1(new_n216), .B2(KEYINPUT1), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n232), .A2(new_n226), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n258), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(new_n256), .A3(KEYINPUT10), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n238), .A2(new_n252), .A3(new_n266), .A4(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n210), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n229), .A2(new_n235), .A3(new_n237), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n266), .B(new_n270), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n252), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT83), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n275), .A2(KEYINPUT83), .A3(new_n276), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n272), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  XNOR2_X1  g095(.A(G110), .B(G140), .ZN(new_n282));
  INV_X1    g096(.A(G953), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n283), .A2(G227), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n282), .B(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n264), .B1(new_n269), .B2(new_n256), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n287), .A2(KEYINPUT12), .A3(new_n276), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT12), .B1(new_n287), .B2(new_n276), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n271), .A2(new_n286), .ZN(new_n291));
  OAI22_X1  g105(.A1(new_n281), .A2(new_n286), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G469), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n292), .A2(new_n293), .A3(new_n189), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n279), .A2(new_n280), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n271), .A2(new_n286), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n271), .B1(new_n288), .B2(new_n289), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n295), .A2(new_n296), .B1(new_n285), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(G469), .B1(new_n298), .B2(G902), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n192), .B1(new_n294), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT20), .ZN(new_n302));
  INV_X1    g116(.A(G214), .ZN(new_n303));
  NOR3_X1   g117(.A1(new_n303), .A2(G237), .A3(G953), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT90), .ZN(new_n305));
  AOI21_X1  g119(.A(KEYINPUT91), .B1(new_n305), .B2(new_n222), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT91), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n307), .A2(G143), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n304), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G237), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(new_n283), .A3(G214), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n307), .B1(KEYINPUT90), .B2(G143), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n309), .A2(new_n245), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT17), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n309), .A2(new_n313), .ZN(new_n316));
  AOI21_X1  g130(.A(KEYINPUT92), .B1(new_n316), .B2(G131), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT92), .ZN(new_n318));
  AOI211_X1 g132(.A(new_n318), .B(new_n245), .C1(new_n309), .C2(new_n313), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n314), .B(new_n315), .C1(new_n317), .C2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT95), .ZN(new_n321));
  INV_X1    g135(.A(G140), .ZN(new_n322));
  INV_X1    g136(.A(G125), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n322), .B1(new_n323), .B2(KEYINPUT72), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT72), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(G125), .A3(G140), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(KEYINPUT16), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT16), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n328), .B1(new_n323), .B2(G140), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G146), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n327), .A2(new_n213), .A3(new_n329), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n317), .A2(new_n319), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n333), .B1(new_n334), .B2(KEYINPUT17), .ZN(new_n335));
  INV_X1    g149(.A(new_n314), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n222), .A2(KEYINPUT91), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n311), .B1(new_n312), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n305), .A2(new_n222), .ZN(new_n339));
  NOR2_X1   g153(.A1(G237), .A2(G953), .ZN(new_n340));
  AOI22_X1  g154(.A1(new_n339), .A2(new_n307), .B1(new_n340), .B2(G214), .ZN(new_n341));
  OAI21_X1  g155(.A(G131), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n318), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n316), .A2(KEYINPUT92), .A3(G131), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n336), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT95), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(new_n346), .A3(new_n315), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n321), .A2(new_n335), .A3(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(G125), .B(G140), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n259), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n324), .A2(new_n326), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n350), .B1(new_n351), .B2(new_n213), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT18), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n353), .A2(new_n245), .ZN(new_n354));
  OAI221_X1 g168(.A(new_n352), .B1(new_n316), .B2(new_n354), .C1(new_n342), .C2(new_n353), .ZN(new_n355));
  XNOR2_X1  g169(.A(G113), .B(G122), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT94), .B(G104), .ZN(new_n357));
  XOR2_X1   g171(.A(new_n356), .B(new_n357), .Z(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n348), .A2(new_n355), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT19), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n349), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n362), .B1(new_n351), .B2(new_n361), .ZN(new_n363));
  INV_X1    g177(.A(new_n259), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n331), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n355), .B1(new_n345), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT93), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n355), .B(KEYINPUT93), .C1(new_n345), .C2(new_n365), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n358), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n360), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(G475), .A2(G902), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n302), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n372), .ZN(new_n374));
  AOI211_X1 g188(.A(KEYINPUT20), .B(new_n374), .C1(new_n360), .C2(new_n370), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n348), .A2(new_n355), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n358), .ZN(new_n377));
  AOI21_X1  g191(.A(G902), .B1(new_n377), .B2(new_n360), .ZN(new_n378));
  INV_X1    g192(.A(G475), .ZN(new_n379));
  OAI22_X1  g193(.A1(new_n373), .A2(new_n375), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT97), .ZN(new_n381));
  INV_X1    g195(.A(G122), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G116), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n197), .B1(new_n383), .B2(KEYINPUT14), .ZN(new_n384));
  INV_X1    g198(.A(G116), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G122), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  OR2_X1    g201(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n384), .A2(new_n387), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n261), .A2(G143), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n391), .B(KEYINPUT96), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n222), .A2(G128), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G134), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n392), .A2(new_n241), .A3(new_n393), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n390), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n396), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n393), .B(KEYINPUT13), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n241), .B1(new_n392), .B2(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n387), .B(new_n197), .ZN(new_n402));
  OR3_X1    g216(.A1(new_n399), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n188), .A2(G217), .A3(new_n283), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n398), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  NOR3_X1   g220(.A1(new_n399), .A2(new_n401), .A3(new_n402), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n404), .B1(new_n407), .B2(new_n397), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n381), .B1(new_n409), .B2(new_n189), .ZN(new_n410));
  INV_X1    g224(.A(G478), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(KEYINPUT15), .ZN(new_n412));
  OR2_X1    g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  AOI211_X1 g227(.A(KEYINPUT97), .B(G902), .C1(new_n406), .C2(new_n408), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n412), .B1(new_n410), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n380), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G952), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n419), .A2(G953), .ZN(new_n420));
  NAND2_X1  g234(.A1(G234), .A2(G237), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n421), .A2(G902), .A3(G953), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT21), .B(G898), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n423), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(G214), .B1(G237), .B2(G902), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(G210), .B1(G237), .B2(G902), .ZN(new_n431));
  XOR2_X1   g245(.A(new_n431), .B(KEYINPUT89), .Z(new_n432));
  XNOR2_X1  g246(.A(G110), .B(G122), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT84), .ZN(new_n435));
  XOR2_X1   g249(.A(KEYINPUT2), .B(G113), .Z(new_n436));
  XNOR2_X1  g250(.A(G116), .B(G119), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G119), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G116), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n385), .A2(G119), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(KEYINPUT2), .B(G113), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n438), .A2(new_n444), .ZN(new_n445));
  AND2_X1   g259(.A1(new_n445), .A2(new_n237), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n210), .A2(new_n435), .A3(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(G113), .B1(new_n440), .B2(KEYINPUT5), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n437), .A2(KEYINPUT5), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n438), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n256), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n447), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n435), .B1(new_n210), .B2(new_n446), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n434), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n210), .A2(new_n446), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(KEYINPUT84), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n459), .A2(new_n433), .A3(new_n454), .A4(new_n447), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n457), .A2(KEYINPUT6), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n233), .A2(new_n234), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(G125), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n323), .B(new_n258), .C1(new_n267), .C2(new_n268), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(KEYINPUT85), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT85), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n283), .A2(G224), .ZN(new_n470));
  XOR2_X1   g284(.A(new_n470), .B(KEYINPUT86), .Z(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n466), .A2(new_n468), .A3(new_n471), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT6), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n476), .B(new_n434), .C1(new_n455), .C2(new_n456), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n461), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT87), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n448), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g294(.A(KEYINPUT87), .B(G113), .C1(new_n440), .C2(KEYINPUT5), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n480), .A2(new_n450), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n438), .ZN(new_n483));
  AND2_X1   g297(.A1(new_n483), .A2(new_n256), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n433), .B(KEYINPUT8), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n485), .B1(new_n256), .B2(new_n452), .ZN(new_n486));
  OAI21_X1  g300(.A(KEYINPUT88), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n255), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n203), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n453), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n483), .A2(new_n256), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT88), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n490), .A2(new_n491), .A3(new_n492), .A4(new_n485), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n487), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n466), .A2(KEYINPUT7), .A3(new_n468), .A4(new_n470), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n470), .A2(KEYINPUT7), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n465), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n494), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n460), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n189), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n432), .B1(new_n478), .B2(new_n500), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n494), .A2(new_n495), .A3(new_n497), .ZN(new_n502));
  AOI21_X1  g316(.A(G902), .B1(new_n502), .B2(new_n460), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n461), .A2(new_n475), .A3(new_n477), .ZN(new_n504));
  INV_X1    g318(.A(new_n432), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n430), .B1(new_n501), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NOR3_X1   g322(.A1(new_n301), .A2(new_n418), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT77), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT32), .ZN(new_n511));
  XOR2_X1   g325(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n512));
  NAND2_X1  g326(.A1(new_n340), .A2(G210), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n512), .B(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT26), .B(G101), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n514), .B(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT28), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT68), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n239), .A2(G134), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n245), .B1(new_n519), .B2(new_n242), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n520), .B1(new_n248), .B2(new_n250), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT67), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n269), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI211_X1 g337(.A(KEYINPUT67), .B(new_n520), .C1(new_n248), .C2(new_n250), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n518), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n233), .A2(KEYINPUT66), .A3(new_n234), .ZN(new_n526));
  AOI21_X1  g340(.A(KEYINPUT66), .B1(new_n233), .B2(new_n234), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n445), .B1(new_n528), .B2(new_n276), .ZN(new_n529));
  INV_X1    g343(.A(new_n520), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n249), .A2(KEYINPUT65), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n249), .A2(KEYINPUT65), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT67), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n521), .A2(new_n522), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n534), .A2(new_n535), .A3(KEYINPUT68), .A4(new_n269), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n525), .A2(new_n529), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n521), .A2(new_n269), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n538), .B1(new_n252), .B2(new_n462), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n445), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n517), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n534), .A2(new_n535), .A3(new_n269), .ZN(new_n542));
  AOI21_X1  g356(.A(KEYINPUT28), .B1(new_n529), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n516), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n516), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n537), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT31), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT30), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n548), .B1(new_n528), .B2(new_n276), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n525), .A2(new_n549), .A3(new_n536), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n539), .A2(new_n548), .B1(new_n444), .B2(new_n438), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n546), .A2(new_n547), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n544), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT70), .ZN(new_n555));
  AOI211_X1 g369(.A(new_n555), .B(new_n547), .C1(new_n546), .C2(new_n552), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n552), .A2(new_n537), .A3(new_n545), .ZN(new_n557));
  AOI21_X1  g371(.A(KEYINPUT70), .B1(new_n557), .B2(KEYINPUT31), .ZN(new_n558));
  NOR3_X1   g372(.A1(new_n554), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(G472), .A2(G902), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n511), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n550), .A2(new_n551), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n537), .A2(new_n545), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT31), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n555), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n557), .A2(KEYINPUT70), .A3(KEYINPUT31), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n566), .A2(new_n544), .A3(new_n553), .A4(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n561), .A2(new_n511), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT29), .ZN(new_n570));
  NOR3_X1   g384(.A1(new_n543), .A2(new_n570), .A3(new_n516), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n525), .A2(new_n536), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n528), .A2(new_n276), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n525), .A2(new_n573), .A3(new_n536), .ZN(new_n574));
  AOI22_X1  g388(.A1(new_n572), .A2(new_n529), .B1(new_n574), .B2(new_n445), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n571), .B1(new_n575), .B2(new_n517), .ZN(new_n576));
  AOI22_X1  g390(.A1(new_n572), .A2(new_n529), .B1(new_n550), .B2(new_n551), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n570), .B1(new_n577), .B2(new_n545), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n529), .A2(new_n542), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n517), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n545), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n581), .A2(new_n541), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n189), .B(new_n576), .C1(new_n578), .C2(new_n582), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n568), .A2(new_n569), .B1(new_n583), .B2(G472), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n562), .A2(new_n584), .ZN(new_n585));
  XOR2_X1   g399(.A(KEYINPUT24), .B(G110), .Z(new_n586));
  XNOR2_X1  g400(.A(G119), .B(G128), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT23), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n589), .B1(new_n439), .B2(G128), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n261), .A2(KEYINPUT23), .A3(G119), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n590), .B(new_n591), .C1(G119), .C2(new_n261), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT71), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n593), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(G110), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n333), .B(new_n588), .C1(new_n594), .C2(new_n596), .ZN(new_n597));
  OAI22_X1  g411(.A1(new_n592), .A2(G110), .B1(new_n586), .B2(new_n587), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n331), .A2(new_n598), .A3(new_n350), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(KEYINPUT22), .B(G137), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(G221), .A2(G234), .ZN(new_n603));
  OR3_X1    g417(.A1(new_n603), .A2(KEYINPUT73), .A3(G953), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT74), .ZN(new_n605));
  OAI21_X1  g419(.A(KEYINPUT73), .B1(new_n603), .B2(G953), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n605), .B1(new_n604), .B2(new_n606), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n602), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n609), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n611), .A2(new_n601), .A3(new_n607), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n610), .A2(new_n612), .A3(KEYINPUT75), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT75), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n601), .B1(new_n611), .B2(new_n607), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n608), .A2(new_n602), .A3(new_n609), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n600), .A2(new_n613), .A3(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n599), .A2(new_n597), .A3(new_n612), .A4(new_n610), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT76), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(G217), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n623), .B1(G234), .B2(new_n189), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n622), .A2(G902), .A3(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n624), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n618), .A2(new_n189), .A3(new_n619), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT25), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n618), .A2(KEYINPUT25), .A3(new_n189), .A4(new_n619), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n626), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n625), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n510), .B1(new_n585), .B2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n632), .ZN(new_n634));
  AOI211_X1 g448(.A(KEYINPUT77), .B(new_n634), .C1(new_n562), .C2(new_n584), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n509), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G101), .ZN(G3));
  INV_X1    g451(.A(new_n429), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n505), .B1(new_n503), .B2(new_n504), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT99), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n501), .A2(KEYINPUT99), .A3(new_n506), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT33), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n644), .B1(new_n404), .B2(KEYINPUT100), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n409), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n406), .A2(new_n408), .A3(new_n645), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n411), .A2(G902), .ZN(new_n649));
  AND4_X1   g463(.A1(KEYINPUT101), .A2(new_n647), .A3(new_n648), .A4(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n409), .A2(new_n189), .ZN(new_n652));
  AOI21_X1  g466(.A(KEYINPUT101), .B1(new_n652), .B2(new_n411), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n650), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n380), .A2(new_n654), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n643), .A2(new_n427), .A3(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  OAI211_X1 g471(.A(KEYINPUT98), .B(G472), .C1(new_n559), .C2(G902), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT98), .ZN(new_n659));
  INV_X1    g473(.A(G472), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n568), .B(new_n189), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n658), .A2(new_n632), .A3(new_n661), .A4(new_n300), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n657), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT34), .B(G104), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G6));
  INV_X1    g479(.A(new_n380), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n416), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n643), .A2(new_n667), .A3(new_n427), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n662), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT35), .B(G107), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G9));
  NAND2_X1  g486(.A1(new_n658), .A2(new_n661), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n617), .A2(new_n613), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT36), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n600), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n674), .A2(new_n675), .A3(new_n597), .A4(new_n599), .ZN(new_n678));
  AND4_X1   g492(.A1(new_n189), .A2(new_n677), .A3(new_n626), .A4(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n631), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n300), .A2(new_n417), .A3(new_n507), .A4(new_n681), .ZN(new_n682));
  OR2_X1    g496(.A1(new_n673), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT37), .B(G110), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G12));
  INV_X1    g499(.A(new_n192), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n290), .A2(new_n291), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n225), .A2(new_n227), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n257), .B1(new_n259), .B2(G143), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n688), .B1(new_n689), .B2(new_n261), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n265), .B1(new_n690), .B2(new_n258), .ZN(new_n691));
  AOI22_X1  g505(.A1(new_n256), .A2(new_n691), .B1(new_n264), .B2(new_n265), .ZN(new_n692));
  AOI211_X1 g506(.A(new_n278), .B(new_n252), .C1(new_n692), .C2(new_n238), .ZN(new_n693));
  AOI21_X1  g507(.A(KEYINPUT83), .B1(new_n275), .B2(new_n276), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n271), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n687), .B1(new_n695), .B2(new_n285), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n696), .A2(G469), .A3(G902), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n296), .B1(new_n693), .B2(new_n694), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n297), .A2(new_n285), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n293), .B1(new_n700), .B2(new_n189), .ZN(new_n701));
  OAI211_X1 g515(.A(new_n686), .B(new_n681), .C1(new_n697), .C2(new_n701), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n702), .B1(new_n562), .B2(new_n584), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n641), .A2(new_n642), .ZN(new_n704));
  INV_X1    g518(.A(G900), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n423), .B1(new_n425), .B2(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n667), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n703), .A2(new_n704), .A3(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(KEYINPUT102), .B(G128), .Z(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G30));
  XOR2_X1   g524(.A(new_n706), .B(KEYINPUT39), .Z(new_n711));
  NAND2_X1  g525(.A1(new_n300), .A2(new_n711), .ZN(new_n712));
  XOR2_X1   g526(.A(new_n712), .B(KEYINPUT40), .Z(new_n713));
  NAND2_X1  g527(.A1(new_n575), .A2(new_n516), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n552), .A2(new_n537), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n545), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n714), .A2(new_n716), .A3(new_n189), .ZN(new_n717));
  AOI22_X1  g531(.A1(new_n568), .A2(new_n569), .B1(G472), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n562), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(new_n506), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n721), .B1(new_n722), .B2(new_n639), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n501), .A2(new_n506), .A3(new_n720), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n416), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n666), .A2(new_n726), .ZN(new_n727));
  AND4_X1   g541(.A1(new_n429), .A2(new_n725), .A3(new_n727), .A4(new_n680), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n713), .A2(new_n719), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G143), .ZN(G45));
  INV_X1    g544(.A(new_n706), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n380), .A2(new_n654), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT104), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(new_n703), .A3(new_n704), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G146), .ZN(G48));
  AOI21_X1  g550(.A(new_n634), .B1(new_n562), .B2(new_n584), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n293), .A2(KEYINPUT105), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n292), .A2(new_n189), .A3(new_n739), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n738), .B1(new_n696), .B2(G902), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n740), .A2(new_n741), .A3(new_n191), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n737), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n744), .A2(new_n657), .ZN(new_n745));
  XOR2_X1   g559(.A(KEYINPUT41), .B(G113), .Z(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(G15));
  NOR2_X1   g561(.A1(new_n744), .A2(new_n669), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(new_n385), .ZN(G18));
  NOR4_X1   g563(.A1(new_n380), .A2(new_n680), .A3(new_n416), .A4(new_n427), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n545), .B1(new_n552), .B2(new_n537), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n582), .A2(new_n751), .A3(KEYINPUT29), .ZN(new_n752));
  INV_X1    g566(.A(new_n571), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n574), .A2(new_n445), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n517), .B1(new_n754), .B2(new_n537), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n189), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g570(.A(G472), .B1(new_n752), .B2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n569), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n757), .B1(new_n559), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(KEYINPUT32), .B1(new_n568), .B2(new_n560), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n750), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n704), .A2(new_n743), .ZN(new_n762));
  OAI21_X1  g576(.A(KEYINPUT106), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n643), .A2(new_n742), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT106), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n585), .A2(new_n764), .A3(new_n765), .A4(new_n750), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G119), .ZN(G21));
  AOI21_X1  g582(.A(new_n660), .B1(new_n568), .B2(new_n189), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n565), .A2(new_n553), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n516), .B1(new_n755), .B2(new_n543), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n561), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n769), .A2(new_n634), .A3(new_n772), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n643), .A2(new_n666), .A3(new_n726), .ZN(new_n774));
  AND4_X1   g588(.A1(new_n428), .A2(new_n740), .A3(new_n741), .A4(new_n191), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n773), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G122), .ZN(G24));
  NOR3_X1   g591(.A1(new_n769), .A2(new_n680), .A3(new_n772), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n734), .A2(new_n764), .A3(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(KEYINPUT107), .B(G125), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n779), .B(new_n780), .ZN(G27));
  OAI21_X1  g595(.A(KEYINPUT108), .B1(new_n697), .B2(new_n701), .ZN(new_n782));
  AND4_X1   g596(.A1(new_n501), .A2(new_n506), .A3(new_n429), .A4(new_n191), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT108), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n294), .A2(new_n299), .A3(new_n784), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n782), .A2(new_n783), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n734), .A2(new_n737), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT42), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n734), .A2(new_n737), .A3(KEYINPUT42), .A4(new_n786), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G131), .ZN(G33));
  NAND3_X1  g606(.A1(new_n737), .A2(new_n707), .A3(new_n786), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT109), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT109), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n737), .A2(new_n786), .A3(new_n795), .A4(new_n707), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G134), .ZN(G36));
  INV_X1    g612(.A(new_n654), .ZN(new_n799));
  OAI21_X1  g613(.A(KEYINPUT43), .B1(new_n799), .B2(new_n380), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT43), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n666), .A2(new_n801), .A3(new_n654), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n803), .A2(new_n673), .A3(new_n681), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT44), .ZN(new_n805));
  OAI211_X1 g619(.A(KEYINPUT110), .B(G469), .C1(new_n298), .C2(KEYINPUT45), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT110), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT45), .B1(new_n698), .B2(new_n699), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n807), .B1(new_n808), .B2(new_n293), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n298), .A2(KEYINPUT45), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n806), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(G469), .A2(G902), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT46), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT111), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n811), .A2(KEYINPUT46), .A3(new_n812), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n818), .A2(new_n294), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n813), .A2(KEYINPUT111), .A3(new_n814), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n817), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(new_n191), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n501), .A2(new_n506), .A3(new_n429), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(KEYINPUT112), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n805), .A2(new_n823), .A3(new_n711), .A4(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(G137), .ZN(G39));
  NOR3_X1   g641(.A1(new_n585), .A2(new_n632), .A3(new_n824), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n821), .A2(KEYINPUT47), .A3(new_n191), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT47), .B1(new_n821), .B2(new_n191), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n734), .B(new_n828), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(G140), .ZN(G42));
  INV_X1    g646(.A(KEYINPUT114), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n834));
  AOI22_X1  g648(.A1(new_n789), .A2(new_n790), .B1(new_n794), .B2(new_n796), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n585), .A2(new_n632), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT77), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n737), .A2(new_n510), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI22_X1  g653(.A1(new_n839), .A2(new_n509), .B1(new_n766), .B2(new_n763), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n737), .B(new_n743), .C1(new_n668), .C2(new_n656), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n301), .A2(new_n634), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n508), .B1(new_n667), .B2(new_n655), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n842), .A2(new_n843), .A3(new_n661), .A4(new_n658), .ZN(new_n844));
  AND4_X1   g658(.A1(new_n683), .A2(new_n841), .A3(new_n776), .A4(new_n844), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n732), .A2(KEYINPUT104), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n732), .A2(KEYINPUT104), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n778), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n418), .A2(new_n706), .A3(new_n824), .ZN(new_n849));
  AOI22_X1  g663(.A1(new_n848), .A2(new_n786), .B1(new_n703), .B2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n835), .A2(new_n840), .A3(new_n845), .A4(new_n850), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n680), .A2(new_n191), .A3(new_n731), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n782), .A2(new_n852), .A3(new_n785), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n774), .A2(new_n853), .A3(new_n719), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n735), .A2(new_n779), .A3(new_n708), .A4(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT52), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n704), .B(new_n703), .C1(new_n734), .C2(new_n707), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT52), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n857), .A2(new_n858), .A3(new_n779), .A4(new_n854), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n834), .B1(new_n851), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n791), .A2(new_n797), .A3(new_n850), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n704), .A2(new_n775), .A3(new_n727), .ZN(new_n863));
  OAI21_X1  g677(.A(G472), .B1(new_n559), .B2(G902), .ZN(new_n864));
  INV_X1    g678(.A(new_n772), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n864), .A2(new_n632), .A3(new_n865), .ZN(new_n866));
  OAI22_X1  g680(.A1(new_n863), .A2(new_n866), .B1(new_n673), .B2(new_n682), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n655), .B1(new_n380), .B2(new_n726), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(new_n507), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n662), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n871), .A2(new_n636), .A3(new_n767), .A4(new_n841), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n862), .A2(new_n872), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n856), .A2(new_n859), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n873), .A2(KEYINPUT53), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n833), .B1(new_n861), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT53), .B1(new_n873), .B2(new_n874), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n877), .A2(KEYINPUT114), .ZN(new_n878));
  OAI21_X1  g692(.A(KEYINPUT54), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n742), .A2(new_n824), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n803), .A2(new_n778), .A3(new_n423), .A4(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n719), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n882), .A2(new_n632), .A3(new_n423), .A4(new_n880), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n666), .A2(new_n799), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT118), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n886), .A2(KEYINPUT50), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n742), .A2(new_n429), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT117), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n888), .A2(new_n889), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n724), .B(new_n723), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n803), .A2(new_n773), .A3(new_n423), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n887), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n888), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(KEYINPUT117), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n725), .B1(new_n897), .B2(new_n890), .ZN(new_n898));
  INV_X1    g712(.A(new_n894), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n898), .B(new_n899), .C1(new_n886), .C2(KEYINPUT50), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n885), .B1(new_n895), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n740), .A2(new_n741), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n902), .A2(new_n686), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n829), .A2(new_n830), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n899), .A2(new_n825), .ZN(new_n905));
  OAI211_X1 g719(.A(KEYINPUT51), .B(new_n901), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  AND4_X1   g720(.A1(new_n737), .A2(new_n803), .A3(new_n423), .A4(new_n880), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n907), .A2(KEYINPUT119), .A3(KEYINPUT48), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n420), .B1(new_n883), .B2(new_n655), .ZN(new_n909));
  XNOR2_X1  g723(.A(KEYINPUT119), .B(KEYINPUT48), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  AOI211_X1 g725(.A(new_n909), .B(new_n911), .C1(new_n764), .C2(new_n899), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n906), .A2(new_n908), .A3(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT115), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n914), .B1(new_n829), .B2(new_n830), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT47), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n822), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n821), .A2(KEYINPUT47), .A3(new_n191), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n917), .A2(KEYINPUT115), .A3(new_n918), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n903), .B(KEYINPUT116), .Z(new_n920));
  AND3_X1   g734(.A1(new_n915), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n901), .B1(new_n921), .B2(new_n905), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT51), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n913), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n861), .A2(new_n875), .ZN(new_n925));
  OR2_X1    g739(.A1(new_n925), .A2(KEYINPUT54), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n879), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n419), .A2(new_n283), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n632), .A2(new_n429), .A3(new_n686), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT113), .ZN(new_n931));
  NOR4_X1   g745(.A1(new_n931), .A2(new_n380), .A3(new_n799), .A4(new_n725), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n902), .B(KEYINPUT49), .Z(new_n933));
  NAND3_X1  g747(.A1(new_n932), .A2(new_n882), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n929), .A2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT120), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n929), .A2(KEYINPUT120), .A3(new_n934), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(G75));
  AOI21_X1  g753(.A(new_n189), .B1(new_n861), .B2(new_n875), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n940), .A2(KEYINPUT122), .A3(new_n432), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT56), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n461), .A2(new_n477), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(new_n475), .ZN(new_n944));
  XOR2_X1   g758(.A(KEYINPUT121), .B(KEYINPUT55), .Z(new_n945));
  XNOR2_X1  g759(.A(new_n944), .B(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n941), .A2(new_n942), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(KEYINPUT122), .B1(new_n940), .B2(new_n432), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n283), .A2(G952), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT56), .B1(new_n940), .B2(new_n432), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n951), .B1(new_n952), .B2(new_n946), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n949), .A2(new_n953), .ZN(G51));
  XNOR2_X1  g768(.A(new_n925), .B(KEYINPUT54), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n812), .B(KEYINPUT57), .Z(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n292), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n811), .B(KEYINPUT123), .Z(new_n959));
  NAND2_X1  g773(.A1(new_n940), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n950), .B1(new_n958), .B2(new_n960), .ZN(G54));
  NAND3_X1  g775(.A1(new_n940), .A2(KEYINPUT58), .A3(G475), .ZN(new_n962));
  INV_X1    g776(.A(new_n371), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n962), .A2(new_n963), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n964), .A2(new_n965), .A3(new_n950), .ZN(G60));
  INV_X1    g780(.A(KEYINPUT124), .ZN(new_n967));
  NAND2_X1  g781(.A1(G478), .A2(G902), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT59), .Z(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n879), .B2(new_n926), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n647), .A2(new_n648), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n967), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n971), .A2(new_n969), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n950), .B1(new_n955), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  NOR3_X1   g790(.A1(new_n970), .A2(new_n967), .A3(new_n972), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n976), .A2(new_n977), .ZN(G63));
  AND2_X1   g792(.A1(new_n677), .A2(new_n678), .ZN(new_n979));
  NAND2_X1  g793(.A1(G217), .A2(G902), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT60), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(KEYINPUT126), .B1(new_n925), .B2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT126), .ZN(new_n984));
  AOI211_X1 g798(.A(new_n984), .B(new_n981), .C1(new_n861), .C2(new_n875), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n979), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  NOR4_X1   g800(.A1(new_n860), .A2(new_n862), .A3(new_n872), .A4(new_n834), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n982), .B1(new_n877), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n984), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n925), .A2(KEYINPUT126), .A3(new_n982), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n989), .A2(new_n622), .A3(new_n990), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n986), .A2(new_n991), .A3(new_n951), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT125), .ZN(new_n993));
  XNOR2_X1  g807(.A(KEYINPUT127), .B(KEYINPUT61), .ZN(new_n994));
  AND3_X1   g808(.A1(new_n992), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n994), .B1(new_n992), .B2(new_n993), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n995), .A2(new_n996), .ZN(G66));
  INV_X1    g811(.A(G224), .ZN(new_n998));
  OAI21_X1  g812(.A(G953), .B1(new_n426), .B2(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(new_n872), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n999), .B1(new_n1000), .B2(G953), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n943), .B1(G898), .B2(new_n283), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1001), .B(new_n1002), .ZN(G69));
  NAND2_X1  g817(.A1(new_n539), .A2(new_n548), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n550), .A2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(new_n363), .ZN(new_n1006));
  NAND2_X1  g820(.A1(G900), .A2(G953), .ZN(new_n1007));
  AND2_X1   g821(.A1(new_n831), .A2(new_n826), .ZN(new_n1008));
  AND2_X1   g822(.A1(new_n857), .A2(new_n779), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n823), .A2(new_n737), .A3(new_n711), .A4(new_n774), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n1008), .A2(new_n835), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n1006), .B(new_n1007), .C1(new_n1011), .C2(G953), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1009), .A2(new_n729), .ZN(new_n1013));
  XOR2_X1   g827(.A(new_n1013), .B(KEYINPUT62), .Z(new_n1014));
  NOR2_X1   g828(.A1(new_n712), .A2(new_n824), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n839), .A2(new_n868), .A3(new_n1015), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1014), .A2(new_n1008), .A3(new_n1016), .ZN(new_n1017));
  AND2_X1   g831(.A1(new_n1017), .A2(new_n283), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1012), .B1(new_n1018), .B2(new_n1006), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n283), .B1(G227), .B2(G900), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1019), .B(new_n1020), .ZN(G72));
  NOR2_X1   g835(.A1(new_n876), .A2(new_n878), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n715), .A2(new_n545), .ZN(new_n1023));
  NAND2_X1  g837(.A1(G472), .A2(G902), .ZN(new_n1024));
  XOR2_X1   g838(.A(new_n1024), .B(KEYINPUT63), .Z(new_n1025));
  NAND2_X1  g839(.A1(new_n716), .A2(new_n1025), .ZN(new_n1026));
  NOR3_X1   g840(.A1(new_n1022), .A2(new_n1023), .A3(new_n1026), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1025), .B1(new_n1011), .B2(new_n872), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1028), .A2(new_n1023), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1029), .A2(new_n951), .ZN(new_n1030));
  INV_X1    g844(.A(new_n716), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n1025), .B1(new_n1017), .B2(new_n872), .ZN(new_n1032));
  AOI211_X1 g846(.A(new_n1027), .B(new_n1030), .C1(new_n1031), .C2(new_n1032), .ZN(G57));
endmodule


