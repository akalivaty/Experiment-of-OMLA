//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 1 1 0 1 1 1 0 1 0 1 0 1 0 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1244, new_n1245, new_n1246, new_n1247, new_n1249,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1310, new_n1311,
    new_n1312;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(KEYINPUT64), .ZN(new_n212));
  INV_X1    g0012(.A(KEYINPUT64), .ZN(new_n213));
  NAND3_X1  g0013(.A1(new_n213), .A2(G1), .A3(G13), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G20), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n202), .A2(new_n203), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G50), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n219));
  INV_X1    g0019(.A(G232), .ZN(new_n220));
  INV_X1    g0020(.A(G97), .ZN(new_n221));
  INV_X1    g0021(.A(G257), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n219), .B1(new_n202), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n207), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n210), .B1(new_n216), .B2(new_n218), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G226), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G97), .B(G107), .Z(new_n239));
  XNOR2_X1  g0039(.A(G87), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n201), .A2(G68), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n203), .A2(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n241), .B(new_n246), .ZN(G351));
  XNOR2_X1  g0047(.A(KEYINPUT3), .B(G33), .ZN(new_n248));
  INV_X1    g0048(.A(G1698), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n248), .A2(G222), .A3(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G77), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n248), .A2(G1698), .ZN(new_n252));
  INV_X1    g0052(.A(G223), .ZN(new_n253));
  OAI221_X1 g0053(.A(new_n250), .B1(new_n251), .B2(new_n248), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  AND2_X1   g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n255), .B1(new_n212), .B2(new_n214), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G41), .ZN(new_n258));
  INV_X1    g0058(.A(G45), .ZN(new_n259));
  AOI21_X1  g0059(.A(G1), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G41), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G1), .A3(G13), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n260), .A2(new_n262), .A3(G274), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n265), .B1(G41), .B2(G45), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n262), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n264), .B1(G226), .B2(new_n268), .ZN(new_n269));
  AND2_X1   g0069(.A1(new_n257), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G190), .ZN(new_n271));
  INV_X1    g0071(.A(G200), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n204), .A2(G20), .ZN(new_n273));
  NOR2_X1   g0073(.A1(G20), .A2(G33), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n273), .A2(KEYINPUT67), .B1(G150), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT8), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n202), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT66), .B(G58), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n277), .B1(new_n278), .B2(new_n276), .ZN(new_n279));
  INV_X1    g0079(.A(G20), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G33), .ZN(new_n281));
  OAI221_X1 g0081(.A(new_n275), .B1(KEYINPUT67), .B2(new_n273), .C1(new_n279), .C2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n212), .A2(new_n214), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n265), .A2(G13), .A3(G20), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n212), .A2(new_n214), .A3(new_n286), .A4(new_n283), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n265), .A2(G20), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NOR3_X1   g0089(.A1(new_n287), .A2(new_n201), .A3(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n286), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n290), .B1(new_n201), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n285), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  OAI221_X1 g0094(.A(new_n271), .B1(new_n272), .B2(new_n270), .C1(new_n294), .C2(KEYINPUT9), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT10), .ZN(new_n297));
  AND3_X1   g0097(.A1(new_n285), .A2(KEYINPUT9), .A3(new_n292), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n298), .B(KEYINPUT70), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n296), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT70), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n298), .B(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT10), .B1(new_n302), .B2(new_n295), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n248), .A2(G232), .A3(G1698), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n248), .A2(G226), .A3(new_n249), .ZN(new_n306));
  NAND2_X1  g0106(.A1(G33), .A2(G97), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n256), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n264), .B1(G238), .B2(new_n268), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT13), .ZN(new_n311));
  AND3_X1   g0111(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n311), .B1(new_n309), .B2(new_n310), .ZN(new_n313));
  OAI21_X1  g0113(.A(G200), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n309), .A2(new_n310), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT13), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(G190), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n274), .ZN(new_n319));
  OAI22_X1  g0119(.A1(new_n319), .A2(new_n201), .B1(new_n280), .B2(G68), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n281), .A2(new_n251), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n284), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  XOR2_X1   g0122(.A(new_n322), .B(KEYINPUT11), .Z(new_n323));
  OAI22_X1  g0123(.A1(new_n286), .A2(G68), .B1(KEYINPUT71), .B2(KEYINPUT12), .ZN(new_n324));
  NAND2_X1  g0124(.A1(KEYINPUT71), .A2(KEYINPUT12), .ZN(new_n325));
  XNOR2_X1  g0125(.A(new_n324), .B(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n287), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n327), .A2(G68), .A3(new_n288), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n323), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n314), .A2(new_n318), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n312), .A2(new_n313), .ZN(new_n333));
  INV_X1    g0133(.A(G169), .ZN(new_n334));
  OAI21_X1  g0134(.A(KEYINPUT14), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(G179), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT14), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n337), .B(G169), .C1(new_n312), .C2(new_n313), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n335), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n330), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n332), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G179), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n270), .A2(new_n342), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n343), .B(new_n293), .C1(G169), .C2(new_n270), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n248), .A2(G232), .A3(new_n249), .ZN(new_n345));
  INV_X1    g0145(.A(G33), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(KEYINPUT3), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT3), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(G33), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(G107), .ZN(new_n351));
  INV_X1    g0151(.A(G238), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n345), .B(new_n351), .C1(new_n252), .C2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n256), .ZN(new_n354));
  INV_X1    g0154(.A(G244), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n263), .B1(new_n355), .B2(new_n267), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(G200), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n288), .A2(G77), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n287), .A2(new_n360), .ZN(new_n361));
  XNOR2_X1  g0161(.A(new_n361), .B(KEYINPUT68), .ZN(new_n362));
  NAND2_X1  g0162(.A1(G20), .A2(G77), .ZN(new_n363));
  XNOR2_X1  g0163(.A(KEYINPUT15), .B(G87), .ZN(new_n364));
  XNOR2_X1  g0164(.A(KEYINPUT8), .B(G58), .ZN(new_n365));
  OAI221_X1 g0165(.A(new_n363), .B1(new_n364), .B2(new_n281), .C1(new_n319), .C2(new_n365), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n366), .A2(new_n284), .B1(new_n251), .B2(new_n291), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n356), .B1(new_n353), .B2(new_n256), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(G190), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n359), .A2(new_n362), .A3(new_n367), .A4(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n358), .A2(new_n334), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n362), .A2(new_n367), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n368), .A2(new_n342), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n375), .B(KEYINPUT69), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n304), .A2(new_n341), .A3(new_n344), .A4(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT7), .B1(new_n350), .B2(new_n280), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT7), .ZN(new_n379));
  AOI211_X1 g0179(.A(new_n379), .B(G20), .C1(new_n347), .C2(new_n349), .ZN(new_n380));
  OAI21_X1  g0180(.A(G68), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n217), .B1(new_n278), .B2(new_n203), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n382), .A2(G20), .B1(G159), .B2(new_n274), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n381), .A2(new_n383), .A3(KEYINPUT16), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT72), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n381), .A2(new_n383), .A3(KEYINPUT72), .A4(KEYINPUT16), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT16), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n381), .A2(KEYINPUT73), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n379), .B1(new_n248), .B2(G20), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n348), .A2(G33), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n346), .A2(KEYINPUT3), .ZN(new_n393));
  OAI211_X1 g0193(.A(KEYINPUT7), .B(new_n280), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n203), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT73), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n383), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n389), .B1(new_n390), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n388), .A2(new_n398), .A3(new_n284), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n279), .A2(new_n289), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n327), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n279), .A2(new_n291), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n399), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT18), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n263), .B1(new_n220), .B2(new_n267), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n248), .A2(G226), .A3(G1698), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n248), .A2(G223), .A3(new_n249), .ZN(new_n409));
  NAND2_X1  g0209(.A1(G33), .A2(G87), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT74), .ZN(new_n411));
  XNOR2_X1  g0211(.A(new_n410), .B(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n408), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n407), .B1(new_n413), .B2(new_n256), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n414), .A2(new_n334), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n415), .B1(G179), .B2(new_n414), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n405), .A2(new_n406), .A3(new_n417), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n212), .A2(new_n214), .A3(new_n283), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n419), .B1(new_n386), .B2(new_n387), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n403), .B1(new_n420), .B2(new_n398), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT18), .B1(new_n421), .B2(new_n416), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT75), .ZN(new_n424));
  INV_X1    g0224(.A(G190), .ZN(new_n425));
  AND3_X1   g0225(.A1(new_n414), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  OR2_X1    g0226(.A1(new_n414), .A2(G200), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n424), .B1(new_n414), .B2(new_n425), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n399), .A2(new_n429), .A3(new_n404), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT17), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n421), .A2(KEYINPUT17), .A3(new_n429), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  OR2_X1    g0234(.A1(new_n423), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n265), .A2(G33), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n419), .A2(G116), .A3(new_n286), .A4(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(G116), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n291), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(G20), .B1(G33), .B2(G283), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n346), .A2(G97), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n440), .A2(new_n441), .B1(G20), .B2(new_n438), .ZN(new_n442));
  AND3_X1   g0242(.A1(new_n442), .A2(new_n284), .A3(KEYINPUT20), .ZN(new_n443));
  AOI21_X1  g0243(.A(KEYINPUT20), .B1(new_n442), .B2(new_n284), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n437), .B(new_n439), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n347), .A2(new_n349), .A3(G264), .A4(G1698), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n347), .A2(new_n349), .A3(G257), .A4(new_n249), .ZN(new_n447));
  XOR2_X1   g0247(.A(KEYINPUT79), .B(G303), .Z(new_n448));
  OAI211_X1 g0248(.A(new_n446), .B(new_n447), .C1(new_n448), .C2(new_n248), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n256), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n259), .A2(G1), .ZN(new_n451));
  NAND2_X1  g0251(.A1(KEYINPUT5), .A2(G41), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(KEYINPUT5), .A2(G41), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n451), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(G274), .B1(new_n255), .B2(new_n211), .ZN(new_n456));
  OAI21_X1  g0256(.A(KEYINPUT77), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n265), .A2(G45), .ZN(new_n458));
  OR2_X1    g0258(.A1(KEYINPUT5), .A2(G41), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n458), .B1(new_n459), .B2(new_n452), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT77), .ZN(new_n461));
  INV_X1    g0261(.A(G274), .ZN(new_n462));
  AND2_X1   g0262(.A1(G1), .A2(G13), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n462), .B1(new_n463), .B2(new_n261), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n460), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n457), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n459), .A2(new_n452), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n467), .A2(new_n451), .B1(new_n463), .B2(new_n261), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G270), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n450), .A2(new_n466), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n445), .B1(new_n470), .B2(G200), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n457), .A2(new_n465), .B1(new_n468), .B2(G270), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n472), .A2(G190), .A3(new_n450), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n470), .A2(G169), .A3(new_n445), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT21), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n445), .A2(G179), .A3(new_n450), .A4(new_n472), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n470), .A2(new_n445), .A3(KEYINPUT21), .A4(G169), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n474), .A2(new_n477), .A3(new_n478), .A4(new_n479), .ZN(new_n480));
  XNOR2_X1  g0280(.A(new_n480), .B(KEYINPUT80), .ZN(new_n481));
  INV_X1    g0281(.A(G250), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(new_n259), .B2(G1), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n265), .A2(new_n462), .A3(G45), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n262), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n352), .A2(new_n249), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n355), .A2(G1698), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n347), .A2(new_n486), .A3(new_n349), .A4(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n346), .A2(new_n438), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  AOI211_X1 g0291(.A(G179), .B(new_n485), .C1(new_n491), .C2(new_n256), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n256), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n262), .A2(new_n483), .A3(new_n484), .ZN(new_n494));
  AOI21_X1  g0294(.A(G169), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n347), .A2(new_n349), .A3(new_n280), .A4(G68), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT19), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(new_n281), .B2(new_n221), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g0300(.A(KEYINPUT78), .B(G87), .ZN(new_n501));
  NOR2_X1   g0301(.A1(G97), .A2(G107), .ZN(new_n502));
  NAND3_X1  g0302(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n501), .A2(new_n502), .B1(new_n280), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n284), .B1(new_n500), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n364), .A2(new_n291), .ZN(new_n506));
  INV_X1    g0306(.A(new_n364), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n327), .A2(new_n507), .A3(new_n436), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n505), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n327), .A2(G87), .A3(new_n436), .ZN(new_n510));
  AND3_X1   g0310(.A1(new_n505), .A2(new_n506), .A3(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(G238), .A2(G1698), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n512), .B1(new_n355), .B2(G1698), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n489), .B1(new_n513), .B2(new_n248), .ZN(new_n514));
  INV_X1    g0314(.A(new_n256), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n425), .B(new_n494), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n485), .B1(new_n491), .B2(new_n256), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n516), .B1(new_n517), .B2(G200), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n496), .A2(new_n509), .B1(new_n511), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n327), .A2(G97), .A3(new_n436), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n265), .A2(new_n221), .A3(G13), .A4(G20), .ZN(new_n521));
  OR2_X1    g0321(.A1(new_n521), .A2(KEYINPUT76), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(KEYINPUT76), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(G107), .B1(new_n378), .B2(new_n380), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT6), .ZN(new_n527));
  AND2_X1   g0327(.A1(G97), .A2(G107), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n527), .B1(new_n528), .B2(new_n502), .ZN(new_n529));
  INV_X1    g0329(.A(G107), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n530), .A2(KEYINPUT6), .A3(G97), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n532), .A2(G20), .B1(G77), .B2(new_n274), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n526), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n525), .B1(new_n534), .B2(new_n284), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n457), .A2(new_n465), .B1(new_n468), .B2(G257), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n347), .A2(new_n349), .A3(G244), .A4(new_n249), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT4), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(G250), .A2(G1698), .ZN(new_n540));
  NAND2_X1  g0340(.A1(KEYINPUT4), .A2(G244), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n540), .B1(new_n541), .B2(G1698), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n248), .A2(new_n542), .B1(G33), .B2(G283), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n256), .ZN(new_n545));
  AND3_X1   g0345(.A1(new_n536), .A2(new_n545), .A3(new_n425), .ZN(new_n546));
  AOI21_X1  g0346(.A(G200), .B1(new_n536), .B2(new_n545), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n535), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n530), .A2(KEYINPUT6), .A3(G97), .ZN(new_n549));
  XNOR2_X1  g0349(.A(G97), .B(G107), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n549), .B1(new_n550), .B2(new_n527), .ZN(new_n551));
  OAI22_X1  g0351(.A1(new_n551), .A2(new_n280), .B1(new_n251), .B2(new_n319), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n530), .B1(new_n391), .B2(new_n394), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n284), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n520), .A2(new_n524), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR3_X1   g0356(.A1(new_n455), .A2(new_n456), .A3(KEYINPUT77), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n461), .B1(new_n460), .B2(new_n464), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n455), .A2(new_n262), .ZN(new_n559));
  OAI22_X1  g0359(.A1(new_n557), .A2(new_n558), .B1(new_n222), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n515), .B1(new_n539), .B2(new_n543), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n334), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n536), .A2(new_n545), .A3(new_n342), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n556), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n519), .A2(new_n548), .A3(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n347), .A2(new_n349), .A3(new_n280), .A4(G87), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT22), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT22), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n248), .A2(new_n568), .A3(new_n280), .A4(G87), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT24), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n281), .A2(new_n438), .ZN(new_n572));
  OAI21_X1  g0372(.A(KEYINPUT81), .B1(new_n280), .B2(G107), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT23), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT23), .ZN(new_n575));
  OAI211_X1 g0375(.A(KEYINPUT81), .B(new_n575), .C1(new_n280), .C2(G107), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n572), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n570), .A2(new_n571), .A3(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n571), .B1(new_n570), .B2(new_n577), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n284), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n287), .B1(new_n265), .B2(G33), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT25), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n286), .B2(G107), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n291), .A2(KEYINPUT25), .A3(new_n530), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n582), .A2(G107), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n222), .A2(G1698), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(G250), .B2(G1698), .ZN(new_n588));
  INV_X1    g0388(.A(G294), .ZN(new_n589));
  OAI22_X1  g0389(.A1(new_n588), .A2(new_n350), .B1(new_n346), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n256), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n455), .A2(G264), .A3(new_n262), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n466), .A2(new_n591), .A3(new_n425), .A4(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n466), .A2(new_n591), .A3(new_n592), .ZN(new_n594));
  AOI22_X1  g0394(.A1(KEYINPUT83), .A2(new_n593), .B1(new_n594), .B2(new_n272), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n594), .A2(KEYINPUT83), .A3(new_n272), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n581), .B(new_n586), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT82), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n557), .A2(new_n558), .ZN(new_n599));
  NOR2_X1   g0399(.A1(G250), .A2(G1698), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n600), .B1(new_n222), .B2(G1698), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n601), .A2(new_n248), .B1(G33), .B2(G294), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n592), .B1(new_n602), .B2(new_n515), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n598), .B(G169), .C1(new_n599), .C2(new_n603), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n590), .A2(new_n256), .B1(new_n468), .B2(G264), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n605), .A2(G179), .A3(new_n466), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n598), .B1(new_n594), .B2(G169), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n570), .A2(new_n577), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(KEYINPUT24), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n419), .B1(new_n610), .B2(new_n578), .ZN(new_n611));
  INV_X1    g0411(.A(new_n586), .ZN(new_n612));
  OAI22_X1  g0412(.A1(new_n607), .A2(new_n608), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT84), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n597), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n614), .B1(new_n597), .B2(new_n613), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n565), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NOR4_X1   g0417(.A1(new_n377), .A2(new_n435), .A3(new_n481), .A4(new_n617), .ZN(G372));
  NAND2_X1  g0418(.A1(new_n316), .A2(new_n317), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n338), .B1(new_n342), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n337), .B1(new_n619), .B2(G169), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n340), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OR2_X1    g0422(.A1(new_n332), .A2(new_n374), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n434), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n304), .B1(new_n624), .B2(new_n423), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n625), .A2(new_n344), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n377), .A2(new_n435), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n479), .A2(new_n478), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n334), .B1(new_n472), .B2(new_n450), .ZN(new_n630));
  AOI21_X1  g0430(.A(KEYINPUT21), .B1(new_n630), .B2(new_n445), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n613), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n633), .A2(new_n565), .A3(new_n597), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n556), .A2(new_n562), .A3(new_n563), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n519), .ZN(new_n636));
  NOR2_X1   g0436(.A1(KEYINPUT85), .A2(KEYINPUT26), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n636), .A2(new_n637), .B1(new_n509), .B2(new_n496), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT85), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT26), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n635), .A2(new_n519), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n511), .A2(new_n518), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n494), .B1(new_n514), .B2(new_n515), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n334), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n517), .A2(new_n342), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n509), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(KEYINPUT26), .B1(new_n648), .B2(new_n564), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n640), .B1(new_n642), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n639), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n626), .B1(new_n628), .B2(new_n651), .ZN(G369));
  INV_X1    g0452(.A(new_n632), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n265), .A2(new_n280), .A3(G13), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(G213), .A3(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(G343), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n445), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n660), .B(KEYINPUT86), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n653), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n481), .B2(new_n661), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(G330), .ZN(new_n664));
  INV_X1    g0464(.A(new_n659), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n613), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n616), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n597), .A2(new_n613), .A3(new_n614), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n659), .B1(new_n611), .B2(new_n612), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n666), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n664), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n669), .A2(new_n653), .A3(new_n665), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n613), .A2(new_n659), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n673), .A2(new_n676), .ZN(G399));
  INV_X1    g0477(.A(new_n208), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(G41), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n501), .A2(new_n438), .A3(new_n502), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n679), .A2(new_n680), .A3(new_n265), .ZN(new_n681));
  INV_X1    g0481(.A(new_n218), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n681), .B1(new_n682), .B2(new_n679), .ZN(new_n683));
  XOR2_X1   g0483(.A(new_n683), .B(KEYINPUT87), .Z(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT28), .ZN(new_n685));
  AND4_X1   g0485(.A1(new_n605), .A2(new_n536), .A3(new_n545), .A4(new_n517), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT30), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n472), .A2(G179), .A3(new_n450), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n686), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n605), .A2(new_n536), .A3(new_n545), .A4(new_n517), .ZN(new_n691));
  OAI21_X1  g0491(.A(KEYINPUT30), .B1(new_n691), .B2(new_n688), .ZN(new_n692));
  AND4_X1   g0492(.A1(new_n342), .A2(new_n470), .A3(new_n594), .A4(new_n644), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n536), .A2(new_n545), .ZN(new_n694));
  AOI22_X1  g0494(.A1(new_n690), .A2(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT31), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n695), .A2(new_n696), .A3(new_n665), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n690), .A2(new_n692), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n693), .A2(new_n694), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(KEYINPUT88), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT88), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n695), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n701), .A2(new_n703), .A3(new_n659), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n697), .B1(new_n704), .B2(new_n696), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(KEYINPUT89), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT89), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n665), .B1(new_n700), .B2(KEYINPUT88), .ZN(new_n708));
  AOI21_X1  g0508(.A(KEYINPUT31), .B1(new_n708), .B2(new_n703), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n707), .B1(new_n709), .B2(new_n697), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT80), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n480), .B(new_n711), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n669), .A2(new_n712), .A3(new_n565), .A4(new_n665), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n706), .A2(new_n710), .A3(new_n713), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n714), .A2(G330), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT91), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n642), .A2(new_n649), .A3(new_n647), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n634), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n716), .B1(new_n718), .B2(new_n665), .ZN(new_n719));
  AOI211_X1 g0519(.A(KEYINPUT91), .B(new_n659), .C1(new_n717), .C2(new_n634), .ZN(new_n720));
  OAI21_X1  g0520(.A(KEYINPUT29), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n665), .B1(new_n639), .B2(new_n650), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(KEYINPUT90), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT29), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT90), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n724), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n715), .B1(new_n721), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n685), .B1(new_n729), .B2(G1), .ZN(G364));
  NOR2_X1   g0530(.A1(new_n280), .A2(new_n342), .ZN(new_n731));
  NOR2_X1   g0531(.A1(G190), .A2(G200), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(G311), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n280), .A2(G179), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n732), .ZN(new_n736));
  INV_X1    g0536(.A(G329), .ZN(new_n737));
  OAI22_X1  g0537(.A1(new_n733), .A2(new_n734), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n731), .A2(G190), .A3(new_n272), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  AOI211_X1 g0540(.A(new_n248), .B(new_n738), .C1(G322), .C2(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n735), .A2(new_n425), .A3(G200), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT95), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G283), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n731), .A2(G200), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n425), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(G190), .ZN(new_n747));
  XNOR2_X1  g0547(.A(KEYINPUT33), .B(G317), .ZN(new_n748));
  AOI22_X1  g0548(.A1(G326), .A2(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n425), .A2(G179), .A3(G200), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n280), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n735), .A2(G190), .A3(G200), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n752), .A2(G294), .B1(new_n754), .B2(G303), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n741), .A2(new_n744), .A3(new_n749), .A4(new_n755), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n739), .A2(new_n278), .B1(new_n733), .B2(new_n251), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n757), .B1(G50), .B2(new_n746), .ZN(new_n758));
  XOR2_X1   g0558(.A(new_n758), .B(KEYINPUT94), .Z(new_n759));
  NAND2_X1  g0559(.A1(new_n743), .A2(G107), .ZN(new_n760));
  OAI211_X1 g0560(.A(new_n760), .B(new_n248), .C1(new_n501), .C2(new_n753), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT96), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G159), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n736), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT32), .ZN(new_n766));
  AOI22_X1  g0566(.A1(G97), .A2(new_n752), .B1(new_n747), .B2(G68), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n759), .A2(new_n763), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n761), .A2(new_n762), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n756), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n215), .B1(new_n280), .B2(G169), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT93), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G13), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(G20), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G45), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT92), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n779), .A2(new_n265), .A3(new_n679), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G13), .A2(G33), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G20), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n773), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n678), .A2(new_n350), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n786), .A2(G355), .B1(new_n438), .B2(new_n678), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n246), .A2(new_n259), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n678), .A2(new_n248), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n789), .B1(G45), .B2(new_n218), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n787), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n781), .B1(new_n785), .B2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n784), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n774), .B(new_n792), .C1(new_n663), .C2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n664), .A2(new_n781), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n663), .A2(G330), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(G396));
  NAND2_X1  g0597(.A1(new_n372), .A2(new_n659), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n370), .A2(new_n374), .A3(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(KEYINPUT99), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n374), .A2(new_n665), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n370), .A2(new_n374), .A3(KEYINPUT99), .A4(new_n798), .ZN(new_n803));
  AND3_X1   g0603(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n724), .A2(new_n727), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n801), .A2(new_n803), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n723), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n715), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n780), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n715), .A2(new_n805), .A3(new_n807), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n739), .A2(new_n589), .B1(new_n736), .B2(new_n734), .ZN(new_n812));
  INV_X1    g0612(.A(new_n733), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n248), .B(new_n812), .C1(G116), .C2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n743), .A2(G87), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n752), .A2(G97), .B1(new_n754), .B2(G107), .ZN(new_n816));
  AOI22_X1  g0616(.A1(G283), .A2(new_n747), .B1(new_n746), .B2(G303), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n814), .A2(new_n815), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  XOR2_X1   g0618(.A(new_n818), .B(KEYINPUT97), .Z(new_n819));
  XOR2_X1   g0619(.A(KEYINPUT98), .B(G143), .Z(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n740), .A2(new_n821), .B1(new_n813), .B2(G159), .ZN(new_n822));
  INV_X1    g0622(.A(new_n747), .ZN(new_n823));
  INV_X1    g0623(.A(G150), .ZN(new_n824));
  INV_X1    g0624(.A(G137), .ZN(new_n825));
  INV_X1    g0625(.A(new_n746), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n822), .B1(new_n823), .B2(new_n824), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT34), .ZN(new_n828));
  OR2_X1    g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n827), .A2(new_n828), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n743), .A2(G68), .ZN(new_n831));
  INV_X1    g0631(.A(G132), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n248), .B1(new_n736), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n751), .A2(new_n278), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n833), .B(new_n834), .C1(G50), .C2(new_n754), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n829), .A2(new_n830), .A3(new_n831), .A4(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n772), .B1(new_n819), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n773), .A2(new_n782), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n781), .B(new_n837), .C1(new_n251), .C2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n804), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n839), .B1(new_n783), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n811), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(G384));
  NOR2_X1   g0643(.A1(new_n776), .A2(new_n265), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n340), .A2(new_n659), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n622), .A2(new_n331), .A3(new_n845), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n340), .B(new_n659), .C1(new_n339), .C2(new_n332), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(new_n840), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n659), .B1(new_n695), .B2(new_n702), .ZN(new_n850));
  AND3_X1   g0650(.A1(new_n698), .A2(new_n702), .A3(new_n699), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n696), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n701), .A2(new_n703), .A3(KEYINPUT31), .A4(new_n659), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n849), .B1(new_n854), .B2(new_n713), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n381), .A2(new_n383), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n389), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n403), .B1(new_n420), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n430), .B1(new_n657), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n858), .A2(new_n416), .ZN(new_n860));
  OAI21_X1  g0660(.A(KEYINPUT37), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n405), .A2(new_n417), .ZN(new_n862));
  INV_X1    g0662(.A(new_n657), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n405), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT37), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n862), .A2(new_n864), .A3(new_n865), .A4(new_n430), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n861), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n858), .A2(new_n657), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n423), .B2(new_n434), .ZN(new_n869));
  AND3_X1   g0669(.A1(new_n867), .A2(new_n869), .A3(KEYINPUT38), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n862), .A2(new_n864), .A3(new_n430), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT37), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n866), .ZN(new_n873));
  INV_X1    g0673(.A(new_n864), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n423), .B2(new_n434), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT38), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n855), .B(KEYINPUT40), .C1(new_n870), .C2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n804), .B1(new_n846), .B2(new_n847), .ZN(new_n879));
  NOR3_X1   g0679(.A1(new_n617), .A2(new_n481), .A3(new_n659), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n852), .A2(new_n853), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n867), .A2(new_n869), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT38), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n867), .A2(new_n869), .A3(KEYINPUT38), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n882), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT102), .B1(new_n887), .B2(KEYINPUT40), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT38), .B1(new_n867), .B2(new_n869), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n855), .B1(new_n870), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT102), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT40), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n878), .B1(new_n888), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n854), .A2(new_n713), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n627), .A2(new_n895), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n894), .A2(new_n896), .ZN(new_n898));
  INV_X1    g0698(.A(G330), .ZN(new_n899));
  NOR3_X1   g0699(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  OR2_X1    g0701(.A1(new_n374), .A2(new_n659), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n902), .B(KEYINPUT101), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n723), .B2(new_n806), .ZN(new_n905));
  INV_X1    g0705(.A(new_n848), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n885), .A2(new_n886), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n907), .A2(new_n908), .B1(new_n423), .B2(new_n657), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT39), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n910), .B1(new_n870), .B2(new_n876), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n885), .A2(KEYINPUT39), .A3(new_n886), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n339), .A2(new_n340), .A3(new_n665), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n909), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n728), .A2(new_n627), .A3(new_n721), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n626), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n916), .B(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n844), .B1(new_n901), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n919), .B2(new_n901), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n532), .A2(KEYINPUT35), .ZN(new_n922));
  NOR3_X1   g0722(.A1(new_n922), .A2(new_n438), .A3(new_n216), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n924), .A2(KEYINPUT100), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n532), .A2(KEYINPUT35), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(KEYINPUT100), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT36), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n682), .B(G77), .C1(new_n203), .C2(new_n278), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n242), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n931), .A2(G1), .A3(new_n775), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n921), .A2(new_n929), .A3(new_n932), .ZN(G367));
  OAI22_X1  g0733(.A1(new_n823), .A2(new_n589), .B1(new_n742), .B2(new_n221), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n826), .A2(new_n734), .B1(new_n530), .B2(new_n751), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(G283), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n739), .A2(new_n448), .B1(new_n733), .B2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n736), .ZN(new_n939));
  AOI211_X1 g0739(.A(new_n248), .B(new_n938), .C1(G317), .C2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n754), .A2(KEYINPUT46), .A3(G116), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT46), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n753), .B2(new_n438), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n936), .A2(new_n940), .A3(new_n941), .A4(new_n943), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n753), .A2(new_n278), .B1(new_n736), .B2(new_n825), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT108), .Z(new_n946));
  OAI21_X1  g0746(.A(new_n248), .B1(new_n742), .B2(new_n251), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n947), .B(KEYINPUT107), .Z(new_n948));
  OAI22_X1  g0748(.A1(new_n739), .A2(new_n824), .B1(new_n733), .B2(new_n201), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(G159), .B2(new_n747), .ZN(new_n950));
  AOI22_X1  g0750(.A1(G68), .A2(new_n752), .B1(new_n746), .B2(new_n821), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n946), .A2(new_n948), .A3(new_n950), .A4(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n944), .A2(new_n952), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n953), .B(KEYINPUT109), .Z(new_n954));
  OR2_X1    g0754(.A1(new_n954), .A2(KEYINPUT47), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(KEYINPUT47), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n955), .A2(new_n773), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n519), .B1(new_n511), .B2(new_n665), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT104), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NOR3_X1   g0760(.A1(new_n647), .A2(new_n511), .A3(new_n665), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT103), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n958), .A2(new_n959), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n960), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n964), .A2(new_n793), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n237), .A2(new_n789), .B1(new_n678), .B2(new_n507), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n781), .B1(new_n785), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n957), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n779), .A2(new_n265), .ZN(new_n970));
  INV_X1    g0770(.A(new_n729), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n671), .B1(new_n632), .B2(new_n659), .ZN(new_n972));
  INV_X1    g0772(.A(new_n664), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n972), .B(new_n674), .C1(new_n973), .C2(KEYINPUT105), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(KEYINPUT105), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n974), .B(new_n975), .Z(new_n976));
  AND2_X1   g0776(.A1(new_n976), .A2(new_n729), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n548), .B(new_n564), .C1(new_n535), .C2(new_n665), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n635), .A2(new_n659), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n676), .A2(new_n980), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n981), .B(KEYINPUT45), .Z(new_n982));
  NOR2_X1   g0782(.A1(new_n676), .A2(new_n980), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT44), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n982), .A2(new_n673), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n982), .A2(new_n984), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n672), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n977), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(KEYINPUT106), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT106), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n977), .A2(new_n990), .A3(new_n985), .A4(new_n987), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n971), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n679), .B(KEYINPUT41), .Z(new_n993));
  OAI21_X1  g0793(.A(new_n970), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n980), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n674), .A2(new_n995), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n996), .A2(KEYINPUT42), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n564), .B1(new_n978), .B2(new_n613), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n996), .A2(KEYINPUT42), .B1(new_n665), .B2(new_n998), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n997), .A2(new_n999), .B1(KEYINPUT43), .B2(new_n964), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n672), .A2(new_n980), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1002), .B(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n969), .B1(new_n994), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(G387));
  INV_X1    g0806(.A(new_n789), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(new_n234), .B2(G45), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(new_n680), .B2(new_n786), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n365), .A2(G50), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT50), .Z(new_n1011));
  OAI21_X1  g0811(.A(new_n259), .B1(new_n203), .B2(new_n251), .ZN(new_n1012));
  NOR3_X1   g0812(.A1(new_n1011), .A2(new_n680), .A3(new_n1012), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n1009), .A2(new_n1013), .B1(G107), .B2(new_n208), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n781), .B1(new_n1014), .B2(new_n785), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n740), .A2(G50), .B1(new_n939), .B2(G150), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n350), .B1(new_n813), .B2(G68), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1016), .B(new_n1017), .C1(new_n279), .C2(new_n823), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n753), .A2(new_n251), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(new_n507), .B2(new_n752), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n764), .B2(new_n826), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n1018), .B(new_n1021), .C1(G97), .C2(new_n743), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n751), .A2(new_n937), .B1(new_n753), .B2(new_n589), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n448), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G317), .A2(new_n740), .B1(new_n1024), .B2(new_n813), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n746), .A2(G322), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1025), .B(new_n1026), .C1(new_n734), .C2(new_n823), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT48), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1023), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n1028), .B2(new_n1027), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT110), .Z(new_n1031));
  OR2_X1    g0831(.A1(new_n1031), .A2(KEYINPUT49), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n248), .B1(new_n939), .B2(G326), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n438), .B2(new_n742), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n1031), .B2(KEYINPUT49), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1022), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1015), .B1(new_n1036), .B2(new_n772), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n671), .B2(new_n784), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n970), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1038), .B1(new_n976), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n977), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n679), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n976), .A2(new_n729), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1040), .B1(new_n1042), .B2(new_n1043), .ZN(G393));
  INV_X1    g0844(.A(new_n785), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n241), .A2(new_n1007), .B1(new_n221), .B2(new_n208), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n780), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(G150), .A2(new_n746), .B1(new_n740), .B2(G159), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT112), .ZN(new_n1049));
  XOR2_X1   g0849(.A(KEYINPUT111), .B(KEYINPUT51), .Z(new_n1050));
  OR2_X1    g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n751), .A2(new_n251), .B1(new_n753), .B2(new_n203), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n248), .B1(new_n733), .B2(new_n365), .C1(new_n736), .C2(new_n820), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n1053), .B(new_n1054), .C1(G50), .C2(new_n747), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1051), .A2(new_n815), .A3(new_n1052), .A4(new_n1055), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G317), .A2(new_n746), .B1(new_n740), .B2(G311), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT52), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n823), .A2(new_n448), .B1(new_n753), .B2(new_n937), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(G116), .B2(new_n752), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n350), .B1(new_n733), .B2(new_n589), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(G322), .B2(new_n939), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1060), .A2(new_n760), .A3(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1056), .B1(new_n1058), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1047), .B1(new_n1064), .B2(new_n773), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n980), .B2(new_n793), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n987), .A2(new_n985), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1066), .B1(new_n1067), .B2(new_n970), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n989), .A2(new_n991), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n679), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n1041), .B2(new_n1067), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1068), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(G390));
  NAND3_X1  g0873(.A1(new_n642), .A2(new_n649), .A3(new_n647), .ZN(new_n1074));
  AND4_X1   g0874(.A1(new_n597), .A2(new_n519), .A3(new_n564), .A4(new_n548), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1074), .B1(new_n633), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(KEYINPUT91), .B1(new_n1076), .B2(new_n659), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n718), .A2(new_n716), .A3(new_n665), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n804), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(KEYINPUT113), .B1(new_n1079), .B2(new_n904), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n840), .B1(new_n719), .B2(new_n720), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT113), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1081), .A2(new_n1082), .A3(new_n903), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1080), .A2(new_n848), .A3(new_n1083), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n870), .A2(new_n876), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1085), .A2(new_n914), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n911), .A2(new_n912), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n913), .B1(new_n905), .B2(new_n906), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n899), .B1(new_n854), .B2(new_n713), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n879), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1091), .A2(KEYINPUT114), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT114), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1092), .A2(new_n1096), .A3(new_n879), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n715), .A2(new_n1097), .A3(new_n840), .A4(new_n848), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1087), .A2(new_n1090), .A3(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1095), .A2(new_n1039), .A3(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1088), .A2(new_n782), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n781), .B1(new_n838), .B2(new_n279), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT117), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n739), .A2(new_n438), .B1(new_n736), .B2(new_n589), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n248), .B(new_n1104), .C1(G97), .C2(new_n813), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G77), .A2(new_n752), .B1(new_n747), .B2(G107), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n746), .A2(G283), .B1(new_n754), .B2(G87), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1105), .A2(new_n831), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(KEYINPUT54), .B(G143), .ZN(new_n1109));
  INV_X1    g0909(.A(G125), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n733), .A2(new_n1109), .B1(new_n736), .B2(new_n1110), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n350), .B(new_n1111), .C1(G132), .C2(new_n740), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n753), .A2(new_n824), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT53), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(G159), .A2(new_n752), .B1(new_n747), .B2(G137), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n742), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n746), .A2(G128), .B1(new_n1116), .B2(G50), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1112), .A2(new_n1114), .A3(new_n1115), .A4(new_n1117), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n1108), .A2(new_n1118), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1101), .B(new_n1103), .C1(new_n772), .C2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1100), .A2(new_n1120), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n1084), .A2(new_n1086), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1094), .A2(KEYINPUT114), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1099), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n627), .A2(new_n1092), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n917), .A2(new_n626), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1092), .A2(new_n840), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n906), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n714), .A2(G330), .A3(new_n840), .A4(new_n848), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1083), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1082), .B1(new_n1081), .B2(new_n903), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1129), .B(new_n1130), .C1(new_n1131), .C2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n713), .B1(new_n705), .B2(KEYINPUT89), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n709), .A2(new_n707), .A3(new_n697), .ZN(new_n1136));
  OAI211_X1 g0936(.A(G330), .B(new_n840), .C1(new_n1135), .C2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n906), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n905), .B1(new_n1138), .B2(new_n1093), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1127), .B1(new_n1134), .B2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(KEYINPUT115), .B1(new_n1124), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1138), .A2(new_n1093), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n905), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1126), .B1(new_n1144), .B2(new_n1133), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT115), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1095), .A2(new_n1145), .A3(new_n1146), .A4(new_n1099), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1070), .B1(new_n1141), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1145), .B1(new_n1124), .B2(KEYINPUT116), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(KEYINPUT116), .B2(new_n1124), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1121), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(G378));
  XNOR2_X1  g0952(.A(new_n1126), .B(KEYINPUT121), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(new_n1141), .B2(new_n1147), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT57), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n304), .A2(new_n344), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT119), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1157), .B(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n293), .A2(new_n863), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT55), .ZN(new_n1161));
  OR2_X1    g0961(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1164));
  AND3_X1   g0964(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1163), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1166));
  OR2_X1    g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n887), .A2(KEYINPUT102), .A3(KEYINPUT40), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n891), .B1(new_n890), .B2(new_n892), .ZN(new_n1169));
  OAI211_X1 g0969(.A(G330), .B(new_n877), .C1(new_n1168), .C2(new_n1169), .ZN(new_n1170));
  AND2_X1   g0970(.A1(new_n909), .A2(new_n915), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n916), .B1(new_n894), .B2(G330), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1167), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n894), .A2(G330), .A3(new_n916), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1174), .A2(new_n1178), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n1155), .A2(new_n1156), .A3(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(KEYINPUT122), .B1(new_n1180), .B2(new_n1070), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1141), .A2(new_n1147), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n1153), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1179), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1183), .A2(KEYINPUT57), .A3(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT122), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1185), .A2(new_n1186), .A3(new_n679), .ZN(new_n1187));
  AOI21_X1  g0987(.A(KEYINPUT57), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1181), .A2(new_n1187), .A3(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1177), .A2(new_n783), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n350), .A2(new_n258), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n346), .A2(new_n258), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n1192), .A2(new_n201), .A3(new_n1193), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(G68), .A2(new_n752), .B1(new_n746), .B2(G116), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT118), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1192), .B1(new_n740), .B2(G107), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n507), .A2(new_n813), .B1(new_n939), .B2(G283), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n742), .A2(new_n278), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n1019), .B(new_n1199), .C1(G97), .C2(new_n747), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .A4(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1194), .B1(new_n1202), .B2(KEYINPUT58), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1193), .B1(new_n939), .B2(G124), .ZN(new_n1204));
  INV_X1    g1004(.A(G128), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n739), .A2(new_n1205), .B1(new_n733), .B2(new_n825), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n746), .A2(G125), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1207), .B1(new_n753), .B2(new_n1109), .C1(new_n823), .C2(new_n832), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1206), .B(new_n1208), .C1(G150), .C2(new_n752), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT59), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1204), .B1(new_n764), .B2(new_n742), .C1(new_n1209), .C2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1209), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1212), .A2(KEYINPUT59), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1203), .B1(KEYINPUT58), .B2(new_n1202), .C1(new_n1211), .C2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n773), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n781), .B1(new_n838), .B2(new_n201), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1191), .A2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n1184), .B2(new_n1039), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1190), .A2(new_n1219), .ZN(G375));
  AOI21_X1  g1020(.A(new_n970), .B1(new_n1144), .B2(new_n1133), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n906), .A2(new_n782), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(new_n773), .A2(G68), .A3(new_n782), .ZN(new_n1223));
  OR3_X1    g1023(.A1(new_n826), .A2(KEYINPUT123), .A3(new_n832), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n740), .A2(G137), .B1(new_n813), .B2(G150), .ZN(new_n1225));
  OAI21_X1  g1025(.A(KEYINPUT123), .B1(new_n826), .B2(new_n832), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n350), .B1(new_n939), .B2(G128), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1199), .B1(G159), .B2(new_n754), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1229), .B1(new_n201), .B2(new_n751), .C1(new_n823), .C2(new_n1109), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n743), .A2(G77), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(G116), .A2(new_n747), .B1(new_n746), .B2(G294), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n248), .B1(new_n939), .B2(G303), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n740), .A2(G283), .B1(new_n813), .B2(G107), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n752), .A2(new_n507), .B1(new_n754), .B2(G97), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1232), .A2(new_n1233), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n1228), .A2(new_n1230), .B1(new_n1231), .B2(new_n1236), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n781), .B(new_n1223), .C1(new_n1237), .C2(new_n773), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1221), .B1(new_n1222), .B2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n993), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1144), .A2(new_n1126), .A3(new_n1133), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1140), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1239), .A2(new_n1242), .ZN(G381));
  INV_X1    g1043(.A(G375), .ZN(new_n1244));
  OR2_X1    g1044(.A1(G393), .A2(G396), .ZN(new_n1245));
  NOR4_X1   g1045(.A1(G390), .A2(new_n1245), .A3(G384), .A4(G381), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1244), .A2(new_n1005), .A3(new_n1151), .A4(new_n1246), .ZN(new_n1247));
  XOR2_X1   g1047(.A(new_n1247), .B(KEYINPUT124), .Z(G407));
  NAND3_X1  g1048(.A1(new_n1244), .A2(new_n658), .A3(new_n1151), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(G407), .A2(G213), .A3(new_n1249), .ZN(G409));
  NAND2_X1  g1050(.A1(G387), .A2(new_n1072), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT126), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1005), .A2(G390), .ZN(new_n1253));
  XOR2_X1   g1053(.A(G393), .B(G396), .Z(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1251), .A2(new_n1252), .A3(new_n1253), .A4(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1252), .B1(new_n1005), .B2(G390), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1005), .A2(G390), .ZN(new_n1258));
  AOI211_X1 g1058(.A(new_n969), .B(new_n1072), .C1(new_n994), .C2(new_n1004), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n1257), .A2(new_n1254), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1256), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT127), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1190), .A2(G378), .A3(new_n1219), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT125), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1183), .A2(new_n1240), .A3(new_n1184), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n1219), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1265), .B1(new_n1267), .B2(new_n1151), .ZN(new_n1268));
  NOR3_X1   g1068(.A1(new_n1155), .A2(new_n993), .A3(new_n1179), .ZN(new_n1269));
  OAI22_X1  g1069(.A1(new_n1179), .A2(new_n970), .B1(new_n1191), .B2(new_n1217), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1265), .B(new_n1151), .C1(new_n1269), .C2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1268), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1264), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(G213), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1275), .A2(G343), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1274), .A2(new_n1277), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1140), .A2(KEYINPUT60), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1241), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1070), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1281), .B1(new_n1280), .B2(new_n1279), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1239), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n842), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1282), .A2(G384), .A3(new_n1239), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  AND3_X1   g1086(.A1(new_n1286), .A2(G2897), .A3(new_n1276), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1286), .B1(G2897), .B2(new_n1276), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1278), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT61), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1263), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1286), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1274), .A2(new_n1277), .A3(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(KEYINPUT62), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1276), .B1(new_n1264), .B2(new_n1273), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT62), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1296), .A2(new_n1297), .A3(new_n1293), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1295), .A2(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1262), .B1(new_n1292), .B2(new_n1299), .ZN(new_n1300));
  AND3_X1   g1100(.A1(new_n1296), .A2(KEYINPUT63), .A3(new_n1293), .ZN(new_n1301));
  AOI21_X1  g1101(.A(KEYINPUT63), .B1(new_n1296), .B2(new_n1293), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1261), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1256), .A2(new_n1260), .A3(KEYINPUT127), .ZN(new_n1304));
  OR2_X1    g1104(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1305));
  OAI211_X1 g1105(.A(new_n1304), .B(new_n1291), .C1(new_n1305), .C2(new_n1296), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1303), .A2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1300), .A2(new_n1308), .ZN(G405));
  NAND2_X1  g1109(.A1(G375), .A2(new_n1151), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(new_n1264), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(new_n1311), .B(new_n1293), .ZN(new_n1312));
  XNOR2_X1  g1112(.A(new_n1312), .B(new_n1262), .ZN(G402));
endmodule


