

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X1 U553 ( .A(n622), .Z(n669) );
  NOR2_X1 U554 ( .A1(n734), .A2(n733), .ZN(n518) );
  XOR2_X1 U555 ( .A(KEYINPUT29), .B(n654), .Z(n519) );
  INV_X1 U556 ( .A(KEYINPUT26), .ZN(n619) );
  NOR2_X1 U557 ( .A1(n643), .A2(n934), .ZN(n644) );
  XNOR2_X1 U558 ( .A(n592), .B(KEYINPUT64), .ZN(n622) );
  OR2_X1 U559 ( .A1(n668), .A2(n667), .ZN(n684) );
  XNOR2_X1 U560 ( .A(n523), .B(KEYINPUT68), .ZN(n532) );
  BUF_X1 U561 ( .A(n532), .Z(n891) );
  NOR2_X1 U562 ( .A1(G651), .A2(n584), .ZN(n803) );
  INV_X1 U563 ( .A(KEYINPUT69), .ZN(n528) );
  XNOR2_X1 U564 ( .A(n529), .B(n528), .ZN(n530) );
  NOR2_X1 U565 ( .A1(n531), .A2(n530), .ZN(G160) );
  NOR2_X1 U566 ( .A1(G2105), .A2(G2104), .ZN(n520) );
  XOR2_X1 U567 ( .A(KEYINPUT17), .B(n520), .Z(n890) );
  NAND2_X1 U568 ( .A1(G137), .A2(n890), .ZN(n522) );
  AND2_X1 U569 ( .A1(G2105), .A2(G2104), .ZN(n895) );
  NAND2_X1 U570 ( .A1(G113), .A2(n895), .ZN(n521) );
  NAND2_X1 U571 ( .A1(n522), .A2(n521), .ZN(n531) );
  XNOR2_X1 U572 ( .A(KEYINPUT67), .B(G2104), .ZN(n525) );
  NOR2_X1 U573 ( .A1(n525), .A2(G2105), .ZN(n523) );
  NAND2_X1 U574 ( .A1(G101), .A2(n532), .ZN(n524) );
  XOR2_X1 U575 ( .A(n524), .B(KEYINPUT23), .Z(n527) );
  AND2_X1 U576 ( .A1(n525), .A2(G2105), .ZN(n898) );
  NAND2_X1 U577 ( .A1(n898), .A2(G125), .ZN(n526) );
  NAND2_X1 U578 ( .A1(n527), .A2(n526), .ZN(n529) );
  NAND2_X1 U579 ( .A1(G102), .A2(n891), .ZN(n534) );
  NAND2_X1 U580 ( .A1(n890), .A2(G138), .ZN(n533) );
  NAND2_X1 U581 ( .A1(n534), .A2(n533), .ZN(n538) );
  NAND2_X1 U582 ( .A1(G114), .A2(n895), .ZN(n536) );
  NAND2_X1 U583 ( .A1(G126), .A2(n898), .ZN(n535) );
  NAND2_X1 U584 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U585 ( .A1(n538), .A2(n537), .ZN(G164) );
  XOR2_X1 U586 ( .A(G543), .B(KEYINPUT0), .Z(n584) );
  NAND2_X1 U587 ( .A1(n803), .A2(G52), .ZN(n542) );
  INV_X1 U588 ( .A(G651), .ZN(n543) );
  NOR2_X1 U589 ( .A1(G543), .A2(n543), .ZN(n539) );
  XOR2_X1 U590 ( .A(KEYINPUT1), .B(n539), .Z(n540) );
  XNOR2_X1 U591 ( .A(KEYINPUT70), .B(n540), .ZN(n804) );
  NAND2_X1 U592 ( .A1(G64), .A2(n804), .ZN(n541) );
  NAND2_X1 U593 ( .A1(n542), .A2(n541), .ZN(n550) );
  NOR2_X1 U594 ( .A1(n584), .A2(n543), .ZN(n807) );
  NAND2_X1 U595 ( .A1(n807), .A2(G77), .ZN(n546) );
  NOR2_X1 U596 ( .A1(G543), .A2(G651), .ZN(n544) );
  XNOR2_X1 U597 ( .A(n544), .B(KEYINPUT66), .ZN(n808) );
  NAND2_X1 U598 ( .A1(G90), .A2(n808), .ZN(n545) );
  NAND2_X1 U599 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U600 ( .A(KEYINPUT9), .B(n547), .ZN(n548) );
  XNOR2_X1 U601 ( .A(KEYINPUT73), .B(n548), .ZN(n549) );
  NOR2_X1 U602 ( .A1(n550), .A2(n549), .ZN(G171) );
  INV_X1 U603 ( .A(G171), .ZN(G301) );
  NAND2_X1 U604 ( .A1(n803), .A2(G51), .ZN(n552) );
  NAND2_X1 U605 ( .A1(G63), .A2(n804), .ZN(n551) );
  NAND2_X1 U606 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U607 ( .A(KEYINPUT6), .B(n553), .ZN(n560) );
  NAND2_X1 U608 ( .A1(n808), .A2(G89), .ZN(n554) );
  XOR2_X1 U609 ( .A(KEYINPUT81), .B(n554), .Z(n555) );
  XNOR2_X1 U610 ( .A(n555), .B(KEYINPUT4), .ZN(n557) );
  NAND2_X1 U611 ( .A1(G76), .A2(n807), .ZN(n556) );
  NAND2_X1 U612 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U613 ( .A(n558), .B(KEYINPUT5), .Z(n559) );
  NOR2_X1 U614 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U615 ( .A(KEYINPUT7), .B(n561), .Z(n562) );
  XNOR2_X1 U616 ( .A(KEYINPUT82), .B(n562), .ZN(G168) );
  NAND2_X1 U617 ( .A1(n807), .A2(G75), .ZN(n564) );
  NAND2_X1 U618 ( .A1(G88), .A2(n808), .ZN(n563) );
  NAND2_X1 U619 ( .A1(n564), .A2(n563), .ZN(n568) );
  NAND2_X1 U620 ( .A1(n803), .A2(G50), .ZN(n566) );
  NAND2_X1 U621 ( .A1(G62), .A2(n804), .ZN(n565) );
  NAND2_X1 U622 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U623 ( .A1(n568), .A2(n567), .ZN(G166) );
  INV_X1 U624 ( .A(G166), .ZN(G303) );
  XOR2_X1 U625 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U626 ( .A1(G86), .A2(n808), .ZN(n570) );
  NAND2_X1 U627 ( .A1(G61), .A2(n804), .ZN(n569) );
  NAND2_X1 U628 ( .A1(n570), .A2(n569), .ZN(n573) );
  NAND2_X1 U629 ( .A1(n807), .A2(G73), .ZN(n571) );
  XOR2_X1 U630 ( .A(KEYINPUT2), .B(n571), .Z(n572) );
  NOR2_X1 U631 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U632 ( .A1(n803), .A2(G48), .ZN(n574) );
  NAND2_X1 U633 ( .A1(n575), .A2(n574), .ZN(G305) );
  NAND2_X1 U634 ( .A1(n803), .A2(G47), .ZN(n576) );
  XNOR2_X1 U635 ( .A(n576), .B(KEYINPUT72), .ZN(n583) );
  NAND2_X1 U636 ( .A1(n807), .A2(G72), .ZN(n578) );
  NAND2_X1 U637 ( .A1(G85), .A2(n808), .ZN(n577) );
  NAND2_X1 U638 ( .A1(n578), .A2(n577), .ZN(n581) );
  NAND2_X1 U639 ( .A1(G60), .A2(n804), .ZN(n579) );
  XNOR2_X1 U640 ( .A(KEYINPUT71), .B(n579), .ZN(n580) );
  NOR2_X1 U641 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U642 ( .A1(n583), .A2(n582), .ZN(G290) );
  NAND2_X1 U643 ( .A1(G87), .A2(n584), .ZN(n586) );
  NAND2_X1 U644 ( .A1(G74), .A2(G651), .ZN(n585) );
  NAND2_X1 U645 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U646 ( .A1(n804), .A2(n587), .ZN(n589) );
  NAND2_X1 U647 ( .A1(n803), .A2(G49), .ZN(n588) );
  NAND2_X1 U648 ( .A1(n589), .A2(n588), .ZN(G288) );
  NAND2_X1 U649 ( .A1(G160), .A2(G40), .ZN(n693) );
  XNOR2_X1 U650 ( .A(n693), .B(KEYINPUT93), .ZN(n591) );
  NOR2_X1 U651 ( .A1(G164), .A2(G1384), .ZN(n590) );
  XOR2_X1 U652 ( .A(KEYINPUT65), .B(n590), .Z(n694) );
  NAND2_X1 U653 ( .A1(n591), .A2(n694), .ZN(n592) );
  INV_X1 U654 ( .A(n622), .ZN(n645) );
  XNOR2_X1 U655 ( .A(KEYINPUT25), .B(G2078), .ZN(n977) );
  NAND2_X1 U656 ( .A1(n645), .A2(n977), .ZN(n593) );
  XNOR2_X1 U657 ( .A(n593), .B(KEYINPUT95), .ZN(n595) );
  NOR2_X1 U658 ( .A1(n645), .A2(G1961), .ZN(n594) );
  NOR2_X1 U659 ( .A1(n595), .A2(n594), .ZN(n656) );
  OR2_X1 U660 ( .A1(n656), .A2(G301), .ZN(n655) );
  NAND2_X1 U661 ( .A1(G2072), .A2(n645), .ZN(n596) );
  XNOR2_X1 U662 ( .A(KEYINPUT27), .B(n596), .ZN(n599) );
  NAND2_X1 U663 ( .A1(n622), .A2(G1956), .ZN(n597) );
  XOR2_X1 U664 ( .A(KEYINPUT96), .B(n597), .Z(n598) );
  NOR2_X1 U665 ( .A1(n599), .A2(n598), .ZN(n637) );
  NAND2_X1 U666 ( .A1(n803), .A2(G53), .ZN(n601) );
  NAND2_X1 U667 ( .A1(G65), .A2(n804), .ZN(n600) );
  NAND2_X1 U668 ( .A1(n601), .A2(n600), .ZN(n605) );
  NAND2_X1 U669 ( .A1(n807), .A2(G78), .ZN(n603) );
  NAND2_X1 U670 ( .A1(G91), .A2(n808), .ZN(n602) );
  NAND2_X1 U671 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U672 ( .A1(n605), .A2(n604), .ZN(n927) );
  NAND2_X1 U673 ( .A1(n637), .A2(n927), .ZN(n648) );
  INV_X1 U674 ( .A(n648), .ZN(n636) );
  XNOR2_X1 U675 ( .A(KEYINPUT77), .B(KEYINPUT13), .ZN(n611) );
  NAND2_X1 U676 ( .A1(n808), .A2(G81), .ZN(n606) );
  XNOR2_X1 U677 ( .A(n606), .B(KEYINPUT76), .ZN(n607) );
  XNOR2_X1 U678 ( .A(n607), .B(KEYINPUT12), .ZN(n609) );
  NAND2_X1 U679 ( .A1(G68), .A2(n807), .ZN(n608) );
  NAND2_X1 U680 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U681 ( .A(n611), .B(n610), .ZN(n615) );
  NAND2_X1 U682 ( .A1(n804), .A2(G56), .ZN(n612) );
  XNOR2_X1 U683 ( .A(n612), .B(KEYINPUT75), .ZN(n613) );
  XNOR2_X1 U684 ( .A(n613), .B(KEYINPUT14), .ZN(n614) );
  NOR2_X1 U685 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U686 ( .A(n616), .B(KEYINPUT78), .ZN(n618) );
  NAND2_X1 U687 ( .A1(G43), .A2(n803), .ZN(n617) );
  NAND2_X1 U688 ( .A1(n618), .A2(n617), .ZN(n942) );
  NAND2_X1 U689 ( .A1(n645), .A2(G1996), .ZN(n620) );
  XNOR2_X1 U690 ( .A(n620), .B(n619), .ZN(n621) );
  NOR2_X1 U691 ( .A1(n942), .A2(n621), .ZN(n625) );
  NAND2_X1 U692 ( .A1(n669), .A2(G1341), .ZN(n623) );
  XOR2_X1 U693 ( .A(KEYINPUT99), .B(n623), .Z(n624) );
  NAND2_X1 U694 ( .A1(n625), .A2(n624), .ZN(n643) );
  NAND2_X1 U695 ( .A1(G92), .A2(n808), .ZN(n627) );
  NAND2_X1 U696 ( .A1(G66), .A2(n804), .ZN(n626) );
  NAND2_X1 U697 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U698 ( .A(n628), .B(KEYINPUT79), .ZN(n630) );
  NAND2_X1 U699 ( .A1(G54), .A2(n803), .ZN(n629) );
  NAND2_X1 U700 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U701 ( .A1(n807), .A2(G79), .ZN(n631) );
  XOR2_X1 U702 ( .A(KEYINPUT80), .B(n631), .Z(n632) );
  NOR2_X1 U703 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U704 ( .A(KEYINPUT15), .B(n634), .ZN(n934) );
  NAND2_X1 U705 ( .A1(n643), .A2(n934), .ZN(n635) );
  OR2_X1 U706 ( .A1(n636), .A2(n635), .ZN(n642) );
  NOR2_X1 U707 ( .A1(n637), .A2(n927), .ZN(n640) );
  XNOR2_X1 U708 ( .A(KEYINPUT28), .B(KEYINPUT98), .ZN(n638) );
  XNOR2_X1 U709 ( .A(n638), .B(KEYINPUT97), .ZN(n639) );
  XNOR2_X1 U710 ( .A(n640), .B(n639), .ZN(n641) );
  AND2_X1 U711 ( .A1(n642), .A2(n641), .ZN(n653) );
  XOR2_X1 U712 ( .A(n644), .B(KEYINPUT100), .Z(n651) );
  NOR2_X1 U713 ( .A1(G1348), .A2(n645), .ZN(n647) );
  NOR2_X1 U714 ( .A1(G2067), .A2(n669), .ZN(n646) );
  NOR2_X1 U715 ( .A1(n647), .A2(n646), .ZN(n649) );
  AND2_X1 U716 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U717 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U718 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U719 ( .A1(n655), .A2(n519), .ZN(n677) );
  NAND2_X1 U720 ( .A1(n656), .A2(G301), .ZN(n657) );
  XNOR2_X1 U721 ( .A(n657), .B(KEYINPUT101), .ZN(n662) );
  NAND2_X1 U722 ( .A1(n669), .A2(G8), .ZN(n734) );
  NOR2_X1 U723 ( .A1(G1966), .A2(n734), .ZN(n665) );
  NOR2_X1 U724 ( .A1(n669), .A2(G2084), .ZN(n664) );
  NOR2_X1 U725 ( .A1(n665), .A2(n664), .ZN(n658) );
  NAND2_X1 U726 ( .A1(G8), .A2(n658), .ZN(n659) );
  XNOR2_X1 U727 ( .A(KEYINPUT30), .B(n659), .ZN(n660) );
  NOR2_X1 U728 ( .A1(G168), .A2(n660), .ZN(n661) );
  NOR2_X1 U729 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U730 ( .A(KEYINPUT31), .B(n663), .Z(n675) );
  AND2_X1 U731 ( .A1(n677), .A2(n675), .ZN(n668) );
  AND2_X1 U732 ( .A1(G8), .A2(n664), .ZN(n666) );
  OR2_X1 U733 ( .A1(n666), .A2(n665), .ZN(n667) );
  INV_X1 U734 ( .A(G8), .ZN(n674) );
  NOR2_X1 U735 ( .A1(G1971), .A2(n734), .ZN(n671) );
  NOR2_X1 U736 ( .A1(n669), .A2(G2090), .ZN(n670) );
  NOR2_X1 U737 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U738 ( .A1(n672), .A2(G303), .ZN(n673) );
  OR2_X1 U739 ( .A1(n674), .A2(n673), .ZN(n678) );
  AND2_X1 U740 ( .A1(n675), .A2(n678), .ZN(n676) );
  NAND2_X1 U741 ( .A1(n677), .A2(n676), .ZN(n681) );
  INV_X1 U742 ( .A(n678), .ZN(n679) );
  OR2_X1 U743 ( .A1(n679), .A2(G286), .ZN(n680) );
  NAND2_X1 U744 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U745 ( .A(n682), .B(KEYINPUT32), .ZN(n683) );
  NAND2_X1 U746 ( .A1(n684), .A2(n683), .ZN(n729) );
  NOR2_X1 U747 ( .A1(G2090), .A2(G303), .ZN(n685) );
  NAND2_X1 U748 ( .A1(G8), .A2(n685), .ZN(n686) );
  NAND2_X1 U749 ( .A1(n729), .A2(n686), .ZN(n687) );
  NAND2_X1 U750 ( .A1(n687), .A2(n734), .ZN(n692) );
  NOR2_X1 U751 ( .A1(G1981), .A2(G305), .ZN(n688) );
  XOR2_X1 U752 ( .A(n688), .B(KEYINPUT24), .Z(n689) );
  NOR2_X1 U753 ( .A1(n734), .A2(n689), .ZN(n690) );
  XOR2_X1 U754 ( .A(n690), .B(KEYINPUT94), .Z(n691) );
  NAND2_X1 U755 ( .A1(n692), .A2(n691), .ZN(n724) );
  NOR2_X1 U756 ( .A1(n694), .A2(n693), .ZN(n757) );
  XNOR2_X1 U757 ( .A(G2067), .B(KEYINPUT37), .ZN(n754) );
  NAND2_X1 U758 ( .A1(G140), .A2(n890), .ZN(n696) );
  NAND2_X1 U759 ( .A1(G104), .A2(n891), .ZN(n695) );
  NAND2_X1 U760 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U761 ( .A(KEYINPUT34), .B(n697), .ZN(n702) );
  NAND2_X1 U762 ( .A1(G116), .A2(n895), .ZN(n699) );
  NAND2_X1 U763 ( .A1(G128), .A2(n898), .ZN(n698) );
  NAND2_X1 U764 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U765 ( .A(KEYINPUT35), .B(n700), .Z(n701) );
  NOR2_X1 U766 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U767 ( .A(KEYINPUT36), .B(n703), .ZN(n908) );
  NOR2_X1 U768 ( .A1(n754), .A2(n908), .ZN(n1004) );
  NAND2_X1 U769 ( .A1(n757), .A2(n1004), .ZN(n752) );
  NAND2_X1 U770 ( .A1(G131), .A2(n890), .ZN(n705) );
  NAND2_X1 U771 ( .A1(G107), .A2(n895), .ZN(n704) );
  NAND2_X1 U772 ( .A1(n705), .A2(n704), .ZN(n709) );
  NAND2_X1 U773 ( .A1(n898), .A2(G119), .ZN(n707) );
  NAND2_X1 U774 ( .A1(G95), .A2(n891), .ZN(n706) );
  NAND2_X1 U775 ( .A1(n707), .A2(n706), .ZN(n708) );
  OR2_X1 U776 ( .A1(n709), .A2(n708), .ZN(n904) );
  NAND2_X1 U777 ( .A1(G1991), .A2(n904), .ZN(n710) );
  XOR2_X1 U778 ( .A(KEYINPUT90), .B(n710), .Z(n721) );
  NAND2_X1 U779 ( .A1(G117), .A2(n895), .ZN(n712) );
  NAND2_X1 U780 ( .A1(G129), .A2(n898), .ZN(n711) );
  NAND2_X1 U781 ( .A1(n712), .A2(n711), .ZN(n716) );
  NAND2_X1 U782 ( .A1(n891), .A2(G105), .ZN(n713) );
  XNOR2_X1 U783 ( .A(n713), .B(KEYINPUT38), .ZN(n714) );
  XNOR2_X1 U784 ( .A(n714), .B(KEYINPUT91), .ZN(n715) );
  NOR2_X1 U785 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U786 ( .A(KEYINPUT92), .B(n717), .ZN(n719) );
  NAND2_X1 U787 ( .A1(G141), .A2(n890), .ZN(n718) );
  NAND2_X1 U788 ( .A1(n719), .A2(n718), .ZN(n910) );
  AND2_X1 U789 ( .A1(n910), .A2(G1996), .ZN(n720) );
  NOR2_X1 U790 ( .A1(n721), .A2(n720), .ZN(n997) );
  XOR2_X1 U791 ( .A(G1986), .B(G290), .Z(n940) );
  NAND2_X1 U792 ( .A1(n997), .A2(n940), .ZN(n722) );
  NAND2_X1 U793 ( .A1(n722), .A2(n757), .ZN(n725) );
  AND2_X1 U794 ( .A1(n752), .A2(n725), .ZN(n723) );
  AND2_X1 U795 ( .A1(n724), .A2(n723), .ZN(n745) );
  INV_X1 U796 ( .A(n725), .ZN(n743) );
  NOR2_X1 U797 ( .A1(G1976), .A2(G288), .ZN(n732) );
  NOR2_X1 U798 ( .A1(G1971), .A2(G303), .ZN(n726) );
  NOR2_X1 U799 ( .A1(n732), .A2(n726), .ZN(n928) );
  INV_X1 U800 ( .A(KEYINPUT33), .ZN(n727) );
  AND2_X1 U801 ( .A1(n928), .A2(n727), .ZN(n728) );
  NAND2_X1 U802 ( .A1(n729), .A2(n728), .ZN(n741) );
  INV_X1 U803 ( .A(n734), .ZN(n730) );
  NAND2_X1 U804 ( .A1(G1976), .A2(G288), .ZN(n931) );
  AND2_X1 U805 ( .A1(n730), .A2(n931), .ZN(n731) );
  NOR2_X1 U806 ( .A1(KEYINPUT33), .A2(n731), .ZN(n739) );
  NAND2_X1 U807 ( .A1(n732), .A2(KEYINPUT33), .ZN(n733) );
  XOR2_X1 U808 ( .A(G1981), .B(G305), .Z(n924) );
  INV_X1 U809 ( .A(n924), .ZN(n735) );
  OR2_X1 U810 ( .A1(n518), .A2(n735), .ZN(n737) );
  INV_X1 U811 ( .A(n752), .ZN(n736) );
  OR2_X1 U812 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U813 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U814 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U815 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U816 ( .A1(n745), .A2(n744), .ZN(n760) );
  INV_X1 U817 ( .A(n997), .ZN(n748) );
  NOR2_X1 U818 ( .A1(G1986), .A2(G290), .ZN(n746) );
  NOR2_X1 U819 ( .A1(G1991), .A2(n904), .ZN(n1003) );
  NOR2_X1 U820 ( .A1(n746), .A2(n1003), .ZN(n747) );
  NOR2_X1 U821 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U822 ( .A1(G1996), .A2(n910), .ZN(n999) );
  NOR2_X1 U823 ( .A1(n749), .A2(n999), .ZN(n750) );
  XNOR2_X1 U824 ( .A(n750), .B(KEYINPUT102), .ZN(n751) );
  XNOR2_X1 U825 ( .A(n751), .B(KEYINPUT39), .ZN(n753) );
  NAND2_X1 U826 ( .A1(n753), .A2(n752), .ZN(n755) );
  NAND2_X1 U827 ( .A1(n754), .A2(n908), .ZN(n996) );
  NAND2_X1 U828 ( .A1(n755), .A2(n996), .ZN(n756) );
  XOR2_X1 U829 ( .A(KEYINPUT103), .B(n756), .Z(n758) );
  NAND2_X1 U830 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U831 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U832 ( .A(n761), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U833 ( .A(KEYINPUT104), .B(KEYINPUT106), .Z(n763) );
  XNOR2_X1 U834 ( .A(G2446), .B(G2451), .ZN(n762) );
  XNOR2_X1 U835 ( .A(n763), .B(n762), .ZN(n767) );
  XOR2_X1 U836 ( .A(G2435), .B(G2438), .Z(n765) );
  XNOR2_X1 U837 ( .A(G2454), .B(G2430), .ZN(n764) );
  XNOR2_X1 U838 ( .A(n765), .B(n764), .ZN(n766) );
  XOR2_X1 U839 ( .A(n767), .B(n766), .Z(n769) );
  XNOR2_X1 U840 ( .A(G2443), .B(G2427), .ZN(n768) );
  XNOR2_X1 U841 ( .A(n769), .B(n768), .ZN(n772) );
  XOR2_X1 U842 ( .A(G1341), .B(G1348), .Z(n770) );
  XNOR2_X1 U843 ( .A(KEYINPUT105), .B(n770), .ZN(n771) );
  XOR2_X1 U844 ( .A(n772), .B(n771), .Z(n773) );
  AND2_X1 U845 ( .A1(G14), .A2(n773), .ZN(G401) );
  AND2_X1 U846 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U847 ( .A(G120), .ZN(G236) );
  INV_X1 U848 ( .A(G69), .ZN(G235) );
  INV_X1 U849 ( .A(G108), .ZN(G238) );
  NAND2_X1 U850 ( .A1(G7), .A2(G661), .ZN(n774) );
  XNOR2_X1 U851 ( .A(n774), .B(KEYINPUT10), .ZN(n775) );
  XNOR2_X1 U852 ( .A(KEYINPUT74), .B(n775), .ZN(G223) );
  INV_X1 U853 ( .A(G223), .ZN(n839) );
  NAND2_X1 U854 ( .A1(n839), .A2(G567), .ZN(n776) );
  XOR2_X1 U855 ( .A(KEYINPUT11), .B(n776), .Z(G234) );
  INV_X1 U856 ( .A(G860), .ZN(n802) );
  OR2_X1 U857 ( .A1(n942), .A2(n802), .ZN(G153) );
  NAND2_X1 U858 ( .A1(G868), .A2(G301), .ZN(n778) );
  INV_X1 U859 ( .A(G868), .ZN(n779) );
  NAND2_X1 U860 ( .A1(n934), .A2(n779), .ZN(n777) );
  NAND2_X1 U861 ( .A1(n778), .A2(n777), .ZN(G284) );
  INV_X1 U862 ( .A(n927), .ZN(G299) );
  NAND2_X1 U863 ( .A1(G868), .A2(G286), .ZN(n781) );
  NAND2_X1 U864 ( .A1(G299), .A2(n779), .ZN(n780) );
  NAND2_X1 U865 ( .A1(n781), .A2(n780), .ZN(G297) );
  NAND2_X1 U866 ( .A1(G559), .A2(n802), .ZN(n782) );
  XOR2_X1 U867 ( .A(KEYINPUT83), .B(n782), .Z(n783) );
  INV_X1 U868 ( .A(n934), .ZN(n800) );
  NAND2_X1 U869 ( .A1(n783), .A2(n800), .ZN(n784) );
  XNOR2_X1 U870 ( .A(n784), .B(KEYINPUT16), .ZN(n785) );
  XNOR2_X1 U871 ( .A(KEYINPUT84), .B(n785), .ZN(G148) );
  NOR2_X1 U872 ( .A1(G868), .A2(n942), .ZN(n788) );
  NAND2_X1 U873 ( .A1(G868), .A2(n800), .ZN(n786) );
  NOR2_X1 U874 ( .A1(G559), .A2(n786), .ZN(n787) );
  NOR2_X1 U875 ( .A1(n788), .A2(n787), .ZN(G282) );
  NAND2_X1 U876 ( .A1(G135), .A2(n890), .ZN(n790) );
  NAND2_X1 U877 ( .A1(G111), .A2(n895), .ZN(n789) );
  NAND2_X1 U878 ( .A1(n790), .A2(n789), .ZN(n797) );
  NAND2_X1 U879 ( .A1(n891), .A2(G99), .ZN(n791) );
  XNOR2_X1 U880 ( .A(n791), .B(KEYINPUT86), .ZN(n795) );
  XOR2_X1 U881 ( .A(KEYINPUT18), .B(KEYINPUT85), .Z(n793) );
  NAND2_X1 U882 ( .A1(G123), .A2(n898), .ZN(n792) );
  XNOR2_X1 U883 ( .A(n793), .B(n792), .ZN(n794) );
  NAND2_X1 U884 ( .A1(n795), .A2(n794), .ZN(n796) );
  NOR2_X1 U885 ( .A1(n797), .A2(n796), .ZN(n1002) );
  XNOR2_X1 U886 ( .A(n1002), .B(G2096), .ZN(n799) );
  INV_X1 U887 ( .A(G2100), .ZN(n798) );
  NAND2_X1 U888 ( .A1(n799), .A2(n798), .ZN(G156) );
  NAND2_X1 U889 ( .A1(G559), .A2(n800), .ZN(n801) );
  XOR2_X1 U890 ( .A(n942), .B(n801), .Z(n819) );
  NAND2_X1 U891 ( .A1(n802), .A2(n819), .ZN(n813) );
  NAND2_X1 U892 ( .A1(n803), .A2(G55), .ZN(n806) );
  NAND2_X1 U893 ( .A1(G67), .A2(n804), .ZN(n805) );
  NAND2_X1 U894 ( .A1(n806), .A2(n805), .ZN(n812) );
  NAND2_X1 U895 ( .A1(n807), .A2(G80), .ZN(n810) );
  NAND2_X1 U896 ( .A1(G93), .A2(n808), .ZN(n809) );
  NAND2_X1 U897 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U898 ( .A1(n812), .A2(n811), .ZN(n821) );
  XOR2_X1 U899 ( .A(n813), .B(n821), .Z(G145) );
  XNOR2_X1 U900 ( .A(n927), .B(KEYINPUT19), .ZN(n815) );
  XNOR2_X1 U901 ( .A(G288), .B(G166), .ZN(n814) );
  XNOR2_X1 U902 ( .A(n815), .B(n814), .ZN(n816) );
  XOR2_X1 U903 ( .A(n821), .B(n816), .Z(n817) );
  XNOR2_X1 U904 ( .A(G305), .B(n817), .ZN(n818) );
  XNOR2_X1 U905 ( .A(n818), .B(G290), .ZN(n914) );
  XNOR2_X1 U906 ( .A(n819), .B(n914), .ZN(n820) );
  NAND2_X1 U907 ( .A1(n820), .A2(G868), .ZN(n823) );
  OR2_X1 U908 ( .A1(G868), .A2(n821), .ZN(n822) );
  NAND2_X1 U909 ( .A1(n823), .A2(n822), .ZN(G295) );
  NAND2_X1 U910 ( .A1(G2078), .A2(G2084), .ZN(n824) );
  XOR2_X1 U911 ( .A(KEYINPUT20), .B(n824), .Z(n825) );
  NAND2_X1 U912 ( .A1(G2090), .A2(n825), .ZN(n826) );
  XNOR2_X1 U913 ( .A(KEYINPUT21), .B(n826), .ZN(n827) );
  NAND2_X1 U914 ( .A1(n827), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U915 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U916 ( .A1(G235), .A2(G236), .ZN(n828) );
  XNOR2_X1 U917 ( .A(n828), .B(KEYINPUT89), .ZN(n829) );
  NOR2_X1 U918 ( .A1(G238), .A2(n829), .ZN(n830) );
  NAND2_X1 U919 ( .A1(G57), .A2(n830), .ZN(n845) );
  NAND2_X1 U920 ( .A1(G567), .A2(n845), .ZN(n837) );
  XOR2_X1 U921 ( .A(KEYINPUT22), .B(KEYINPUT87), .Z(n832) );
  NAND2_X1 U922 ( .A1(G132), .A2(G82), .ZN(n831) );
  XNOR2_X1 U923 ( .A(n832), .B(n831), .ZN(n833) );
  NOR2_X1 U924 ( .A1(n833), .A2(G218), .ZN(n834) );
  XNOR2_X1 U925 ( .A(KEYINPUT88), .B(n834), .ZN(n835) );
  NAND2_X1 U926 ( .A1(n835), .A2(G96), .ZN(n844) );
  NAND2_X1 U927 ( .A1(G2106), .A2(n844), .ZN(n836) );
  NAND2_X1 U928 ( .A1(n837), .A2(n836), .ZN(n847) );
  NAND2_X1 U929 ( .A1(G661), .A2(G483), .ZN(n838) );
  NOR2_X1 U930 ( .A1(n847), .A2(n838), .ZN(n841) );
  NAND2_X1 U931 ( .A1(n841), .A2(G36), .ZN(G176) );
  NAND2_X1 U932 ( .A1(G2106), .A2(n839), .ZN(G217) );
  AND2_X1 U933 ( .A1(G15), .A2(G2), .ZN(n840) );
  NAND2_X1 U934 ( .A1(G661), .A2(n840), .ZN(G259) );
  NAND2_X1 U935 ( .A1(G3), .A2(G1), .ZN(n842) );
  NAND2_X1 U936 ( .A1(n842), .A2(n841), .ZN(n843) );
  XOR2_X1 U937 ( .A(KEYINPUT107), .B(n843), .Z(G188) );
  INV_X1 U939 ( .A(G132), .ZN(G219) );
  INV_X1 U940 ( .A(G96), .ZN(G221) );
  INV_X1 U941 ( .A(G82), .ZN(G220) );
  NOR2_X1 U942 ( .A1(n845), .A2(n844), .ZN(n846) );
  XNOR2_X1 U943 ( .A(n846), .B(KEYINPUT108), .ZN(G325) );
  INV_X1 U944 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U945 ( .A(KEYINPUT109), .B(n847), .ZN(G319) );
  XOR2_X1 U946 ( .A(G2100), .B(G2096), .Z(n849) );
  XNOR2_X1 U947 ( .A(KEYINPUT42), .B(G2678), .ZN(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U949 ( .A(KEYINPUT43), .B(G2090), .Z(n851) );
  XNOR2_X1 U950 ( .A(G2067), .B(G2072), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U952 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U953 ( .A(G2078), .B(G2084), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(G227) );
  XNOR2_X1 U955 ( .A(G1991), .B(KEYINPUT110), .ZN(n865) );
  XOR2_X1 U956 ( .A(G1961), .B(G1966), .Z(n857) );
  XNOR2_X1 U957 ( .A(G1996), .B(G1981), .ZN(n856) );
  XNOR2_X1 U958 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U959 ( .A(G1956), .B(G1971), .Z(n859) );
  XNOR2_X1 U960 ( .A(G1986), .B(G1976), .ZN(n858) );
  XNOR2_X1 U961 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U962 ( .A(n861), .B(n860), .Z(n863) );
  XNOR2_X1 U963 ( .A(G2474), .B(KEYINPUT41), .ZN(n862) );
  XNOR2_X1 U964 ( .A(n863), .B(n862), .ZN(n864) );
  XNOR2_X1 U965 ( .A(n865), .B(n864), .ZN(G229) );
  NAND2_X1 U966 ( .A1(G124), .A2(n898), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n866), .B(KEYINPUT44), .ZN(n871) );
  NAND2_X1 U968 ( .A1(n895), .A2(G112), .ZN(n868) );
  NAND2_X1 U969 ( .A1(G100), .A2(n891), .ZN(n867) );
  NAND2_X1 U970 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U971 ( .A(KEYINPUT112), .B(n869), .Z(n870) );
  NAND2_X1 U972 ( .A1(n871), .A2(n870), .ZN(n874) );
  NAND2_X1 U973 ( .A1(G136), .A2(n890), .ZN(n872) );
  XNOR2_X1 U974 ( .A(KEYINPUT111), .B(n872), .ZN(n873) );
  NOR2_X1 U975 ( .A1(n874), .A2(n873), .ZN(G162) );
  NAND2_X1 U976 ( .A1(n898), .A2(G127), .ZN(n875) );
  XNOR2_X1 U977 ( .A(n875), .B(KEYINPUT116), .ZN(n877) );
  NAND2_X1 U978 ( .A1(G115), .A2(n895), .ZN(n876) );
  NAND2_X1 U979 ( .A1(n877), .A2(n876), .ZN(n878) );
  XNOR2_X1 U980 ( .A(n878), .B(KEYINPUT47), .ZN(n883) );
  NAND2_X1 U981 ( .A1(G139), .A2(n890), .ZN(n880) );
  NAND2_X1 U982 ( .A1(G103), .A2(n891), .ZN(n879) );
  NAND2_X1 U983 ( .A1(n880), .A2(n879), .ZN(n881) );
  XNOR2_X1 U984 ( .A(KEYINPUT115), .B(n881), .ZN(n882) );
  NAND2_X1 U985 ( .A1(n883), .A2(n882), .ZN(n884) );
  XNOR2_X1 U986 ( .A(n884), .B(KEYINPUT117), .ZN(n1007) );
  XNOR2_X1 U987 ( .A(G164), .B(n1007), .ZN(n885) );
  XNOR2_X1 U988 ( .A(n885), .B(G162), .ZN(n889) );
  XOR2_X1 U989 ( .A(KEYINPUT114), .B(KEYINPUT46), .Z(n887) );
  XNOR2_X1 U990 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n886) );
  XNOR2_X1 U991 ( .A(n887), .B(n886), .ZN(n888) );
  XOR2_X1 U992 ( .A(n889), .B(n888), .Z(n907) );
  NAND2_X1 U993 ( .A1(G142), .A2(n890), .ZN(n893) );
  NAND2_X1 U994 ( .A1(G106), .A2(n891), .ZN(n892) );
  NAND2_X1 U995 ( .A1(n893), .A2(n892), .ZN(n894) );
  XNOR2_X1 U996 ( .A(n894), .B(KEYINPUT45), .ZN(n897) );
  NAND2_X1 U997 ( .A1(G118), .A2(n895), .ZN(n896) );
  NAND2_X1 U998 ( .A1(n897), .A2(n896), .ZN(n901) );
  NAND2_X1 U999 ( .A1(G130), .A2(n898), .ZN(n899) );
  XNOR2_X1 U1000 ( .A(KEYINPUT113), .B(n899), .ZN(n900) );
  NOR2_X1 U1001 ( .A1(n901), .A2(n900), .ZN(n902) );
  XOR2_X1 U1002 ( .A(n1002), .B(n902), .Z(n903) );
  XNOR2_X1 U1003 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(n905), .B(KEYINPUT48), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(n907), .B(n906), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(n909), .B(n908), .ZN(n911) );
  XNOR2_X1 U1007 ( .A(n911), .B(n910), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(n912), .B(G160), .ZN(n913) );
  NOR2_X1 U1009 ( .A1(G37), .A2(n913), .ZN(G395) );
  XNOR2_X1 U1010 ( .A(n914), .B(n942), .ZN(n915) );
  XNOR2_X1 U1011 ( .A(n915), .B(G286), .ZN(n917) );
  XOR2_X1 U1012 ( .A(n934), .B(G171), .Z(n916) );
  XNOR2_X1 U1013 ( .A(n917), .B(n916), .ZN(n918) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n918), .ZN(G397) );
  NOR2_X1 U1015 ( .A1(G227), .A2(G229), .ZN(n919) );
  XNOR2_X1 U1016 ( .A(KEYINPUT49), .B(n919), .ZN(n920) );
  NOR2_X1 U1017 ( .A1(G401), .A2(n920), .ZN(n922) );
  NOR2_X1 U1018 ( .A1(G395), .A2(G397), .ZN(n921) );
  AND2_X1 U1019 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1020 ( .A1(G319), .A2(n923), .ZN(G225) );
  INV_X1 U1021 ( .A(G225), .ZN(G308) );
  INV_X1 U1022 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1023 ( .A(G1966), .B(G168), .ZN(n925) );
  NAND2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1025 ( .A(KEYINPUT57), .B(n926), .ZN(n946) );
  XNOR2_X1 U1026 ( .A(n927), .B(G1956), .ZN(n929) );
  NAND2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n938) );
  NAND2_X1 U1028 ( .A1(G1971), .A2(G303), .ZN(n930) );
  NAND2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n933) );
  XNOR2_X1 U1030 ( .A(G1961), .B(G301), .ZN(n932) );
  NOR2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n936) );
  XOR2_X1 U1032 ( .A(G1348), .B(n934), .Z(n935) );
  NAND2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1036 ( .A(KEYINPUT125), .B(n941), .Z(n944) );
  XNOR2_X1 U1037 ( .A(G1341), .B(n942), .ZN(n943) );
  NOR2_X1 U1038 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1040 ( .A(KEYINPUT126), .B(n947), .ZN(n950) );
  XNOR2_X1 U1041 ( .A(G16), .B(KEYINPUT56), .ZN(n948) );
  XNOR2_X1 U1042 ( .A(n948), .B(KEYINPUT124), .ZN(n949) );
  NAND2_X1 U1043 ( .A1(n950), .A2(n949), .ZN(n1027) );
  XOR2_X1 U1044 ( .A(G1986), .B(G24), .Z(n954) );
  XNOR2_X1 U1045 ( .A(G1976), .B(G23), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(G1971), .B(G22), .ZN(n951) );
  NOR2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(KEYINPUT58), .B(KEYINPUT127), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(n956), .B(n955), .ZN(n960) );
  XNOR2_X1 U1051 ( .A(G1966), .B(G21), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(G1961), .B(G5), .ZN(n957) );
  NOR2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n970) );
  XOR2_X1 U1055 ( .A(G1348), .B(KEYINPUT59), .Z(n961) );
  XNOR2_X1 U1056 ( .A(G4), .B(n961), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(G20), .B(G1956), .ZN(n962) );
  NOR2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n967) );
  XNOR2_X1 U1059 ( .A(G1981), .B(G6), .ZN(n965) );
  XNOR2_X1 U1060 ( .A(G1341), .B(G19), .ZN(n964) );
  NOR2_X1 U1061 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(KEYINPUT60), .B(n968), .ZN(n969) );
  NOR2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(KEYINPUT61), .B(n971), .ZN(n973) );
  INV_X1 U1066 ( .A(G16), .ZN(n972) );
  NAND2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1068 ( .A1(n974), .A2(G11), .ZN(n1025) );
  XNOR2_X1 U1069 ( .A(KEYINPUT121), .B(G2072), .ZN(n975) );
  XNOR2_X1 U1070 ( .A(n975), .B(G33), .ZN(n985) );
  XOR2_X1 U1071 ( .A(G2067), .B(G26), .Z(n976) );
  NAND2_X1 U1072 ( .A1(n976), .A2(G28), .ZN(n983) );
  XNOR2_X1 U1073 ( .A(G27), .B(n977), .ZN(n981) );
  XNOR2_X1 U1074 ( .A(G1996), .B(G32), .ZN(n979) );
  XNOR2_X1 U1075 ( .A(G1991), .B(G25), .ZN(n978) );
  NOR2_X1 U1076 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1079 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1080 ( .A(n986), .B(KEYINPUT53), .ZN(n987) );
  XNOR2_X1 U1081 ( .A(n987), .B(KEYINPUT122), .ZN(n990) );
  XOR2_X1 U1082 ( .A(G2084), .B(KEYINPUT54), .Z(n988) );
  XNOR2_X1 U1083 ( .A(G34), .B(n988), .ZN(n989) );
  NAND2_X1 U1084 ( .A1(n990), .A2(n989), .ZN(n992) );
  XNOR2_X1 U1085 ( .A(G35), .B(G2090), .ZN(n991) );
  NOR2_X1 U1086 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1087 ( .A(KEYINPUT55), .B(n993), .Z(n994) );
  NOR2_X1 U1088 ( .A1(G29), .A2(n994), .ZN(n995) );
  XNOR2_X1 U1089 ( .A(n995), .B(KEYINPUT123), .ZN(n1023) );
  NAND2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n1017) );
  XOR2_X1 U1091 ( .A(G2090), .B(G162), .Z(n998) );
  NOR2_X1 U1092 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1093 ( .A(KEYINPUT51), .B(n1000), .Z(n1015) );
  XOR2_X1 U1094 ( .A(G2084), .B(G160), .Z(n1001) );
  NOR2_X1 U1095 ( .A1(n1002), .A2(n1001), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1013) );
  XOR2_X1 U1098 ( .A(G2072), .B(n1007), .Z(n1009) );
  XOR2_X1 U1099 ( .A(G164), .B(G2078), .Z(n1008) );
  NOR2_X1 U1100 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1101 ( .A(KEYINPUT120), .B(n1010), .Z(n1011) );
  XNOR2_X1 U1102 ( .A(KEYINPUT50), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1106 ( .A(n1018), .B(KEYINPUT52), .ZN(n1020) );
  INV_X1 U1107 ( .A(KEYINPUT55), .ZN(n1019) );
  NAND2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1109 ( .A1(G29), .A2(n1021), .ZN(n1022) );
  NAND2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XOR2_X1 U1113 ( .A(KEYINPUT62), .B(n1028), .Z(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

