//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1 1 1 0 1 1 0 1 0 0 1 0 0 1 1 1 0 1 0 0 1 0 0 1 1 1 1 0 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n753, new_n754, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012;
  INV_X1    g000(.A(G143), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G146), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT81), .ZN(new_n192));
  OAI211_X1 g006(.A(new_n192), .B(KEYINPUT1), .C1(new_n187), .C2(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G128), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n192), .B1(new_n190), .B2(KEYINPUT1), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n191), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT82), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  OR3_X1    g013(.A1(new_n191), .A2(KEYINPUT1), .A3(new_n199), .ZN(new_n200));
  OAI211_X1 g014(.A(KEYINPUT82), .B(new_n191), .C1(new_n194), .C2(new_n195), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n198), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G104), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT3), .B1(new_n203), .B2(G107), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT3), .ZN(new_n205));
  INV_X1    g019(.A(G107), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(G104), .ZN(new_n207));
  INV_X1    g021(.A(G101), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n203), .A2(G107), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n204), .A2(new_n207), .A3(new_n208), .A4(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n206), .A2(G104), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n203), .A2(G107), .ZN(new_n212));
  OAI21_X1  g026(.A(G101), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AND2_X1   g027(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n202), .A2(new_n214), .ZN(new_n215));
  XOR2_X1   g029(.A(KEYINPUT83), .B(KEYINPUT10), .Z(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n199), .B1(new_n190), .B2(KEYINPUT1), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n219), .B1(new_n189), .B2(G143), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n187), .A2(KEYINPUT65), .A3(G146), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT64), .B1(new_n187), .B2(G146), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT64), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n224), .A2(new_n189), .A3(G143), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n218), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  NOR3_X1   g041(.A1(new_n191), .A2(KEYINPUT1), .A3(new_n199), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n214), .B(KEYINPUT10), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT84), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n190), .A2(KEYINPUT1), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G128), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n223), .A2(new_n225), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n220), .A2(new_n221), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(new_n200), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n237), .A2(KEYINPUT84), .A3(KEYINPUT10), .A4(new_n214), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n231), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT11), .ZN(new_n240));
  INV_X1    g054(.A(G134), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n240), .B1(new_n241), .B2(G137), .ZN(new_n242));
  INV_X1    g056(.A(G137), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(KEYINPUT11), .A3(G134), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n241), .A2(G137), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n242), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(KEYINPUT66), .A2(G131), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n242), .A2(new_n244), .A3(new_n247), .A4(new_n245), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  AND4_X1   g066(.A1(KEYINPUT0), .A2(new_n188), .A3(new_n190), .A4(G128), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n224), .B1(G143), .B2(new_n189), .ZN(new_n254));
  NOR3_X1   g068(.A1(new_n187), .A2(KEYINPUT64), .A3(G146), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n220), .B(new_n221), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  XOR2_X1   g070(.A(KEYINPUT0), .B(G128), .Z(new_n257));
  AOI21_X1  g071(.A(new_n253), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n204), .A2(new_n207), .A3(new_n209), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n259), .A2(G101), .ZN(new_n260));
  XOR2_X1   g074(.A(KEYINPUT80), .B(KEYINPUT4), .Z(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n259), .A2(G101), .ZN(new_n263));
  OAI211_X1 g077(.A(KEYINPUT4), .B(new_n210), .C1(new_n263), .C2(KEYINPUT79), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT79), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n265), .B1(new_n259), .B2(G101), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n258), .B(new_n262), .C1(new_n264), .C2(new_n266), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n217), .A2(new_n239), .A3(new_n252), .A4(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT85), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n210), .A2(KEYINPUT4), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n271), .B1(new_n260), .B2(new_n265), .ZN(new_n272));
  INV_X1    g086(.A(new_n266), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n272), .A2(new_n273), .B1(new_n260), .B2(new_n261), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n258), .A2(new_n274), .B1(new_n231), .B2(new_n238), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n275), .A2(KEYINPUT85), .A3(new_n252), .A4(new_n217), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n270), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(G110), .B(G140), .ZN(new_n278));
  INV_X1    g092(.A(G953), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n279), .A2(G227), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n278), .B(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n215), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n237), .A2(new_n214), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n251), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT12), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI211_X1 g101(.A(KEYINPUT12), .B(new_n251), .C1(new_n283), .C2(new_n284), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n277), .A2(new_n282), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT86), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n277), .A2(new_n289), .A3(KEYINPUT86), .A4(new_n282), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n275), .A2(new_n217), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n251), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n277), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(new_n281), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n292), .A2(new_n293), .A3(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G469), .ZN(new_n299));
  INV_X1    g113(.A(G902), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n299), .A2(new_n300), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n282), .B1(new_n277), .B2(new_n289), .ZN(new_n303));
  AND2_X1   g117(.A1(new_n277), .A2(new_n295), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n303), .B1(new_n282), .B2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n302), .B1(new_n305), .B2(G469), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT9), .B(G234), .ZN(new_n308));
  OAI21_X1  g122(.A(G221), .B1(new_n308), .B2(G902), .ZN(new_n309));
  OAI21_X1  g123(.A(G210), .B1(G237), .B2(G902), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(G110), .B(G122), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  OR2_X1    g127(.A1(KEYINPUT68), .A2(G116), .ZN(new_n314));
  NAND2_X1  g128(.A1(KEYINPUT68), .A2(G116), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n314), .A2(G119), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT67), .ZN(new_n317));
  INV_X1    g131(.A(G119), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(KEYINPUT67), .A2(G119), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(G116), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT2), .B(G113), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n323), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(new_n316), .A3(new_n321), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n327), .B(new_n262), .C1(new_n264), .C2(new_n266), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n214), .A2(new_n326), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT5), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n319), .A2(new_n331), .A3(G116), .A4(new_n320), .ZN(new_n332));
  AND2_X1   g146(.A1(new_n332), .A2(G113), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n316), .A2(new_n321), .A3(KEYINPUT5), .ZN(new_n334));
  AOI21_X1  g148(.A(KEYINPUT87), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n333), .A2(KEYINPUT87), .A3(new_n334), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n330), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n313), .B1(new_n329), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n330), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n333), .A2(KEYINPUT87), .A3(new_n334), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n340), .B1(new_n341), .B2(new_n335), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(new_n328), .A3(new_n312), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n339), .A2(KEYINPUT6), .A3(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT76), .B(G125), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n237), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n258), .A2(new_n345), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n279), .A2(G224), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n349), .B(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT6), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n352), .B(new_n313), .C1(new_n329), .C2(new_n338), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n344), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT89), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n350), .A2(KEYINPUT7), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n356), .B1(new_n347), .B2(new_n348), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n347), .A2(new_n348), .A3(new_n356), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n343), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  XOR2_X1   g174(.A(new_n312), .B(KEYINPUT8), .Z(new_n361));
  OAI21_X1  g175(.A(new_n326), .B1(new_n341), .B2(new_n335), .ZN(new_n362));
  INV_X1    g176(.A(new_n214), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n332), .A2(G113), .ZN(new_n365));
  OR2_X1    g179(.A1(new_n365), .A2(KEYINPUT88), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(KEYINPUT88), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(new_n334), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n340), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n361), .B1(new_n364), .B2(new_n369), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n355), .B(new_n300), .C1(new_n360), .C2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n354), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n359), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n373), .A2(new_n357), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n362), .A2(new_n363), .B1(new_n340), .B2(new_n368), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n374), .B(new_n343), .C1(new_n375), .C2(new_n361), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n355), .B1(new_n376), .B2(new_n300), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n311), .B1(new_n372), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n300), .B1(new_n360), .B2(new_n370), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT89), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n380), .A2(new_n310), .A3(new_n354), .A4(new_n371), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT93), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT92), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n187), .A2(G128), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n199), .A2(G143), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n385), .A2(new_n386), .A3(new_n384), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n241), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n389), .ZN(new_n391));
  NOR3_X1   g205(.A1(new_n391), .A2(G134), .A3(new_n387), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n383), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n388), .A2(new_n389), .A3(new_n241), .ZN(new_n394));
  OAI21_X1  g208(.A(G134), .B1(new_n391), .B2(new_n387), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n395), .A3(KEYINPUT93), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n314), .A2(G122), .A3(new_n315), .ZN(new_n397));
  INV_X1    g211(.A(G122), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G116), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n206), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n397), .A2(G107), .A3(new_n399), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n399), .A2(KEYINPUT14), .A3(G107), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n397), .A2(KEYINPUT14), .A3(G107), .A4(new_n399), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n393), .A2(new_n396), .A3(new_n404), .A4(new_n405), .ZN(new_n406));
  XOR2_X1   g220(.A(KEYINPUT91), .B(KEYINPUT13), .Z(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(G128), .A3(new_n187), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n385), .A2(new_n386), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n408), .B(G134), .C1(new_n409), .C2(new_n407), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n410), .A2(new_n394), .A3(new_n401), .A4(new_n402), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n406), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G217), .ZN(new_n413));
  NOR3_X1   g227(.A1(new_n308), .A2(new_n413), .A3(G953), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n406), .A2(new_n411), .A3(new_n414), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n416), .A2(KEYINPUT94), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT94), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n412), .A2(new_n419), .A3(new_n415), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n418), .A2(new_n300), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(G478), .ZN(new_n422));
  NOR2_X1   g236(.A1(KEYINPUT95), .A2(KEYINPUT15), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(KEYINPUT95), .A2(KEYINPUT15), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n422), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n421), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n426), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n418), .A2(new_n300), .A3(new_n420), .A4(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(G234), .A2(G237), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n430), .A2(G952), .A3(new_n279), .ZN(new_n431));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(G898), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n430), .A2(G902), .A3(G953), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n431), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(KEYINPUT96), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT16), .ZN(new_n438));
  INV_X1    g252(.A(G140), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n345), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(G125), .A2(G140), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n441), .B1(new_n345), .B2(G140), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n440), .B1(new_n442), .B2(new_n438), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n189), .ZN(new_n444));
  OAI211_X1 g258(.A(G146), .B(new_n440), .C1(new_n442), .C2(new_n438), .ZN(new_n445));
  NOR2_X1   g259(.A1(G237), .A2(G953), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(G214), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n187), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n446), .A2(G143), .A3(G214), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(KEYINPUT17), .A3(G131), .ZN(new_n451));
  INV_X1    g265(.A(new_n449), .ZN(new_n452));
  AOI21_X1  g266(.A(G143), .B1(new_n446), .B2(G214), .ZN(new_n453));
  OAI21_X1  g267(.A(G131), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT17), .ZN(new_n455));
  INV_X1    g269(.A(G131), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n448), .A2(new_n456), .A3(new_n449), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n454), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n444), .A2(new_n445), .A3(new_n451), .A4(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n441), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT77), .ZN(new_n461));
  NAND2_X1  g275(.A1(G125), .A2(G140), .ZN(new_n462));
  AND3_X1   g276(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n461), .B1(new_n460), .B2(new_n462), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n189), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n442), .A2(G146), .ZN(new_n466));
  NAND2_X1  g280(.A1(KEYINPUT18), .A2(G131), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  AOI22_X1  g282(.A1(new_n465), .A2(new_n466), .B1(new_n450), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(KEYINPUT90), .B1(new_n450), .B2(new_n468), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT90), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n448), .A2(new_n471), .A3(new_n449), .A4(new_n467), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(G113), .B(G122), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n475), .B(new_n203), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n459), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n476), .B1(new_n459), .B2(new_n474), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n300), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n437), .B1(new_n479), .B2(G475), .ZN(new_n480));
  NOR2_X1   g294(.A1(G475), .A2(G902), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n442), .A2(KEYINPUT19), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n463), .A2(new_n464), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n482), .B(new_n189), .C1(new_n483), .C2(KEYINPUT19), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n454), .A2(new_n457), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n445), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n476), .B1(new_n486), .B2(new_n474), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n481), .B1(new_n477), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT20), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n459), .A2(new_n474), .A3(new_n476), .ZN(new_n490));
  AND2_X1   g304(.A1(new_n445), .A2(new_n485), .ZN(new_n491));
  AOI22_X1  g305(.A1(new_n491), .A2(new_n484), .B1(new_n469), .B2(new_n473), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n490), .B1(new_n492), .B2(new_n476), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT20), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(new_n494), .A3(new_n481), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n489), .A2(new_n495), .ZN(new_n496));
  AND4_X1   g310(.A1(new_n427), .A2(new_n429), .A3(new_n480), .A4(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(G214), .B1(G237), .B2(G902), .ZN(new_n498));
  AND3_X1   g312(.A1(new_n382), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n307), .A2(new_n309), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(KEYINPUT97), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n413), .B1(G234), .B2(new_n300), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n279), .A2(G221), .A3(G234), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(KEYINPUT78), .ZN(new_n504));
  XNOR2_X1  g318(.A(KEYINPUT22), .B(G137), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n504), .B(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n444), .A2(new_n445), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n319), .A2(G128), .A3(new_n320), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n318), .A2(G128), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT24), .B(G110), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n508), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT75), .ZN(new_n517));
  AOI21_X1  g331(.A(G128), .B1(new_n319), .B2(new_n320), .ZN(new_n518));
  AOI22_X1  g332(.A1(KEYINPUT74), .A2(new_n518), .B1(new_n509), .B2(KEYINPUT23), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n319), .A2(new_n320), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n199), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT74), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n519), .A2(new_n523), .B1(KEYINPUT23), .B2(new_n511), .ZN(new_n524));
  INV_X1    g338(.A(G110), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n517), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n519), .A2(new_n523), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n511), .A2(KEYINPUT23), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n529), .A2(KEYINPUT75), .A3(G110), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n516), .B1(new_n526), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n445), .A2(new_n465), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n524), .A2(new_n525), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n513), .B1(new_n510), .B2(new_n511), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n507), .B1(new_n531), .B2(new_n535), .ZN(new_n536));
  AOI22_X1  g350(.A1(new_n444), .A2(new_n445), .B1(new_n512), .B2(new_n514), .ZN(new_n537));
  AOI21_X1  g351(.A(KEYINPUT75), .B1(new_n529), .B2(G110), .ZN(new_n538));
  NOR3_X1   g352(.A1(new_n524), .A2(new_n517), .A3(new_n525), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n535), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(new_n541), .A3(new_n506), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n536), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(KEYINPUT25), .B1(new_n543), .B2(new_n300), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT25), .ZN(new_n545));
  AOI211_X1 g359(.A(new_n545), .B(G902), .C1(new_n536), .C2(new_n542), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n502), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n502), .A2(G902), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n543), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT72), .ZN(new_n551));
  INV_X1    g365(.A(new_n327), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n258), .A2(new_n251), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n456), .B1(G134), .B2(new_n243), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n246), .A2(new_n456), .B1(new_n245), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT69), .ZN(new_n556));
  OAI22_X1  g370(.A1(new_n227), .A2(new_n228), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n246), .A2(new_n456), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n554), .A2(new_n245), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n560), .A2(KEYINPUT69), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n552), .B(new_n553), .C1(new_n557), .C2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n563), .A2(KEYINPUT28), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n562), .A2(KEYINPUT71), .ZN(new_n565));
  AOI22_X1  g379(.A1(new_n237), .A2(new_n560), .B1(new_n258), .B2(new_n251), .ZN(new_n566));
  OR2_X1    g380(.A1(new_n566), .A2(new_n552), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n560), .A2(KEYINPUT69), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n555), .A2(new_n556), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(new_n237), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT71), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n570), .A2(new_n571), .A3(new_n552), .A4(new_n553), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n565), .A2(new_n567), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n564), .B1(new_n573), .B2(KEYINPUT28), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n446), .A2(G210), .ZN(new_n575));
  XOR2_X1   g389(.A(new_n575), .B(KEYINPUT27), .Z(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT26), .B(G101), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT70), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n570), .A2(new_n581), .A3(KEYINPUT30), .A4(new_n553), .ZN(new_n582));
  OAI211_X1 g396(.A(KEYINPUT30), .B(new_n553), .C1(new_n557), .C2(new_n561), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(KEYINPUT70), .B1(new_n566), .B2(KEYINPUT30), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n582), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n327), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n565), .A2(new_n572), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n587), .A2(new_n589), .A3(new_n579), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT31), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n588), .B1(new_n586), .B2(new_n327), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n593), .A2(KEYINPUT31), .A3(new_n579), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n580), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(G472), .A2(G902), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n551), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT32), .ZN(new_n599));
  OR2_X1    g413(.A1(new_n574), .A2(new_n579), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT31), .B1(new_n593), .B2(new_n579), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n583), .B(KEYINPUT70), .C1(KEYINPUT30), .C2(new_n566), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n552), .B1(new_n602), .B2(new_n582), .ZN(new_n603));
  NOR4_X1   g417(.A1(new_n603), .A2(new_n591), .A3(new_n588), .A4(new_n578), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n600), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n605), .A2(KEYINPUT72), .A3(new_n596), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n598), .A2(new_n599), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n592), .A2(new_n594), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n597), .B1(new_n608), .B2(new_n600), .ZN(new_n609));
  OAI21_X1  g423(.A(KEYINPUT73), .B1(new_n593), .B2(new_n579), .ZN(new_n610));
  AOI21_X1  g424(.A(KEYINPUT29), .B1(new_n574), .B2(new_n579), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT73), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n612), .B(new_n578), .C1(new_n603), .C2(new_n588), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n570), .A2(new_n553), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n565), .B(new_n572), .C1(new_n552), .C2(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n564), .B1(new_n616), .B2(KEYINPUT28), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n579), .A2(KEYINPUT29), .ZN(new_n618));
  AOI21_X1  g432(.A(G902), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n609), .A2(KEYINPUT32), .B1(new_n620), .B2(G472), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n550), .B1(new_n607), .B2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n309), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n623), .B1(new_n301), .B2(new_n306), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT97), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n624), .A2(new_n625), .A3(new_n499), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n501), .A2(new_n622), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(G101), .ZN(G3));
  NAND2_X1  g442(.A1(new_n307), .A2(new_n309), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n629), .A2(new_n550), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n381), .A2(KEYINPUT99), .ZN(new_n631));
  INV_X1    g445(.A(new_n498), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n378), .A2(KEYINPUT99), .A3(new_n381), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AOI22_X1  g449(.A1(new_n489), .A2(new_n495), .B1(G475), .B2(new_n479), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT33), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n418), .A2(new_n637), .A3(new_n420), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n416), .A2(KEYINPUT33), .A3(new_n417), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n638), .A2(G478), .A3(new_n300), .A4(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n421), .A2(new_n422), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n636), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n635), .A2(new_n437), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n598), .A2(new_n606), .ZN(new_n645));
  OAI21_X1  g459(.A(G472), .B1(new_n595), .B2(G902), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT98), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OAI211_X1 g462(.A(KEYINPUT98), .B(G472), .C1(new_n595), .C2(G902), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n645), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n630), .A2(new_n644), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT34), .B(G104), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G6));
  INV_X1    g467(.A(KEYINPUT100), .ZN(new_n654));
  INV_X1    g468(.A(new_n495), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n494), .B1(new_n493), .B2(new_n481), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n489), .A2(KEYINPUT100), .A3(new_n495), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n427), .A2(new_n429), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n659), .A2(new_n660), .A3(new_n480), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n635), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n630), .A2(new_n650), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G107), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT101), .B(KEYINPUT35), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G9));
  INV_X1    g480(.A(KEYINPUT102), .ZN(new_n667));
  INV_X1    g481(.A(new_n502), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n540), .A2(new_n541), .A3(new_n506), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n506), .B1(new_n540), .B2(new_n541), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n300), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n545), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n543), .A2(KEYINPUT25), .A3(new_n300), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n668), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n540), .A2(new_n541), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n506), .A2(KEYINPUT36), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n548), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n667), .B1(new_n674), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n547), .A2(KEYINPUT102), .A3(new_n678), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n501), .A2(new_n626), .A3(new_n650), .A4(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT37), .B(G110), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G12));
  NAND2_X1  g500(.A1(new_n607), .A2(new_n621), .ZN(new_n687));
  INV_X1    g501(.A(new_n635), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n434), .A2(G900), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n431), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n691), .B1(new_n479), .B2(G475), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n659), .A2(new_n660), .A3(new_n692), .ZN(new_n693));
  AND3_X1   g507(.A1(new_n680), .A2(new_n681), .A3(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n687), .A2(new_n624), .A3(new_n688), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G128), .ZN(G30));
  XNOR2_X1  g510(.A(new_n690), .B(KEYINPUT39), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n624), .A2(new_n697), .ZN(new_n698));
  OR2_X1    g512(.A1(new_n698), .A2(KEYINPUT40), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(KEYINPUT40), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n605), .A2(KEYINPUT32), .A3(new_n596), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n593), .A2(new_n578), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n300), .B1(new_n616), .B2(new_n579), .ZN(new_n703));
  OAI21_X1  g517(.A(G472), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  AND2_X1   g518(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n607), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n382), .B(KEYINPUT38), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n547), .A2(new_n678), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n636), .B1(new_n427), .B2(new_n429), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n708), .A2(new_n710), .A3(new_n632), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n706), .A2(new_n707), .A3(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n699), .A2(new_n700), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(KEYINPUT103), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(new_n187), .ZN(G45));
  AOI211_X1 g529(.A(new_n691), .B(new_n636), .C1(new_n640), .C2(new_n641), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n680), .A2(new_n681), .A3(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n687), .A2(new_n624), .A3(new_n688), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G146), .ZN(G48));
  AND3_X1   g533(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n299), .B1(new_n298), .B2(new_n300), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n720), .A2(new_n721), .A3(new_n623), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n622), .A2(new_n644), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(KEYINPUT41), .B(G113), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G15));
  NAND3_X1  g539(.A1(new_n622), .A2(new_n722), .A3(new_n662), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT104), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n622), .A2(new_n722), .A3(KEYINPUT104), .A4(new_n662), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G116), .ZN(G18));
  AND3_X1   g545(.A1(new_n680), .A2(new_n681), .A3(new_n497), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n722), .A2(new_n687), .A3(new_n688), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(KEYINPUT105), .B(G119), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(G21));
  OAI22_X1  g549(.A1(new_n601), .A2(new_n604), .B1(new_n579), .B2(new_n617), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n596), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n646), .A2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n550), .ZN(new_n739));
  AND3_X1   g553(.A1(new_n738), .A2(new_n739), .A3(new_n436), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT106), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n372), .A2(new_n377), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT99), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n743), .A3(new_n310), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n634), .A2(new_n744), .A3(new_n498), .A4(new_n709), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n740), .A2(new_n741), .A3(new_n722), .A4(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n738), .A2(new_n746), .A3(new_n739), .A4(new_n436), .ZN(new_n748));
  INV_X1    g562(.A(new_n722), .ZN(new_n749));
  OAI21_X1  g563(.A(KEYINPUT106), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G122), .ZN(G24));
  AND4_X1   g566(.A1(new_n646), .A2(new_n708), .A3(new_n716), .A4(new_n737), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n722), .A2(new_n688), .A3(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G125), .ZN(G27));
  NAND3_X1  g569(.A1(new_n378), .A2(new_n498), .A3(new_n381), .ZN(new_n756));
  AOI211_X1 g570(.A(new_n623), .B(new_n756), .C1(new_n301), .C2(new_n306), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n622), .A2(new_n757), .A3(new_n716), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT42), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n756), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n642), .A2(new_n690), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n762), .A2(new_n759), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n624), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n620), .A2(G472), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n599), .B1(new_n595), .B2(new_n597), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(new_n766), .A3(new_n701), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(KEYINPUT107), .A3(new_n739), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(KEYINPUT107), .B1(new_n767), .B2(new_n739), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n764), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n760), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G131), .ZN(G33));
  NAND3_X1  g587(.A1(new_n622), .A2(new_n757), .A3(new_n693), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G134), .ZN(G36));
  NAND3_X1  g589(.A1(new_n277), .A2(new_n282), .A3(new_n295), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n277), .A2(new_n289), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n776), .B1(new_n777), .B2(new_n282), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT45), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n299), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI211_X1 g594(.A(KEYINPUT45), .B(new_n776), .C1(new_n777), .C2(new_n282), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(KEYINPUT108), .A3(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(KEYINPUT108), .B1(new_n780), .B2(new_n781), .ZN(new_n784));
  OAI22_X1  g598(.A1(new_n783), .A2(new_n784), .B1(new_n299), .B2(new_n300), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT46), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(KEYINPUT109), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT109), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n778), .A2(new_n779), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(G469), .A3(new_n781), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT108), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n302), .B1(new_n792), .B2(new_n782), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n788), .B1(new_n793), .B2(KEYINPUT46), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n720), .B1(new_n793), .B2(KEYINPUT46), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n787), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n796), .A2(new_n309), .A3(new_n697), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n640), .A2(new_n641), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n636), .ZN(new_n799));
  XOR2_X1   g613(.A(new_n799), .B(KEYINPUT43), .Z(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n708), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n801), .A2(new_n650), .ZN(new_n802));
  OR3_X1    g616(.A1(new_n802), .A2(KEYINPUT110), .A3(KEYINPUT44), .ZN(new_n803));
  OAI21_X1  g617(.A(KEYINPUT110), .B1(new_n802), .B2(KEYINPUT44), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n756), .B1(new_n802), .B2(KEYINPUT44), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n797), .A2(new_n803), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G137), .ZN(G39));
  NOR4_X1   g621(.A1(new_n687), .A2(new_n739), .A3(new_n762), .A4(new_n756), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n796), .A2(KEYINPUT47), .A3(new_n309), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT47), .B1(new_n796), .B2(new_n309), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n808), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G140), .ZN(G42));
  NOR2_X1   g626(.A1(new_n720), .A2(new_n721), .ZN(new_n813));
  XOR2_X1   g627(.A(new_n813), .B(KEYINPUT49), .Z(new_n814));
  OR4_X1    g628(.A1(new_n550), .A2(new_n799), .A3(new_n623), .A4(new_n632), .ZN(new_n815));
  OR4_X1    g629(.A1(new_n706), .A2(new_n814), .A3(new_n707), .A4(new_n815), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n723), .A2(new_n733), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n730), .A2(new_n751), .A3(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n660), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n819), .A2(new_n659), .A3(new_n692), .ZN(new_n820));
  AOI211_X1 g634(.A(new_n820), .B(new_n682), .C1(new_n607), .C2(new_n621), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n757), .B1(new_n821), .B2(new_n753), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n772), .A2(new_n822), .A3(new_n774), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n818), .A2(new_n823), .ZN(new_n824));
  XOR2_X1   g638(.A(new_n690), .B(KEYINPUT114), .Z(new_n825));
  NAND3_X1  g639(.A1(new_n547), .A2(new_n678), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n745), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n706), .A2(new_n624), .A3(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n695), .A2(new_n718), .A3(new_n828), .A4(new_n754), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n829), .A2(KEYINPUT52), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n695), .A2(new_n754), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT113), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n695), .A2(new_n754), .A3(KEYINPUT113), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n833), .A2(new_n718), .A3(new_n828), .A4(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n830), .B1(new_n835), .B2(KEYINPUT52), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n632), .B1(new_n378), .B2(new_n381), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n436), .A3(new_n642), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT111), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n660), .A2(new_n636), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n837), .A2(new_n840), .A3(new_n436), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT111), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n837), .A2(new_n842), .A3(new_n436), .A4(new_n642), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n839), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n630), .A2(new_n650), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n684), .A2(new_n627), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT112), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n684), .A2(new_n627), .A3(new_n845), .A4(KEYINPUT112), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n824), .A2(new_n836), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n851), .A2(KEYINPUT115), .A3(new_n852), .ZN(new_n853));
  XOR2_X1   g667(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT52), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n829), .B(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n824), .A2(new_n850), .A3(new_n855), .A4(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n853), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT115), .B1(new_n851), .B2(new_n852), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT54), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n769), .A2(new_n770), .ZN(new_n862));
  INV_X1    g676(.A(new_n431), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n800), .A2(new_n722), .A3(new_n863), .A4(new_n761), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  XOR2_X1   g679(.A(new_n865), .B(KEYINPUT48), .Z(new_n866));
  INV_X1    g680(.A(G952), .ZN(new_n867));
  AND4_X1   g681(.A1(new_n739), .A2(new_n800), .A3(new_n863), .A4(new_n738), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n749), .A2(new_n635), .ZN(new_n869));
  AOI211_X1 g683(.A(new_n867), .B(G953), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n722), .A2(new_n761), .ZN(new_n871));
  OR4_X1    g685(.A1(new_n550), .A2(new_n871), .A3(new_n431), .A4(new_n706), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n866), .B(new_n870), .C1(new_n643), .C2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n707), .A2(new_n498), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n868), .A2(new_n722), .A3(new_n874), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT50), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n640), .A2(new_n636), .A3(new_n641), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n738), .A2(new_n708), .ZN(new_n878));
  OAI22_X1  g692(.A1(new_n872), .A2(new_n877), .B1(new_n878), .B2(new_n864), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n720), .A2(new_n721), .A3(new_n309), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n809), .A2(new_n810), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n868), .A2(new_n761), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n880), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(KEYINPUT51), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT51), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n880), .B(new_n886), .C1(new_n882), .C2(new_n883), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n873), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n730), .A2(new_n751), .A3(new_n817), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n772), .A2(new_n774), .A3(new_n822), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n850), .A2(new_n857), .A3(new_n889), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n854), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT54), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n824), .A2(new_n836), .A3(KEYINPUT53), .A4(new_n850), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n861), .A2(new_n888), .A3(KEYINPUT117), .A4(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n867), .A2(new_n279), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n895), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n850), .A2(new_n890), .A3(new_n889), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n835), .A2(KEYINPUT52), .ZN(new_n901));
  INV_X1    g715(.A(new_n830), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n852), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT115), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(new_n858), .A3(new_n853), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n899), .B1(new_n907), .B2(KEYINPUT54), .ZN(new_n908));
  AOI21_X1  g722(.A(KEYINPUT117), .B1(new_n908), .B2(new_n888), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n816), .B1(new_n898), .B2(new_n909), .ZN(G75));
  NAND2_X1  g724(.A1(new_n344), .A2(new_n353), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(new_n351), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT55), .Z(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n300), .B1(new_n892), .B2(new_n894), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(G210), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT56), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT119), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n279), .A2(G952), .ZN(new_n921));
  XNOR2_X1  g735(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n913), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n921), .B1(new_n916), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n919), .A2(new_n920), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n916), .A2(new_n923), .ZN(new_n926));
  INV_X1    g740(.A(new_n921), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT119), .B1(new_n928), .B2(new_n918), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n925), .A2(new_n929), .ZN(G51));
  NAND2_X1  g744(.A1(new_n892), .A2(new_n894), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n931), .A2(G902), .A3(new_n792), .A4(new_n782), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT121), .Z(new_n933));
  XNOR2_X1  g747(.A(new_n931), .B(new_n893), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n302), .B(KEYINPUT120), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT57), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n298), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n921), .B1(new_n933), .B2(new_n937), .ZN(G54));
  AND3_X1   g752(.A1(new_n915), .A2(KEYINPUT58), .A3(G475), .ZN(new_n939));
  OAI21_X1  g753(.A(KEYINPUT122), .B1(new_n939), .B2(new_n493), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n921), .B1(new_n939), .B2(new_n493), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n939), .A2(KEYINPUT122), .A3(new_n493), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n942), .A2(new_n943), .ZN(G60));
  NAND2_X1  g758(.A1(G478), .A2(G902), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT59), .Z(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n638), .A2(new_n639), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n927), .B1(new_n934), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n638), .A2(new_n639), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n861), .A2(new_n895), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n947), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n949), .B1(new_n950), .B2(new_n952), .ZN(G63));
  XNOR2_X1  g767(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n413), .A2(new_n300), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n954), .B(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n931), .A2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n543), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n921), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n956), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n892), .B2(new_n894), .ZN(new_n961));
  AND3_X1   g775(.A1(new_n961), .A2(KEYINPUT124), .A3(new_n677), .ZN(new_n962));
  AOI21_X1  g776(.A(KEYINPUT124), .B1(new_n961), .B2(new_n677), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n959), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT125), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n965), .B1(new_n962), .B2(new_n963), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT61), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n964), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  OAI221_X1 g782(.A(new_n959), .B1(new_n965), .B2(KEYINPUT61), .C1(new_n962), .C2(new_n963), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(G66));
  INV_X1    g784(.A(G224), .ZN(new_n971));
  OAI21_X1  g785(.A(G953), .B1(new_n432), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n850), .A2(new_n889), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n972), .B1(new_n974), .B2(G953), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n911), .B1(G898), .B2(new_n279), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT126), .Z(new_n977));
  XNOR2_X1  g791(.A(new_n975), .B(new_n977), .ZN(G69));
  AOI21_X1  g792(.A(new_n279), .B1(G227), .B2(G900), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n811), .A2(new_n806), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n797), .B(new_n746), .C1(new_n770), .C2(new_n769), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n772), .A2(new_n774), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n833), .A2(new_n718), .A3(new_n834), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n980), .A2(new_n981), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n482), .B1(new_n483), .B2(KEYINPUT19), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n586), .B(new_n986), .Z(new_n987));
  NAND3_X1  g801(.A1(new_n985), .A2(new_n279), .A3(new_n987), .ZN(new_n988));
  OR3_X1    g802(.A1(new_n840), .A2(KEYINPUT127), .A3(new_n642), .ZN(new_n989));
  OAI21_X1  g803(.A(KEYINPUT127), .B1(new_n840), .B2(new_n642), .ZN(new_n990));
  AND3_X1   g804(.A1(new_n989), .A2(new_n761), .A3(new_n990), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n991), .A2(new_n622), .A3(new_n624), .A4(new_n697), .ZN(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT62), .ZN(new_n994));
  OR3_X1    g808(.A1(new_n714), .A2(new_n994), .A3(new_n983), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n994), .B1(new_n714), .B2(new_n983), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n993), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(G953), .B1(new_n997), .B2(new_n980), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n988), .B1(new_n998), .B2(new_n987), .ZN(new_n999));
  INV_X1    g813(.A(G900), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n979), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n1001), .B1(new_n979), .B2(new_n999), .ZN(G72));
  NAND2_X1  g816(.A1(G472), .A2(G902), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1003), .B(KEYINPUT63), .Z(new_n1004));
  OAI21_X1  g818(.A(new_n1004), .B1(new_n985), .B2(new_n973), .ZN(new_n1005));
  NOR3_X1   g819(.A1(new_n603), .A2(new_n588), .A3(new_n579), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n921), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n997), .A2(new_n974), .A3(new_n980), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1008), .A2(new_n1004), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(new_n702), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n610), .A2(new_n590), .A3(new_n613), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n907), .A2(new_n1004), .A3(new_n1011), .ZN(new_n1012));
  AND3_X1   g826(.A1(new_n1007), .A2(new_n1010), .A3(new_n1012), .ZN(G57));
endmodule


