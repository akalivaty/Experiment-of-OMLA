//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 0 1 0 1 1 0 1 0 0 0 1 1 1 1 0 1 1 1 1 0 1 1 0 0 0 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1216, new_n1217, new_n1218,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1282, new_n1283, new_n1284;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  XOR2_X1   g0017(.A(KEYINPUT64), .B(G238), .Z(new_n218));
  INV_X1    g0018(.A(G68), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G107), .A2(G264), .ZN(new_n224));
  NAND4_X1  g0024(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n209), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n202), .A2(G68), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n219), .A2(G50), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n240), .B(new_n245), .ZN(G351));
  NAND3_X1  g0046(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n219), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT12), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  AOI22_X1  g0051(.A1(new_n251), .A2(G50), .B1(G20), .B2(new_n219), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(G20), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G77), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n252), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n215), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n257), .A2(KEYINPUT11), .A3(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n248), .A2(new_n259), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n206), .A2(G20), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n261), .A2(G68), .A3(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n250), .A2(new_n260), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(KEYINPUT11), .B1(new_n257), .B2(new_n259), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT14), .ZN(new_n268));
  INV_X1    g0068(.A(G41), .ZN(new_n269));
  INV_X1    g0069(.A(G45), .ZN(new_n270));
  AOI21_X1  g0070(.A(G1), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n272), .A2(G1), .A3(G13), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n271), .A2(new_n273), .A3(G274), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G238), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n274), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(new_n278), .B(KEYINPUT68), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT3), .B(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n230), .A2(G1698), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n280), .B(new_n281), .C1(G226), .C2(G1698), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G33), .A2(G97), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT67), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n273), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n282), .A2(KEYINPUT67), .A3(new_n283), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT13), .ZN(new_n290));
  AND3_X1   g0090(.A1(new_n279), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n290), .B1(new_n279), .B2(new_n289), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n268), .B(G169), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n279), .A2(new_n289), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT13), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n279), .A2(new_n289), .A3(new_n290), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n295), .A2(G179), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(new_n296), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n268), .B1(new_n299), .B2(G169), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n267), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT69), .ZN(new_n302));
  OAI21_X1  g0102(.A(G200), .B1(new_n291), .B2(new_n292), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n295), .A2(G190), .A3(new_n296), .ZN(new_n304));
  AND3_X1   g0104(.A1(new_n303), .A2(new_n304), .A3(new_n266), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  AND3_X1   g0106(.A1(new_n301), .A2(new_n302), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n302), .B1(new_n301), .B2(new_n306), .ZN(new_n308));
  INV_X1    g0108(.A(G226), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n274), .B1(new_n276), .B2(new_n309), .ZN(new_n310));
  OR2_X1    g0110(.A1(KEYINPUT3), .A2(G33), .ZN(new_n311));
  NAND2_X1  g0111(.A1(KEYINPUT3), .A2(G33), .ZN(new_n312));
  AOI21_X1  g0112(.A(G1698), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  AND2_X1   g0113(.A1(KEYINPUT3), .A2(G33), .ZN(new_n314));
  NOR2_X1   g0114(.A1(KEYINPUT3), .A2(G33), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n313), .A2(G222), .B1(new_n316), .B2(G77), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n280), .A2(G1698), .ZN(new_n318));
  XOR2_X1   g0118(.A(KEYINPUT65), .B(G223), .Z(new_n319));
  OAI21_X1  g0119(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n310), .B1(new_n320), .B2(new_n287), .ZN(new_n321));
  XOR2_X1   g0121(.A(KEYINPUT66), .B(G200), .Z(new_n322));
  OR2_X1    g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n261), .A2(G50), .A3(new_n262), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(G50), .B2(new_n247), .ZN(new_n325));
  INV_X1    g0125(.A(new_n259), .ZN(new_n326));
  XOR2_X1   g0126(.A(KEYINPUT8), .B(G58), .Z(new_n327));
  AOI22_X1  g0127(.A1(new_n327), .A2(new_n254), .B1(G150), .B2(new_n251), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n203), .A2(G20), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n326), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  OR2_X1    g0131(.A1(new_n331), .A2(KEYINPUT9), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n321), .A2(G190), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n331), .A2(KEYINPUT9), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n323), .A2(new_n332), .A3(new_n333), .A4(new_n334), .ZN(new_n335));
  OR2_X1    g0135(.A1(new_n335), .A2(KEYINPUT10), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(KEYINPUT10), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G244), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n274), .B1(new_n276), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G1698), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n280), .A2(G232), .A3(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(G107), .ZN(new_n343));
  OAI221_X1 g0143(.A(new_n342), .B1(new_n343), .B2(new_n280), .C1(new_n318), .C2(new_n218), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n340), .B1(new_n344), .B2(new_n287), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n345), .A2(G169), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n261), .A2(G77), .A3(new_n262), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(G77), .B2(new_n247), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n327), .A2(new_n251), .B1(G20), .B2(G77), .ZN(new_n349));
  XOR2_X1   g0149(.A(KEYINPUT15), .B(G87), .Z(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n254), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n326), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n346), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G179), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n345), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n345), .A2(G190), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n358), .B(new_n353), .C1(new_n322), .C2(new_n345), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n321), .A2(new_n355), .ZN(new_n360));
  OAI221_X1 g0160(.A(new_n360), .B1(G169), .B2(new_n321), .C1(new_n330), .C2(new_n325), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n338), .A2(new_n357), .A3(new_n359), .A4(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT17), .ZN(new_n363));
  XNOR2_X1  g0163(.A(KEYINPUT8), .B(G58), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n364), .B1(new_n206), .B2(G20), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n365), .A2(new_n261), .B1(new_n248), .B2(new_n364), .ZN(new_n366));
  AOI21_X1  g0166(.A(KEYINPUT7), .B1(new_n316), .B2(new_n207), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n311), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n312), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(G68), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(G58), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n371), .A2(new_n219), .ZN(new_n372));
  OAI21_X1  g0172(.A(G20), .B1(new_n372), .B2(new_n201), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n251), .A2(G159), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(KEYINPUT16), .B1(new_n370), .B2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n311), .A2(new_n207), .A3(new_n312), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT7), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n219), .B1(new_n380), .B2(new_n368), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n373), .A2(KEYINPUT16), .A3(new_n374), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n259), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n366), .B1(new_n377), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n309), .A2(G1698), .ZN(new_n385));
  OAI221_X1 g0185(.A(new_n385), .B1(G223), .B2(G1698), .C1(new_n314), .C2(new_n315), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G33), .A2(G87), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n273), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n274), .B1(new_n276), .B2(new_n230), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(G190), .ZN(new_n391));
  AND2_X1   g0191(.A1(new_n391), .A2(KEYINPUT72), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n391), .A2(KEYINPUT72), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(G200), .B1(new_n388), .B2(new_n389), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI211_X1 g0198(.A(KEYINPUT73), .B(new_n363), .C1(new_n384), .C2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n397), .ZN(new_n400));
  NOR3_X1   g0200(.A1(new_n388), .A2(new_n389), .A3(new_n394), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n366), .ZN(new_n403));
  INV_X1    g0203(.A(new_n382), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n326), .B1(new_n370), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT16), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(new_n381), .B2(new_n375), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n403), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  OR2_X1    g0208(.A1(new_n363), .A2(KEYINPUT73), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n363), .A2(KEYINPUT73), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n402), .A2(new_n408), .A3(new_n409), .A4(new_n410), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n399), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT70), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n384), .A2(new_n413), .ZN(new_n414));
  OAI211_X1 g0214(.A(KEYINPUT70), .B(new_n366), .C1(new_n377), .C2(new_n383), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n390), .A2(G179), .ZN(new_n416));
  INV_X1    g0216(.A(G169), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n416), .B1(new_n417), .B2(new_n390), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n414), .A2(new_n415), .A3(new_n418), .ZN(new_n419));
  XOR2_X1   g0219(.A(KEYINPUT71), .B(KEYINPUT18), .Z(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NOR2_X1   g0221(.A1(KEYINPUT71), .A2(KEYINPUT18), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n414), .A2(new_n415), .A3(new_n418), .A4(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n412), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  NOR4_X1   g0224(.A1(new_n307), .A2(new_n308), .A3(new_n362), .A4(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT81), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT20), .ZN(new_n427));
  INV_X1    g0227(.A(G97), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n207), .B1(new_n428), .B2(G33), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT75), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n430), .A2(G33), .A3(G283), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G33), .A2(G283), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT75), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n429), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(G116), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n258), .A2(new_n215), .B1(G20), .B2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n427), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n433), .A2(new_n431), .ZN(new_n439));
  OAI211_X1 g0239(.A(KEYINPUT20), .B(new_n436), .C1(new_n439), .C2(new_n429), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n247), .A2(G116), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n253), .A2(G1), .ZN(new_n443));
  NOR3_X1   g0243(.A1(new_n248), .A2(new_n259), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n442), .B1(new_n444), .B2(G116), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n417), .B1(new_n441), .B2(new_n445), .ZN(new_n446));
  OAI211_X1 g0246(.A(G264), .B(G1698), .C1(new_n314), .C2(new_n315), .ZN(new_n447));
  OAI211_X1 g0247(.A(G257), .B(new_n341), .C1(new_n314), .C2(new_n315), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n311), .A2(G303), .A3(new_n312), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  AND2_X1   g0250(.A1(new_n450), .A2(new_n287), .ZN(new_n451));
  XNOR2_X1  g0251(.A(KEYINPUT5), .B(G41), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n206), .A2(G45), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n455), .A2(G270), .A3(new_n273), .ZN(new_n456));
  OR2_X1    g0256(.A1(KEYINPUT5), .A2(G41), .ZN(new_n457));
  NAND2_X1  g0257(.A1(KEYINPUT5), .A2(G41), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n453), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(G274), .ZN(new_n460));
  INV_X1    g0260(.A(new_n215), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n460), .B1(new_n461), .B2(new_n272), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n456), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(KEYINPUT80), .B1(new_n451), .B2(new_n464), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n452), .A2(new_n454), .B1(new_n461), .B2(new_n272), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n466), .A2(G270), .B1(new_n459), .B2(new_n462), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n450), .A2(new_n287), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT80), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n446), .A2(new_n465), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT21), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n441), .A2(new_n445), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n467), .A2(new_n468), .A3(G179), .ZN(new_n475));
  OR2_X1    g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n446), .A2(new_n465), .A3(KEYINPUT21), .A4(new_n470), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n473), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n470), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n469), .B1(new_n467), .B2(new_n468), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n395), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n465), .A2(G200), .A3(new_n470), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n481), .A2(new_n474), .A3(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n426), .B1(new_n478), .B2(new_n483), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n476), .A2(new_n477), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n481), .A2(new_n482), .A3(new_n474), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n485), .A2(KEYINPUT81), .A3(new_n473), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT77), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n251), .A2(G77), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT6), .ZN(new_n492));
  AND2_X1   g0292(.A1(G97), .A2(G107), .ZN(new_n493));
  NOR2_X1   g0293(.A1(G97), .A2(G107), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n343), .A2(KEYINPUT6), .A3(G97), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n491), .B1(new_n497), .B2(G20), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n380), .A2(new_n368), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n498), .A2(KEYINPUT74), .B1(new_n499), .B2(G107), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT74), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n207), .B1(new_n495), .B2(new_n496), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n501), .B1(new_n502), .B2(new_n491), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n326), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n247), .A2(G97), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n505), .B1(new_n444), .B2(G97), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n489), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n498), .A2(KEYINPUT74), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n499), .A2(G107), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n509), .A2(new_n503), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n259), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n512), .A2(KEYINPUT77), .A3(new_n506), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n455), .A2(G257), .A3(new_n273), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n463), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  OAI211_X1 g0316(.A(G244), .B(new_n341), .C1(new_n314), .C2(new_n315), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT4), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n280), .A2(KEYINPUT4), .A3(G244), .A4(new_n341), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n433), .A2(new_n431), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n280), .A2(G250), .A3(G1698), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n519), .A2(new_n520), .A3(new_n521), .A4(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT76), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n523), .A2(new_n524), .A3(new_n287), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n524), .B1(new_n523), .B2(new_n287), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n355), .B(new_n516), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n515), .B1(new_n287), .B2(new_n523), .ZN(new_n529));
  OR2_X1    g0329(.A1(new_n529), .A2(G169), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n508), .A2(new_n513), .A3(new_n528), .A4(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n504), .A2(new_n507), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n529), .A2(G190), .ZN(new_n533));
  INV_X1    g0333(.A(new_n527), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n515), .B1(new_n534), .B2(new_n525), .ZN(new_n535));
  INV_X1    g0335(.A(G200), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n532), .B(new_n533), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(G244), .B(G1698), .C1(new_n314), .C2(new_n315), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT78), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT78), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n280), .A2(new_n540), .A3(G244), .A4(G1698), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n280), .A2(G238), .A3(new_n341), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n253), .A2(new_n435), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n539), .A2(new_n541), .A3(new_n542), .A4(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT79), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n543), .B1(new_n313), .B2(G238), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n548), .A2(KEYINPUT79), .A3(new_n541), .A4(new_n539), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n287), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n462), .A2(new_n454), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n273), .A2(G250), .A3(new_n453), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n550), .A2(new_n355), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n254), .A2(G97), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT19), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n207), .B1(new_n283), .B2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(G87), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n494), .A2(new_n559), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n556), .A2(new_n557), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n280), .A2(new_n207), .A3(G68), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n259), .ZN(new_n564));
  INV_X1    g0364(.A(new_n350), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n248), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n444), .A2(new_n350), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n273), .B1(new_n545), .B2(new_n546), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n553), .B1(new_n571), .B2(new_n549), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n555), .B(new_n570), .C1(G169), .C2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n550), .A2(G190), .A3(new_n554), .ZN(new_n574));
  INV_X1    g0374(.A(new_n444), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n575), .A2(new_n559), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n567), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n574), .B(new_n577), .C1(new_n572), .C2(new_n322), .ZN(new_n578));
  AND4_X1   g0378(.A1(new_n531), .A2(new_n537), .A3(new_n573), .A4(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n559), .A2(KEYINPUT82), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n280), .A2(new_n207), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT22), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n280), .A2(KEYINPUT22), .A3(new_n207), .A4(new_n580), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT23), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n207), .B2(G107), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n343), .A2(KEYINPUT23), .A3(G20), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n586), .A2(new_n587), .B1(new_n543), .B2(new_n207), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n583), .A2(new_n584), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT24), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT24), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n583), .A2(new_n591), .A3(new_n584), .A4(new_n588), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n326), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(KEYINPUT25), .B1(new_n248), .B2(new_n343), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n248), .A2(KEYINPUT25), .A3(new_n343), .ZN(new_n595));
  OAI22_X1  g0395(.A1(new_n575), .A2(new_n343), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n313), .A2(G250), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n280), .A2(G257), .A3(G1698), .ZN(new_n599));
  NAND2_X1  g0399(.A1(G33), .A2(G294), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n601), .A2(new_n287), .B1(G264), .B2(new_n466), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n602), .A2(G190), .A3(new_n463), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n463), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(G200), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n597), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(new_n417), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n602), .A2(new_n355), .A3(new_n463), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n607), .B(new_n608), .C1(new_n593), .C2(new_n596), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n425), .A2(new_n488), .A3(new_n579), .A4(new_n610), .ZN(new_n611));
  XOR2_X1   g0411(.A(new_n611), .B(KEYINPUT83), .Z(G372));
  NAND2_X1  g0412(.A1(new_n578), .A2(new_n573), .ZN(new_n613));
  OAI21_X1  g0413(.A(KEYINPUT26), .B1(new_n613), .B2(new_n531), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n609), .A2(new_n473), .A3(new_n476), .A4(new_n477), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n606), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n531), .A2(new_n537), .A3(new_n573), .A4(new_n578), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n614), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n573), .A2(KEYINPUT84), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n550), .A2(new_n554), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n417), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT84), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n622), .A2(new_n623), .A3(new_n555), .A4(new_n570), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n528), .A2(new_n530), .ZN(new_n625));
  INV_X1    g0425(.A(new_n532), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n625), .A2(new_n573), .A3(new_n578), .A4(new_n626), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n620), .B(new_n624), .C1(new_n627), .C2(KEYINPUT26), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n619), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n425), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT85), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n338), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n336), .A2(KEYINPUT85), .A3(new_n337), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n412), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n305), .A2(new_n357), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n636), .B1(new_n637), .B2(new_n301), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n418), .A2(new_n384), .ZN(new_n639));
  OR2_X1    g0439(.A1(new_n639), .A2(KEYINPUT18), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(KEYINPUT18), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n635), .B1(new_n638), .B2(new_n642), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n643), .A2(new_n361), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n631), .A2(new_n644), .ZN(G369));
  NAND3_X1  g0445(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(G213), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(G343), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n474), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT86), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n653), .B1(new_n488), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n484), .A2(new_n487), .A3(KEYINPUT86), .ZN(new_n656));
  INV_X1    g0456(.A(new_n478), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n655), .A2(new_n656), .B1(new_n657), .B2(new_n653), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n651), .B1(new_n593), .B2(new_n596), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT87), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(new_n606), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n609), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n609), .A2(new_n651), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n658), .A2(G330), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n478), .A2(new_n652), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n664), .A2(new_n671), .A3(new_n666), .ZN(new_n672));
  AOI21_X1  g0472(.A(KEYINPUT88), .B1(new_n672), .B2(new_n666), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n672), .A2(KEYINPUT88), .A3(new_n666), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n669), .B1(new_n673), .B2(new_n674), .ZN(G399));
  INV_X1    g0475(.A(new_n210), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(G41), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n560), .A2(G116), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(G1), .A3(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(new_n213), .B2(new_n678), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT28), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n578), .A2(new_n573), .ZN(new_n683));
  INV_X1    g0483(.A(new_n531), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT26), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n627), .A2(KEYINPUT26), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n686), .B(new_n687), .C1(new_n617), .C2(new_n616), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n620), .A2(new_n624), .A3(KEYINPUT90), .ZN(new_n689));
  AOI21_X1  g0489(.A(KEYINPUT90), .B1(new_n620), .B2(new_n624), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI211_X1 g0491(.A(KEYINPUT29), .B(new_n652), .C1(new_n688), .C2(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n651), .B1(new_n619), .B2(new_n629), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n692), .B1(new_n693), .B2(KEYINPUT29), .ZN(new_n694));
  INV_X1    g0494(.A(G330), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT30), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n475), .A2(KEYINPUT89), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT89), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n467), .A2(new_n468), .A3(new_n698), .A4(G179), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n550), .A2(new_n529), .A3(new_n554), .A4(new_n602), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n696), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n529), .A2(new_n602), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n697), .A2(new_n699), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n703), .A2(new_n704), .A3(KEYINPUT30), .A4(new_n572), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n516), .B1(new_n526), .B2(new_n527), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n479), .A2(new_n480), .ZN(new_n707));
  AOI21_X1  g0507(.A(G179), .B1(new_n602), .B2(new_n463), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n706), .A2(new_n707), .A3(new_n621), .A4(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n702), .A2(new_n705), .A3(new_n709), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n710), .A2(KEYINPUT31), .A3(new_n651), .ZN(new_n711));
  AOI21_X1  g0511(.A(KEYINPUT31), .B1(new_n710), .B2(new_n651), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n488), .A2(new_n579), .A3(new_n610), .A4(new_n652), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n695), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n694), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n682), .B1(new_n717), .B2(G1), .ZN(G364));
  NAND2_X1  g0518(.A1(new_n658), .A2(G330), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n207), .A2(G13), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT91), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(G45), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n678), .A2(G1), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n719), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n658), .A2(G330), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(G13), .A2(G33), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(G20), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n658), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n676), .A2(new_n316), .ZN(new_n732));
  AOI22_X1  g0532(.A1(new_n732), .A2(G355), .B1(new_n435), .B2(new_n676), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n676), .A2(new_n280), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(G45), .B2(new_n213), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n245), .A2(new_n270), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n733), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n215), .B1(G20), .B2(new_n417), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n729), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n723), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g0540(.A(new_n740), .B(KEYINPUT92), .ZN(new_n741));
  INV_X1    g0541(.A(new_n738), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n207), .A2(G190), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G179), .A2(G200), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n280), .B1(new_n746), .B2(G329), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n207), .A2(new_n355), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n536), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G190), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(G311), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n394), .A2(new_n749), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(G322), .ZN(new_n755));
  OAI221_X1 g0555(.A(new_n747), .B1(new_n751), .B2(new_n752), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n748), .A2(G200), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n394), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(G326), .ZN(new_n760));
  INV_X1    g0560(.A(G294), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n744), .A2(G190), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G20), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n759), .A2(new_n760), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n756), .B1(KEYINPUT94), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n757), .A2(G190), .ZN(new_n767));
  XNOR2_X1  g0567(.A(KEYINPUT33), .B(G317), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT95), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n770), .B1(new_n769), .B2(new_n768), .ZN(new_n771));
  INV_X1    g0571(.A(G283), .ZN(new_n772));
  INV_X1    g0572(.A(new_n322), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n773), .A2(new_n355), .A3(new_n743), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n207), .A2(new_n391), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n773), .A2(new_n355), .A3(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G303), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n772), .A2(new_n774), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n771), .A2(new_n778), .ZN(new_n779));
  OAI211_X1 g0579(.A(new_n766), .B(new_n779), .C1(KEYINPUT94), .C2(new_n765), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n759), .A2(new_n202), .ZN(new_n781));
  INV_X1    g0581(.A(new_n767), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n746), .A2(G159), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n782), .A2(new_n219), .B1(new_n783), .B2(KEYINPUT32), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n781), .B(new_n784), .C1(KEYINPUT32), .C2(new_n783), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n280), .B1(new_n764), .B2(new_n428), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n776), .A2(new_n559), .ZN(new_n787));
  INV_X1    g0587(.A(new_n774), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n786), .B(new_n787), .C1(G107), .C2(new_n788), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n753), .A2(G58), .B1(new_n750), .B2(G77), .ZN(new_n790));
  OR2_X1    g0590(.A1(new_n790), .A2(KEYINPUT93), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(KEYINPUT93), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n785), .A2(new_n789), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n742), .B1(new_n780), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n741), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n726), .B1(new_n731), .B2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(G396));
  INV_X1    g0597(.A(new_n723), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n359), .B1(new_n353), .B2(new_n652), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(new_n357), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n357), .A2(new_n651), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n803), .B(new_n652), .C1(new_n618), .C2(new_n628), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n803), .B(KEYINPUT99), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n804), .B1(new_n693), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n798), .B1(new_n806), .B2(new_n716), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n716), .B2(new_n806), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n738), .A2(new_n727), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT96), .Z(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n723), .B1(new_n256), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n788), .A2(G87), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n752), .B2(new_n745), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  AND2_X1   g0615(.A1(new_n815), .A2(KEYINPUT98), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n815), .A2(KEYINPUT98), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n280), .B1(new_n763), .B2(G97), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n818), .B1(new_n776), .B2(new_n343), .C1(new_n761), .C2(new_n754), .ZN(new_n819));
  NOR3_X1   g0619(.A1(new_n816), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n758), .A2(G303), .B1(new_n767), .B2(G283), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n435), .B2(new_n751), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n822), .B(KEYINPUT97), .Z(new_n823));
  AOI22_X1  g0623(.A1(new_n758), .A2(G137), .B1(new_n750), .B2(G159), .ZN(new_n824));
  INV_X1    g0624(.A(G143), .ZN(new_n825));
  INV_X1    g0625(.A(G150), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n824), .B1(new_n825), .B2(new_n754), .C1(new_n826), .C2(new_n782), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT34), .ZN(new_n828));
  INV_X1    g0628(.A(G132), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n280), .B1(new_n745), .B2(new_n829), .C1(new_n764), .C2(new_n371), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n776), .A2(new_n202), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n830), .B(new_n831), .C1(G68), .C2(new_n788), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n820), .A2(new_n823), .B1(new_n828), .B2(new_n832), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n812), .B1(new_n833), .B2(new_n742), .C1(new_n803), .C2(new_n728), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n808), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(G384));
  INV_X1    g0636(.A(KEYINPUT38), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT37), .ZN(new_n838));
  INV_X1    g0638(.A(new_n649), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n414), .A2(new_n415), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(KEYINPUT101), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT101), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n414), .A2(new_n415), .A3(new_n842), .A4(new_n839), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n402), .A2(new_n408), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n639), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n838), .B1(new_n844), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n419), .A2(new_n838), .A3(new_n845), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(new_n843), .B2(new_n841), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n642), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n844), .B1(new_n852), .B2(new_n412), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n837), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n408), .A2(new_n649), .ZN(new_n855));
  OAI21_X1  g0655(.A(KEYINPUT37), .B1(new_n846), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n844), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n856), .B1(new_n857), .B2(new_n849), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT100), .ZN(new_n859));
  AND3_X1   g0659(.A1(new_n424), .A2(new_n859), .A3(new_n855), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n859), .B1(new_n424), .B2(new_n855), .ZN(new_n861));
  OAI211_X1 g0661(.A(KEYINPUT38), .B(new_n858), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n854), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT39), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n858), .B1(new_n860), .B2(new_n861), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n837), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n867), .A2(KEYINPUT39), .A3(new_n862), .ZN(new_n868));
  OAI21_X1  g0668(.A(G169), .B1(new_n291), .B2(new_n292), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(KEYINPUT14), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n870), .A2(new_n297), .A3(new_n293), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n871), .A2(new_n267), .A3(new_n652), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n865), .A2(new_n868), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n867), .A2(new_n862), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n267), .A2(new_n651), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n301), .A2(new_n306), .A3(new_n876), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n267), .B(new_n651), .C1(new_n871), .C2(new_n305), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n802), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n879), .B1(new_n804), .B2(new_n880), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n875), .A2(new_n881), .B1(new_n642), .B2(new_n649), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n874), .A2(new_n882), .ZN(new_n883));
  XOR2_X1   g0683(.A(new_n883), .B(KEYINPUT102), .Z(new_n884));
  OAI211_X1 g0684(.A(new_n425), .B(new_n692), .C1(KEYINPUT29), .C2(new_n693), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n644), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n884), .B(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n713), .A2(new_n714), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n877), .A2(new_n878), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n888), .A2(new_n803), .A3(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT103), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(KEYINPUT103), .A2(KEYINPUT40), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n892), .B(new_n875), .C1(new_n890), .C2(new_n893), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n854), .A2(new_n862), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT40), .B1(new_n895), .B2(new_n890), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  AND3_X1   g0697(.A1(new_n897), .A2(new_n425), .A3(new_n888), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n897), .B1(new_n425), .B2(new_n888), .ZN(new_n899));
  NOR3_X1   g0699(.A1(new_n898), .A2(new_n899), .A3(new_n695), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n887), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n887), .A2(new_n900), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n206), .B2(new_n721), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n901), .B1(new_n903), .B2(KEYINPUT104), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(KEYINPUT104), .B2(new_n903), .ZN(new_n905));
  OR2_X1    g0705(.A1(new_n497), .A2(KEYINPUT35), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n497), .A2(KEYINPUT35), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n906), .A2(G116), .A3(new_n216), .A4(new_n907), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n908), .B(KEYINPUT36), .ZN(new_n909));
  NOR3_X1   g0709(.A1(new_n372), .A2(new_n213), .A3(new_n256), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(new_n202), .B2(G68), .ZN(new_n911));
  OR3_X1    g0711(.A1(new_n911), .A2(new_n206), .A3(G13), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n905), .A2(new_n909), .A3(new_n912), .ZN(G367));
  INV_X1    g0713(.A(new_n734), .ZN(new_n914));
  OAI221_X1 g0714(.A(new_n739), .B1(new_n210), .B2(new_n565), .C1(new_n914), .C2(new_n236), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n915), .A2(new_n798), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n776), .A2(new_n435), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT46), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n788), .A2(G97), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n753), .A2(G303), .B1(new_n750), .B2(G283), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n758), .A2(G311), .B1(new_n767), .B2(G294), .ZN(new_n921));
  INV_X1    g0721(.A(G317), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n316), .B1(new_n745), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(G107), .B2(new_n763), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n919), .A2(new_n920), .A3(new_n921), .A4(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n788), .A2(G77), .ZN(new_n926));
  INV_X1    g0726(.A(new_n776), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(G58), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n753), .A2(G150), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n316), .B1(new_n746), .B2(G137), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n926), .A2(new_n928), .A3(new_n929), .A4(new_n930), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n758), .A2(G143), .B1(new_n767), .B2(G159), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n763), .A2(G68), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n932), .B(new_n933), .C1(new_n202), .C2(new_n751), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n918), .A2(new_n925), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n935), .B(KEYINPUT47), .Z(new_n936));
  OAI21_X1  g0736(.A(new_n651), .B1(new_n567), .B2(new_n576), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n683), .A2(new_n937), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n938), .A2(KEYINPUT105), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n937), .B1(new_n620), .B2(new_n624), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n938), .A2(KEYINPUT105), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n916), .B1(new_n742), .B2(new_n936), .C1(new_n943), .C2(new_n730), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n677), .B(KEYINPUT41), .Z(new_n945));
  OAI211_X1 g0745(.A(new_n531), .B(new_n537), .C1(new_n532), .C2(new_n652), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n625), .A2(new_n626), .A3(new_n651), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n674), .B2(new_n673), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT45), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n949), .B(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n674), .ZN(new_n952));
  INV_X1    g0752(.A(new_n673), .ZN(new_n953));
  INV_X1    g0753(.A(new_n948), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT44), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n952), .A2(KEYINPUT44), .A3(new_n953), .A4(new_n954), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n951), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n669), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT108), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n719), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n658), .A2(KEYINPUT108), .A3(G330), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n667), .A2(KEYINPUT107), .A3(new_n670), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n667), .A2(new_n670), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT107), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n967), .A2(new_n672), .A3(new_n968), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n964), .A2(new_n965), .A3(new_n966), .A4(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n966), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n971), .A2(new_n719), .A3(new_n963), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n717), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n951), .A2(new_n959), .A3(new_n669), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n962), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n945), .B1(new_n977), .B2(new_n717), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n722), .A2(G1), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OR3_X1    g0780(.A1(new_n669), .A2(KEYINPUT106), .A3(new_n954), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n943), .A2(KEYINPUT43), .ZN(new_n982));
  OAI21_X1  g0782(.A(KEYINPUT106), .B1(new_n669), .B2(new_n954), .ZN(new_n983));
  AND3_X1   g0783(.A1(new_n981), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n982), .B1(new_n981), .B2(new_n983), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n943), .A2(KEYINPUT43), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n672), .A2(new_n954), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(KEYINPUT42), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n531), .B1(new_n954), .B2(new_n609), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n652), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n988), .A2(KEYINPUT42), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n986), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  OR3_X1    g0794(.A1(new_n984), .A2(new_n985), .A3(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n994), .B1(new_n984), .B2(new_n985), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n944), .B1(new_n980), .B2(new_n997), .ZN(G387));
  OAI21_X1  g0798(.A(new_n316), .B1(new_n745), .B2(new_n760), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n758), .A2(G322), .B1(new_n767), .B2(G311), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n1000), .B1(new_n777), .B2(new_n751), .C1(new_n922), .C2(new_n754), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT48), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n927), .A2(G294), .B1(G283), .B2(new_n763), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT49), .Z(new_n1007));
  AOI211_X1 g0807(.A(new_n999), .B(new_n1007), .C1(G116), .C2(new_n788), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n927), .A2(G77), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n763), .A2(new_n350), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n316), .B1(new_n746), .B2(G150), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n919), .A2(new_n1009), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n758), .A2(G159), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT112), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n753), .A2(G50), .B1(new_n767), .B2(new_n327), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n219), .B2(new_n751), .ZN(new_n1016));
  NOR3_X1   g0816(.A1(new_n1012), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n738), .B1(new_n1008), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n679), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n732), .A2(new_n1019), .B1(new_n343), .B2(new_n676), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n233), .A2(G45), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT110), .Z(new_n1022));
  INV_X1    g0822(.A(KEYINPUT111), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n270), .B1(new_n219), .B2(new_n256), .C1(new_n1019), .C2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(new_n1023), .B2(new_n1019), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n364), .A2(G50), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT50), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n734), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1020), .B1(new_n1022), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n723), .B1(new_n1030), .B2(new_n739), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1018), .B(new_n1031), .C1(new_n668), .C2(new_n730), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n975), .A2(new_n678), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n973), .A2(new_n717), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1033), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n973), .A2(new_n979), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT109), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1036), .A2(new_n1038), .ZN(G393));
  INV_X1    g0839(.A(new_n976), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n669), .B1(new_n951), .B2(new_n959), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n974), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1042), .A2(new_n977), .A3(new_n677), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT113), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n962), .A2(KEYINPUT113), .A3(new_n976), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1045), .A2(new_n1046), .A3(new_n979), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n739), .B1(new_n428), .B2(new_n210), .C1(new_n914), .C2(new_n240), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n798), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G150), .A2(new_n758), .B1(new_n753), .B2(G159), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT51), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n280), .B1(new_n825), .B2(new_n745), .C1(new_n782), .C2(new_n202), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n751), .A2(new_n364), .B1(new_n764), .B2(new_n256), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n813), .B1(new_n219), .B2(new_n776), .ZN(new_n1054));
  NOR4_X1   g0854(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1056), .A2(KEYINPUT114), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G311), .A2(new_n753), .B1(new_n758), .B2(G317), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT52), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n316), .B1(new_n755), .B2(new_n745), .C1(new_n782), .C2(new_n777), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n751), .A2(new_n761), .B1(new_n764), .B2(new_n435), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n343), .A2(new_n774), .B1(new_n776), .B2(new_n772), .ZN(new_n1062));
  OR4_X1    g0862(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1056), .A2(KEYINPUT114), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1057), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1049), .B1(new_n1065), .B2(new_n738), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n948), .B2(new_n730), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1043), .A2(new_n1047), .A3(new_n1067), .ZN(G390));
  NAND2_X1  g0868(.A1(new_n865), .A2(new_n868), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n804), .A2(new_n880), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n889), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n872), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1069), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n863), .A2(new_n872), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n652), .B(new_n800), .C1(new_n688), .C2(new_n691), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n879), .B1(new_n1075), .B2(new_n880), .ZN(new_n1076));
  OR2_X1    g0876(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n888), .A2(G330), .A3(new_n803), .A4(new_n889), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT115), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OR2_X1    g0880(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1073), .A2(new_n1077), .A3(new_n1080), .A4(new_n1081), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n865), .A2(new_n868), .B1(new_n1071), .B2(new_n872), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1079), .B(new_n1078), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n425), .A2(new_n715), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n885), .A2(new_n644), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT116), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1078), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n889), .B1(new_n715), .B2(new_n803), .ZN(new_n1091));
  OR2_X1    g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1089), .B(new_n889), .C1(new_n715), .C2(new_n803), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1092), .A2(new_n1070), .A3(new_n1094), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n1075), .A2(new_n880), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n805), .A2(new_n715), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1096), .B(new_n1078), .C1(new_n1097), .C2(new_n889), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1088), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1086), .A2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1070), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1098), .B1(new_n1101), .B2(new_n1093), .ZN(new_n1102));
  AND3_X1   g0902(.A1(new_n885), .A2(new_n644), .A3(new_n1087), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1104), .A2(new_n1085), .A3(new_n1082), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1100), .A2(new_n677), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n316), .B1(new_n746), .B2(G125), .ZN(new_n1107));
  INV_X1    g0907(.A(G128), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n1107), .B1(new_n774), .B2(new_n202), .C1(new_n1108), .C2(new_n759), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(KEYINPUT54), .B(G143), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n754), .A2(new_n829), .B1(new_n751), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(G137), .ZN(new_n1112));
  INV_X1    g0912(.A(G159), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n782), .A2(new_n1112), .B1(new_n764), .B2(new_n1113), .ZN(new_n1114));
  NOR3_X1   g0914(.A1(new_n1109), .A2(new_n1111), .A3(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n776), .A2(new_n826), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT53), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n316), .B1(new_n745), .B2(new_n761), .C1(new_n764), .C2(new_n256), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n1118), .B(new_n787), .C1(G68), .C2(new_n788), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n759), .A2(new_n772), .B1(new_n751), .B2(new_n428), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n754), .A2(new_n435), .B1(new_n782), .B2(new_n343), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n1115), .A2(new_n1117), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n798), .B1(new_n327), .B2(new_n810), .C1(new_n1123), .C2(new_n742), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(new_n1069), .B2(new_n727), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(new_n1086), .B2(new_n979), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1106), .A2(new_n1126), .ZN(G378));
  NAND2_X1  g0927(.A1(new_n897), .A2(G330), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n633), .A2(new_n361), .A3(new_n634), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n331), .A2(new_n649), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1130), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  OR2_X1    g0936(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1137), .A2(new_n1133), .A3(new_n1129), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n874), .A2(new_n1139), .A3(new_n882), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1139), .B1(new_n874), .B2(new_n882), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1128), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1139), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n883), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n874), .A2(new_n1139), .A3(new_n882), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n695), .B1(new_n894), .B2(new_n896), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1142), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1104), .B1(new_n1085), .B2(new_n1082), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1088), .B(KEYINPUT119), .ZN(new_n1150));
  OAI211_X1 g0950(.A(KEYINPUT57), .B(new_n1148), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(KEYINPUT120), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1150), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1100), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT120), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1154), .A2(new_n1155), .A3(KEYINPUT57), .A4(new_n1148), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT57), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1150), .B1(new_n1086), .B2(new_n1099), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n1142), .A2(new_n1147), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1157), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1152), .A2(new_n677), .A3(new_n1156), .A4(new_n1160), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(G33), .A2(G41), .ZN(new_n1162));
  AOI211_X1 g0962(.A(G50), .B(new_n1162), .C1(new_n316), .C2(new_n269), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n753), .A2(G107), .B1(new_n767), .B2(G97), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1164), .B1(new_n435), .B2(new_n759), .C1(new_n565), .C2(new_n751), .ZN(new_n1165));
  AOI211_X1 g0965(.A(G41), .B(new_n280), .C1(new_n746), .C2(G283), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1009), .A2(new_n933), .A3(new_n1166), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n774), .A2(new_n371), .ZN(new_n1168));
  NOR3_X1   g0968(.A1(new_n1165), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT117), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT58), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1163), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n1171), .B2(new_n1170), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n753), .A2(G128), .B1(new_n767), .B2(G132), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n776), .B2(new_n1110), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n758), .A2(G125), .B1(G150), .B2(new_n763), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n1112), .B2(new_n751), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT59), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT118), .ZN(new_n1180));
  AND2_X1   g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n746), .A2(G124), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1162), .B(new_n1183), .C1(new_n774), .C2(new_n1113), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n1181), .A2(new_n1182), .A3(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n738), .B1(new_n1173), .B2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n723), .B1(new_n202), .B2(new_n809), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(new_n1143), .B2(new_n727), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(new_n1148), .B2(new_n979), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1161), .A2(new_n1190), .ZN(G375));
  INV_X1    g0991(.A(new_n1102), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(new_n1088), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n945), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1193), .A2(new_n1194), .A3(new_n1104), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n879), .A2(new_n727), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n798), .B1(G68), .B2(new_n810), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n280), .B1(new_n746), .B2(G303), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n926), .A2(new_n1010), .A3(new_n1198), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n758), .A2(G294), .B1(new_n750), .B2(G107), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1200), .B1(new_n435), .B2(new_n782), .C1(new_n772), .C2(new_n754), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1199), .B(new_n1201), .C1(G97), .C2(new_n927), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  OR2_X1    g1003(.A1(new_n1203), .A2(KEYINPUT121), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n280), .B1(new_n745), .B2(new_n1108), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1205), .B(new_n1168), .C1(G132), .C2(new_n758), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n754), .A2(new_n1112), .B1(new_n202), .B2(new_n764), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n1110), .A2(new_n782), .B1(new_n751), .B2(new_n826), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1206), .B(new_n1209), .C1(new_n1113), .C2(new_n776), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1203), .A2(KEYINPUT121), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1204), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1197), .B1(new_n1212), .B2(new_n738), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1102), .A2(new_n979), .B1(new_n1196), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1195), .A2(new_n1214), .ZN(G381));
  XNOR2_X1  g1015(.A(G375), .B(KEYINPUT122), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1036), .A2(new_n796), .A3(new_n1038), .ZN(new_n1217));
  OR4_X1    g1017(.A1(G384), .A2(G390), .A3(new_n1217), .A4(G381), .ZN(new_n1218));
  OR4_X1    g1018(.A1(G387), .A2(new_n1216), .A3(G378), .A4(new_n1218), .ZN(G407));
  INV_X1    g1019(.A(G378), .ZN(new_n1220));
  INV_X1    g1020(.A(G213), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1221), .A2(G343), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1220), .A2(new_n1222), .ZN(new_n1223));
  OAI211_X1 g1023(.A(G407), .B(G213), .C1(new_n1216), .C2(new_n1223), .ZN(G409));
  INV_X1    g1024(.A(KEYINPUT124), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1161), .A2(G378), .A3(new_n1190), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1154), .A2(new_n1194), .A3(new_n1148), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(KEYINPUT123), .B2(new_n1190), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n1190), .A2(KEYINPUT123), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1220), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1226), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1222), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1095), .A2(KEYINPUT60), .A3(new_n1088), .A4(new_n1098), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n677), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1104), .A2(KEYINPUT60), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1234), .B1(new_n1193), .B2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1214), .ZN(new_n1237));
  OR3_X1    g1037(.A1(new_n1236), .A2(new_n835), .A3(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n835), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1231), .A2(KEYINPUT63), .A3(new_n1232), .A4(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT61), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1222), .B1(new_n1226), .B2(new_n1230), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1222), .A2(G2897), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1240), .B(new_n1246), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1242), .B(new_n1243), .C1(new_n1244), .C2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(G393), .A2(G396), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n1217), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n995), .B(new_n996), .C1(new_n978), .C2(new_n979), .ZN(new_n1251));
  AND3_X1   g1051(.A1(new_n1251), .A2(new_n944), .A3(G390), .ZN(new_n1252));
  AOI21_X1  g1052(.A(G390), .B1(new_n1251), .B2(new_n944), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1250), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(G390), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(G387), .A2(new_n1255), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1249), .A2(new_n1217), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1251), .A2(new_n944), .A3(G390), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1256), .A2(new_n1257), .A3(new_n1258), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1254), .A2(new_n1259), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n1222), .B(new_n1240), .C1(new_n1226), .C2(new_n1230), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1260), .B1(new_n1261), .B2(KEYINPUT63), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1225), .B1(new_n1248), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1254), .A2(new_n1259), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1244), .A2(new_n1241), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT63), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1264), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1244), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(new_n1240), .B(new_n1245), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT61), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1267), .A2(new_n1270), .A3(KEYINPUT124), .A4(new_n1242), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1263), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1270), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1274), .B1(new_n1244), .B2(new_n1241), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT126), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(new_n1275), .A2(new_n1276), .B1(KEYINPUT62), .B2(new_n1261), .ZN(new_n1277));
  OAI21_X1  g1077(.A(KEYINPUT126), .B1(new_n1261), .B2(new_n1274), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1273), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1264), .B(KEYINPUT127), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1272), .B1(new_n1279), .B2(new_n1280), .ZN(G405));
  NAND2_X1  g1081(.A1(G375), .A2(new_n1220), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1226), .ZN(new_n1283));
  XNOR2_X1  g1083(.A(new_n1283), .B(new_n1241), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(new_n1284), .B(new_n1264), .ZN(G402));
endmodule


