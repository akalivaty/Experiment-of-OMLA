//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 0 1 1 0 0 1 0 1 0 1 0 0 1 0 0 1 0 1 0 0 1 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 0 0 1 1 0 0 1 1 0 1 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n623,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT64), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT66), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n463), .A2(new_n464), .A3(G101), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n466), .A2(G101), .A3(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT67), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  OAI211_X1 g046(.A(G137), .B(new_n466), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g048(.A(G125), .B1(new_n470), .B2(new_n471), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n466), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n473), .A2(new_n476), .ZN(G160));
  NOR2_X1   g052(.A1(new_n470), .A2(new_n471), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(new_n466), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n480), .B(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n478), .A2(G2105), .ZN(new_n483));
  MUX2_X1   g058(.A(G100), .B(G112), .S(G2105), .Z(new_n484));
  AOI22_X1  g059(.A1(new_n483), .A2(G136), .B1(G2104), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT69), .ZN(G162));
  INV_X1    g062(.A(G126), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT3), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(new_n462), .ZN(new_n490));
  NAND2_X1  g065(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n488), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AND2_X1   g067(.A1(G114), .A2(G2104), .ZN(new_n493));
  OAI21_X1  g068(.A(G2105), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(KEYINPUT4), .A2(G138), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n495), .B1(new_n490), .B2(new_n491), .ZN(new_n496));
  NAND2_X1  g071(.A1(G102), .A2(G2104), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n466), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  OAI211_X1 g074(.A(G138), .B(new_n466), .C1(new_n470), .C2(new_n471), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n494), .A2(new_n499), .A3(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT70), .B1(new_n507), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(new_n505), .A3(KEYINPUT5), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n506), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT6), .B(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  INV_X1    g092(.A(G50), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n515), .A2(G543), .ZN(new_n519));
  OAI22_X1  g094(.A1(new_n516), .A2(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n514), .A2(new_n520), .ZN(G166));
  INV_X1    g096(.A(new_n519), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G51), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  AND3_X1   g101(.A1(new_n523), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n516), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G89), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n527), .A2(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  AOI22_X1  g106(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n513), .ZN(new_n533));
  XNOR2_X1  g108(.A(KEYINPUT71), .B(G90), .ZN(new_n534));
  INV_X1    g109(.A(G52), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n516), .A2(new_n534), .B1(new_n535), .B2(new_n519), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n533), .A2(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  INV_X1    g113(.A(G81), .ZN(new_n539));
  INV_X1    g114(.A(G43), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n516), .A2(new_n539), .B1(new_n540), .B2(new_n519), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n541), .A2(KEYINPUT73), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(KEYINPUT73), .ZN(new_n543));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n508), .A2(new_n510), .ZN(new_n545));
  INV_X1    g120(.A(new_n506), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n544), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(KEYINPUT72), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n513), .B1(new_n549), .B2(KEYINPUT72), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n542), .A2(new_n543), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  AND3_X1   g128(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G36), .ZN(G176));
  XOR2_X1   g130(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n556));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n556), .B(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT75), .ZN(G188));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G65), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n547), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G651), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n528), .A2(G91), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n515), .A2(G53), .A3(G543), .ZN(new_n566));
  NAND2_X1  g141(.A1(KEYINPUT76), .A2(KEYINPUT9), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n515), .A2(G53), .A3(G543), .A4(new_n567), .ZN(new_n570));
  AND3_X1   g145(.A1(new_n569), .A2(KEYINPUT77), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g146(.A(KEYINPUT77), .B1(new_n569), .B2(new_n570), .ZN(new_n572));
  OAI211_X1 g147(.A(new_n564), .B(new_n565), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(KEYINPUT78), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n511), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G91), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n575), .A2(new_n513), .B1(new_n576), .B2(new_n516), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n578), .B(new_n579), .C1(new_n572), .C2(new_n571), .ZN(new_n580));
  AND2_X1   g155(.A1(new_n574), .A2(new_n580), .ZN(G299));
  INV_X1    g156(.A(G166), .ZN(G303));
  NAND2_X1  g157(.A1(new_n522), .A2(G49), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n511), .A2(G87), .A3(new_n515), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(G288));
  NAND3_X1  g161(.A1(new_n515), .A2(G48), .A3(G543), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n545), .A2(G61), .A3(new_n546), .ZN(new_n589));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n588), .B1(new_n591), .B2(G651), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n545), .A2(G86), .A3(new_n546), .A4(new_n515), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(KEYINPUT79), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT79), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n511), .A2(new_n595), .A3(G86), .A4(new_n515), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n592), .A2(new_n597), .ZN(G305));
  AOI22_X1  g173(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n599), .A2(new_n513), .ZN(new_n600));
  INV_X1    g175(.A(G85), .ZN(new_n601));
  INV_X1    g176(.A(G47), .ZN(new_n602));
  OAI22_X1  g177(.A1(new_n516), .A2(new_n601), .B1(new_n602), .B2(new_n519), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT80), .ZN(new_n604));
  OR3_X1    g179(.A1(new_n600), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n600), .B2(new_n603), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(G290));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  NOR2_X1   g183(.A1(G301), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n511), .A2(G92), .A3(new_n515), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(G79), .A2(G543), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT81), .ZN(new_n614));
  INV_X1    g189(.A(G66), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n547), .B2(new_n615), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n616), .A2(G651), .B1(G54), .B2(new_n522), .ZN(new_n617));
  AND2_X1   g192(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n609), .B1(new_n608), .B2(new_n618), .ZN(G284));
  AOI21_X1  g194(.A(new_n609), .B1(new_n608), .B2(new_n618), .ZN(G321));
  NAND2_X1  g195(.A1(G286), .A2(G868), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT82), .Z(new_n622));
  NAND2_X1  g197(.A1(G299), .A2(new_n608), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(G297));
  XNOR2_X1  g199(.A(G297), .B(KEYINPUT83), .ZN(G280));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n618), .B1(new_n626), .B2(G860), .ZN(G148));
  INV_X1    g202(.A(new_n552), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n628), .A2(G868), .ZN(new_n629));
  INV_X1    g204(.A(new_n618), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n630), .A2(G559), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n629), .B1(G868), .B2(new_n631), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g208(.A1(new_n483), .A2(G2104), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT12), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  INV_X1    g211(.A(G2100), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n483), .A2(G135), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n479), .A2(G123), .ZN(new_n641));
  MUX2_X1   g216(.A(G99), .B(G111), .S(G2105), .Z(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(G2104), .ZN(new_n643));
  AND3_X1   g218(.A1(new_n640), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2096), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n638), .A2(new_n639), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT84), .Z(G156));
  INV_X1    g222(.A(KEYINPUT14), .ZN(new_n648));
  XOR2_X1   g223(.A(KEYINPUT15), .B(G2435), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2438), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2427), .ZN(new_n651));
  INV_X1    g226(.A(G2430), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n648), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(new_n652), .B2(new_n651), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2451), .B(G2454), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT16), .ZN(new_n656));
  XOR2_X1   g231(.A(G2443), .B(G2446), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1341), .B(G1348), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT85), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n658), .B(new_n660), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n654), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n654), .A2(new_n661), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n662), .A2(G14), .A3(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(G401));
  XNOR2_X1  g240(.A(G2072), .B(G2078), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT17), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2084), .B(G2090), .ZN(new_n669));
  NOR3_X1   g244(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT88), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT87), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n669), .B1(new_n666), .B2(new_n668), .ZN(new_n673));
  AOI22_X1  g248(.A1(new_n667), .A2(new_n668), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n674), .B1(new_n672), .B2(new_n673), .ZN(new_n675));
  INV_X1    g250(.A(new_n669), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n676), .A2(new_n666), .A3(new_n668), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT86), .B(KEYINPUT18), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n671), .A2(new_n675), .A3(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(G2096), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n682), .A2(G2100), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(G2100), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(G227));
  XNOR2_X1  g261(.A(G1961), .B(G1966), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT89), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G1956), .B(G2474), .Z(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1971), .B(G1976), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT19), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT90), .B(KEYINPUT20), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n689), .A2(new_n690), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n697), .A2(new_n693), .A3(new_n691), .ZN(new_n698));
  OAI211_X1 g273(.A(new_n696), .B(new_n698), .C1(new_n693), .C2(new_n697), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(G1991), .B(G1996), .Z(new_n702));
  XNOR2_X1  g277(.A(G1981), .B(G1986), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n702), .B(new_n703), .Z(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n701), .B(new_n705), .ZN(G229));
  MUX2_X1   g281(.A(G6), .B(G305), .S(G16), .Z(new_n707));
  XOR2_X1   g282(.A(KEYINPUT32), .B(G1981), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G23), .ZN(new_n711));
  INV_X1    g286(.A(G288), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(new_n712), .B2(new_n710), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT33), .B(G1976), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(G16), .A2(G22), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G166), .B2(G16), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(G1971), .Z(new_n718));
  AND3_X1   g293(.A1(new_n709), .A2(new_n715), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT92), .B(KEYINPUT34), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  MUX2_X1   g297(.A(G95), .B(G107), .S(G2105), .Z(new_n723));
  AOI22_X1  g298(.A1(new_n479), .A2(G119), .B1(G2104), .B2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G131), .ZN(new_n725));
  INV_X1    g300(.A(new_n483), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  MUX2_X1   g302(.A(G25), .B(new_n727), .S(G29), .Z(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT35), .B(G1991), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT91), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n728), .B(new_n730), .Z(new_n731));
  INV_X1    g306(.A(G290), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G16), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G16), .B2(G24), .ZN(new_n734));
  INV_X1    g309(.A(G1986), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n731), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n735), .B2(new_n734), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n721), .A2(new_n722), .A3(new_n737), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT36), .Z(new_n739));
  MUX2_X1   g314(.A(G104), .B(G116), .S(G2105), .Z(new_n740));
  AOI22_X1  g315(.A1(new_n479), .A2(G128), .B1(G2104), .B2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(G140), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n741), .B1(new_n742), .B2(new_n726), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G29), .ZN(new_n744));
  INV_X1    g319(.A(G29), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(G26), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT28), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(G2067), .Z(new_n749));
  NOR2_X1   g324(.A1(G168), .A2(new_n710), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n710), .B2(G21), .ZN(new_n751));
  INV_X1    g326(.A(G1966), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n749), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n745), .A2(G32), .ZN(new_n754));
  AOI22_X1  g329(.A1(G129), .A2(new_n479), .B1(new_n483), .B2(G141), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n463), .A2(G105), .ZN(new_n756));
  NAND3_X1  g331(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT26), .Z(new_n758));
  NAND3_X1  g333(.A1(new_n755), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n754), .B1(new_n760), .B2(new_n745), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT27), .B(G1996), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  AND2_X1   g338(.A1(KEYINPUT24), .A2(G34), .ZN(new_n764));
  NOR2_X1   g339(.A1(KEYINPUT24), .A2(G34), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n745), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(G160), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n766), .B1(new_n767), .B2(new_n745), .ZN(new_n768));
  INV_X1    g343(.A(G2084), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n644), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n771), .A2(new_n745), .ZN(new_n772));
  OR2_X1    g347(.A1(KEYINPUT30), .A2(G28), .ZN(new_n773));
  NAND2_X1  g348(.A1(KEYINPUT30), .A2(G28), .ZN(new_n774));
  AOI21_X1  g349(.A(G29), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT31), .B(G11), .Z(new_n776));
  NOR4_X1   g351(.A1(new_n770), .A2(new_n772), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n710), .A2(G5), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G171), .B2(new_n710), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n763), .B(new_n777), .C1(G1961), .C2(new_n779), .ZN(new_n780));
  AOI211_X1 g355(.A(new_n753), .B(new_n780), .C1(new_n752), .C2(new_n751), .ZN(new_n781));
  NOR2_X1   g356(.A1(G29), .A2(G33), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT94), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n490), .A2(new_n491), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n784), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n785), .A2(new_n466), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n786), .A2(KEYINPUT95), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(KEYINPUT95), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n463), .A2(G103), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT25), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n463), .A2(KEYINPUT25), .A3(G103), .ZN(new_n792));
  AOI22_X1  g367(.A1(G139), .A2(new_n483), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n787), .A2(new_n788), .A3(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n783), .B1(new_n794), .B2(new_n745), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G2072), .ZN(new_n796));
  NOR2_X1   g371(.A1(G4), .A2(G16), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n618), .B2(G16), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT93), .B(G1348), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(G27), .A2(G29), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G164), .B2(G29), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G2078), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n768), .A2(new_n769), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT96), .Z(new_n805));
  AOI211_X1 g380(.A(new_n803), .B(new_n805), .C1(G1961), .C2(new_n779), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n781), .A2(new_n796), .A3(new_n800), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(G299), .A2(G16), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n710), .A2(G20), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT23), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(G1956), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n807), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(G16), .A2(G19), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(new_n552), .B2(G16), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(G1341), .Z(new_n816));
  NAND2_X1  g391(.A1(new_n745), .A2(G35), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G162), .B2(new_n745), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT29), .ZN(new_n819));
  INV_X1    g394(.A(G2090), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n813), .A2(new_n816), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n739), .A2(new_n822), .ZN(G311));
  INV_X1    g398(.A(G311), .ZN(G150));
  NAND2_X1  g399(.A1(G80), .A2(G543), .ZN(new_n825));
  INV_X1    g400(.A(G67), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n547), .B2(new_n826), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n827), .A2(KEYINPUT98), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n513), .B1(new_n827), .B2(KEYINPUT98), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT99), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n828), .A2(KEYINPUT99), .A3(new_n829), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n528), .A2(G93), .B1(G55), .B2(new_n522), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(G860), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT37), .Z(new_n838));
  AND3_X1   g413(.A1(new_n834), .A2(new_n552), .A3(new_n835), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n552), .B1(new_n834), .B2(new_n835), .ZN(new_n840));
  NOR4_X1   g415(.A1(new_n839), .A2(new_n840), .A3(new_n626), .A4(new_n630), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n836), .A2(new_n628), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n834), .A2(new_n552), .A3(new_n835), .ZN(new_n843));
  AOI22_X1  g418(.A1(new_n842), .A2(new_n843), .B1(G559), .B2(new_n618), .ZN(new_n844));
  XOR2_X1   g419(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n845));
  OR3_X1    g420(.A1(new_n841), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n845), .B1(new_n841), .B2(new_n844), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT39), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(G860), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n848), .B1(new_n846), .B2(new_n847), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n838), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT100), .ZN(G145));
  XNOR2_X1  g429(.A(new_n743), .B(G164), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n794), .A2(KEYINPUT101), .A3(new_n759), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n759), .B1(new_n794), .B2(KEYINPUT101), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n855), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n858), .ZN(new_n860));
  INV_X1    g435(.A(new_n855), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n860), .A2(new_n856), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n635), .B(new_n727), .ZN(new_n864));
  MUX2_X1   g439(.A(G106), .B(G118), .S(G2105), .Z(new_n865));
  AOI22_X1  g440(.A1(new_n479), .A2(G130), .B1(G2104), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(G142), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n866), .B1(new_n867), .B2(new_n726), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n864), .B(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n863), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n869), .A2(new_n862), .A3(new_n859), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(G162), .A2(new_n767), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT69), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n486), .B(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(G160), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n771), .B1(new_n874), .B2(new_n877), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n874), .A2(new_n877), .A3(new_n771), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n873), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n878), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT102), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n869), .A2(new_n882), .A3(new_n862), .A4(new_n859), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n872), .A2(KEYINPUT102), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n881), .A2(new_n883), .A3(new_n884), .A4(new_n871), .ZN(new_n885));
  INV_X1    g460(.A(G37), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n880), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT103), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT103), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n880), .A2(new_n885), .A3(new_n889), .A4(new_n886), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g467(.A1(new_n836), .A2(new_n608), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n618), .B1(new_n574), .B2(new_n580), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n894), .A2(KEYINPUT104), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(KEYINPUT104), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n574), .A2(new_n580), .A3(new_n618), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n631), .B1(new_n839), .B2(new_n840), .ZN(new_n899));
  INV_X1    g474(.A(new_n631), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n842), .A2(new_n900), .A3(new_n843), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n898), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT105), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n898), .A2(new_n899), .A3(new_n901), .A4(KEYINPUT105), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n899), .A2(new_n901), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT41), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n895), .A2(new_n908), .A3(new_n896), .A4(new_n897), .ZN(new_n909));
  INV_X1    g484(.A(new_n896), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n897), .B1(new_n894), .B2(KEYINPUT104), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT41), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n907), .A2(new_n909), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT106), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n907), .A2(new_n912), .A3(new_n909), .A4(KEYINPUT106), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n732), .A2(new_n712), .ZN(new_n917));
  NAND2_X1  g492(.A1(G290), .A2(G288), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(G305), .B(G166), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n917), .A2(new_n918), .A3(new_n920), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT42), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT42), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n922), .A2(new_n926), .A3(new_n923), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n906), .A2(new_n915), .A3(new_n916), .A4(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT107), .ZN(new_n930));
  AOI22_X1  g505(.A1(new_n904), .A2(new_n905), .B1(new_n913), .B2(new_n914), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT107), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n931), .A2(new_n932), .A3(new_n916), .A4(new_n928), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n906), .A2(new_n916), .A3(new_n915), .ZN(new_n934));
  INV_X1    g509(.A(new_n928), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n930), .A2(new_n933), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n893), .B1(new_n937), .B2(new_n608), .ZN(G295));
  OAI21_X1  g513(.A(new_n893), .B1(new_n937), .B2(new_n608), .ZN(G331));
  XOR2_X1   g514(.A(G301), .B(G286), .Z(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n941), .B1(new_n839), .B2(new_n840), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n842), .A2(new_n940), .A3(new_n843), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n898), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT109), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT109), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n898), .A2(new_n942), .A3(new_n943), .A4(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n942), .A2(new_n943), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n948), .A2(new_n912), .A3(new_n909), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n945), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n950), .A2(new_n922), .A3(new_n923), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT43), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n945), .A2(new_n949), .A3(new_n947), .A4(new_n924), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n951), .A2(new_n952), .A3(new_n886), .A4(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n886), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n924), .B1(new_n949), .B2(new_n944), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT43), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n954), .A2(new_n957), .A3(KEYINPUT44), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n951), .A2(KEYINPUT43), .A3(new_n886), .A4(new_n953), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n952), .B1(new_n955), .B2(new_n956), .ZN(new_n960));
  XOR2_X1   g535(.A(KEYINPUT108), .B(KEYINPUT44), .Z(new_n961));
  NAND3_X1  g536(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n958), .A2(new_n962), .ZN(G397));
  INV_X1    g538(.A(G1384), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n503), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT45), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n476), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n968), .A2(G40), .A3(new_n469), .A4(new_n472), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G1996), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n972), .B(KEYINPUT111), .ZN(new_n973));
  OR2_X1    g548(.A1(new_n973), .A2(KEYINPUT46), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(KEYINPUT46), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n743), .B(G2067), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n970), .B1(new_n976), .B2(new_n759), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n974), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n978), .B(KEYINPUT47), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n970), .A2(G1996), .A3(new_n759), .ZN(new_n980));
  OR2_X1    g555(.A1(new_n980), .A2(KEYINPUT112), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(KEYINPUT112), .ZN(new_n982));
  AOI22_X1  g557(.A1(new_n981), .A2(new_n982), .B1(new_n970), .B2(new_n976), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n973), .A2(new_n760), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n985), .A2(new_n730), .A3(new_n727), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n743), .A2(G2067), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n970), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n727), .B(new_n730), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n985), .B1(new_n970), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n732), .A2(new_n735), .ZN(new_n991));
  INV_X1    g566(.A(new_n970), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  XOR2_X1   g568(.A(new_n993), .B(KEYINPUT48), .Z(new_n994));
  NAND2_X1  g569(.A1(new_n990), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n979), .A2(new_n988), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT126), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT126), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n979), .A2(new_n988), .A3(new_n998), .A4(new_n995), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G1981), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n592), .A2(new_n1001), .A3(new_n597), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n590), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1004), .B1(new_n511), .B2(G61), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n587), .B(new_n593), .C1(new_n1005), .C2(new_n513), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(G1981), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT115), .B1(new_n1002), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT49), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  AOI211_X1 g585(.A(KEYINPUT115), .B(KEYINPUT49), .C1(new_n1002), .C2(new_n1007), .ZN(new_n1011));
  INV_X1    g586(.A(G8), .ZN(new_n1012));
  INV_X1    g587(.A(new_n495), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1013), .B1(new_n470), .B2(new_n471), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n497), .ZN(new_n1015));
  AOI22_X1  g590(.A1(new_n1015), .A2(new_n466), .B1(new_n501), .B2(new_n500), .ZN(new_n1016));
  AOI21_X1  g591(.A(G1384), .B1(new_n1016), .B2(new_n494), .ZN(new_n1017));
  INV_X1    g592(.A(G40), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n473), .A2(new_n476), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1012), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  OR3_X1    g596(.A1(new_n1010), .A2(new_n1011), .A3(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(G288), .A2(G1976), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1003), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n583), .A2(new_n584), .A3(G1976), .A4(new_n585), .ZN(new_n1026));
  INV_X1    g601(.A(G1976), .ZN(new_n1027));
  NAND2_X1  g602(.A1(G288), .A2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1020), .A2(new_n1025), .A3(new_n1026), .A4(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1025), .B1(new_n1020), .B2(new_n1026), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1029), .B1(new_n1030), .B2(KEYINPUT114), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1019), .A2(new_n964), .A3(new_n503), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n1032), .A2(G8), .A3(new_n1026), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1033), .A2(new_n1034), .A3(new_n1025), .A4(new_n1028), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1022), .A2(new_n1031), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1037), .B1(G166), .B2(new_n1012), .ZN(new_n1038));
  OAI211_X1 g613(.A(KEYINPUT55), .B(G8), .C1(new_n514), .C2(new_n520), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n503), .A2(KEYINPUT50), .A3(new_n964), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT50), .B1(new_n503), .B2(new_n964), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n820), .B(new_n1019), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g619(.A(KEYINPUT113), .B(G1971), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n969), .B1(new_n965), .B2(new_n966), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n964), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1045), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  OAI211_X1 g623(.A(G8), .B(new_n1040), .C1(new_n1044), .C2(new_n1048), .ZN(new_n1049));
  OAI22_X1  g624(.A1(new_n1024), .A2(new_n1021), .B1(new_n1036), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(KEYINPUT116), .ZN(new_n1051));
  OAI21_X1  g626(.A(G8), .B1(new_n1044), .B2(new_n1048), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1040), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1031), .A2(new_n1035), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n1010), .A2(new_n1011), .A3(new_n1021), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1052), .A2(KEYINPUT116), .A3(new_n1053), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n967), .A2(new_n1019), .A3(new_n1047), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(new_n752), .ZN(new_n1061));
  XOR2_X1   g636(.A(KEYINPUT117), .B(G2084), .Z(new_n1062));
  OAI211_X1 g637(.A(new_n1019), .B(new_n1062), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(G8), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1065), .A2(G286), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1055), .A2(new_n1058), .A3(new_n1059), .A4(new_n1066), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT118), .B(KEYINPUT63), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AND2_X1   g644(.A1(new_n1053), .A2(KEYINPUT119), .ZN(new_n1070));
  OR2_X1    g645(.A1(new_n1070), .A2(new_n1052), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT63), .ZN(new_n1072));
  NOR3_X1   g647(.A1(new_n1065), .A2(new_n1072), .A3(G286), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1070), .A2(new_n1052), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1071), .A2(new_n1073), .A3(new_n1058), .A4(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1050), .B1(new_n1069), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G2078), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n967), .A2(new_n1077), .A3(new_n1019), .A4(new_n1047), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1019), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1081));
  INV_X1    g656(.A(G1961), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1046), .A2(KEYINPUT53), .A3(new_n1077), .A4(new_n1047), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1080), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(G171), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1055), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1088));
  AOI211_X1 g663(.A(new_n1012), .B(G168), .C1(new_n1061), .C2(new_n1063), .ZN(new_n1089));
  NAND2_X1  g664(.A1(G286), .A2(G8), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1091), .B1(new_n1064), .B2(G8), .ZN(new_n1092));
  AOI21_X1  g667(.A(KEYINPUT51), .B1(new_n1090), .B2(KEYINPUT123), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1089), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  OAI211_X1 g670(.A(G8), .B(new_n1093), .C1(new_n1064), .C2(G286), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1095), .A2(KEYINPUT62), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT62), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1087), .B(new_n1088), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1032), .A2(G2067), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1100), .B1(new_n1081), .B2(new_n799), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1101), .A2(new_n630), .ZN(new_n1102));
  INV_X1    g677(.A(G1956), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1081), .A2(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(KEYINPUT56), .B(G2072), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1046), .A2(new_n1047), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT121), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1104), .A2(new_n1106), .A3(KEYINPUT121), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT120), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n577), .A2(new_n1112), .ZN(new_n1113));
  OAI221_X1 g688(.A(KEYINPUT120), .B1(new_n516), .B2(new_n576), .C1(new_n575), .C2(new_n513), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(KEYINPUT57), .B1(new_n569), .B2(new_n570), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n1115), .A2(new_n1116), .B1(new_n573), .B2(KEYINPUT57), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1102), .B1(new_n1111), .B2(new_n1118), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1117), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT61), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1117), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1122), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1124));
  AOI211_X1 g699(.A(new_n618), .B(new_n1100), .C1(new_n799), .C2(new_n1081), .ZN(new_n1125));
  OAI21_X1  g700(.A(KEYINPUT60), .B1(new_n1102), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT60), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1101), .A2(new_n1127), .A3(new_n618), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1124), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(KEYINPUT61), .B1(new_n1107), .B2(new_n1118), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1130), .B1(new_n1111), .B2(new_n1118), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(KEYINPUT58), .B(G1341), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1133), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1046), .A2(new_n971), .A3(new_n1047), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1134), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  OR3_X1    g714(.A1(new_n1139), .A2(KEYINPUT59), .A3(new_n628), .ZN(new_n1140));
  OAI21_X1  g715(.A(KEYINPUT59), .B1(new_n1139), .B2(new_n628), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1121), .B1(new_n1132), .B2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1080), .A2(new_n1083), .A3(G301), .A4(new_n1084), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1086), .A2(KEYINPUT54), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(KEYINPUT124), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT124), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1086), .A2(new_n1147), .A3(KEYINPUT54), .A4(new_n1144), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1086), .A2(new_n1144), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT54), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1149), .A2(new_n1088), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1076), .B(new_n1099), .C1(new_n1143), .C2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(G290), .A2(G1986), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n992), .B1(new_n991), .B2(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1157), .B(KEYINPUT110), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n990), .A2(new_n1158), .ZN(new_n1159));
  AND3_X1   g734(.A1(new_n1155), .A2(KEYINPUT125), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(KEYINPUT125), .B1(new_n1155), .B2(new_n1159), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1000), .B1(new_n1160), .B2(new_n1161), .ZN(G329));
  assign    G231 = 1'b0;
  NAND4_X1  g737(.A1(new_n683), .A2(G319), .A3(new_n664), .A4(new_n684), .ZN(new_n1164));
  OAI21_X1  g738(.A(KEYINPUT127), .B1(G229), .B2(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g739(.A(new_n701), .B(new_n704), .ZN(new_n1166));
  INV_X1    g740(.A(KEYINPUT127), .ZN(new_n1167));
  AND2_X1   g741(.A1(new_n664), .A2(G319), .ZN(new_n1168));
  NAND4_X1  g742(.A1(new_n1166), .A2(new_n685), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  NAND2_X1  g743(.A1(new_n1165), .A2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g744(.A(new_n1170), .B1(new_n888), .B2(new_n890), .ZN(new_n1171));
  AND3_X1   g745(.A1(new_n1171), .A2(new_n960), .A3(new_n959), .ZN(G308));
  NAND3_X1  g746(.A1(new_n1171), .A2(new_n960), .A3(new_n959), .ZN(G225));
endmodule


