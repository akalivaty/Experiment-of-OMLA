//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 0 1 0 1 1 1 1 1 0 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 1 1 1 1 0 1 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n818, new_n819, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n955, new_n956, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1016, new_n1017, new_n1018, new_n1019;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(G141gat), .ZN(new_n204));
  INV_X1    g003(.A(G148gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT2), .ZN(new_n207));
  NAND2_X1  g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G162gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G155gat), .ZN(new_n211));
  INV_X1    g010(.A(G155gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G162gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n209), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(KEYINPUT77), .B(G162gat), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n207), .B1(new_n216), .B2(G155gat), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n206), .A2(new_n211), .A3(new_n213), .A4(new_n208), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n215), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AND2_X1   g018(.A1(KEYINPUT68), .A2(G120gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(KEYINPUT68), .A2(G120gat), .ZN(new_n221));
  OAI21_X1  g020(.A(G113gat), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G113gat), .ZN(new_n223));
  INV_X1    g022(.A(G120gat), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT1), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G127gat), .B(G134gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n222), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G134gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G127gat), .ZN(new_n229));
  INV_X1    g028(.A(G127gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G134gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n223), .A2(new_n224), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT1), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n234), .B1(G113gat), .B2(G120gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n232), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n227), .A2(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n219), .A2(new_n237), .ZN(new_n238));
  AND2_X1   g037(.A1(new_n206), .A2(new_n208), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n211), .A2(new_n213), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT77), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(new_n210), .ZN(new_n242));
  NAND2_X1  g041(.A1(KEYINPUT77), .A2(G162gat), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n212), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n239), .B(new_n240), .C1(new_n244), .C2(new_n207), .ZN(new_n245));
  AOI22_X1  g044(.A1(new_n245), .A2(new_n215), .B1(new_n236), .B2(new_n227), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n203), .B1(new_n238), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT79), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XOR2_X1   g048(.A(KEYINPUT78), .B(KEYINPUT3), .Z(new_n250));
  OAI211_X1 g049(.A(new_n215), .B(new_n250), .C1(new_n217), .C2(new_n218), .ZN(new_n251));
  AND2_X1   g050(.A1(KEYINPUT77), .A2(G162gat), .ZN(new_n252));
  NOR2_X1   g051(.A1(KEYINPUT77), .A2(G162gat), .ZN(new_n253));
  OAI21_X1  g052(.A(G155gat), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT2), .ZN(new_n255));
  AND4_X1   g054(.A1(new_n211), .A2(new_n206), .A3(new_n213), .A4(new_n208), .ZN(new_n256));
  AOI22_X1  g055(.A1(new_n255), .A2(new_n256), .B1(new_n214), .B2(new_n209), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT3), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n251), .B(new_n237), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n260), .B1(new_n219), .B2(new_n237), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n232), .A2(new_n235), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n225), .B1(new_n223), .B2(new_n224), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n262), .A2(new_n222), .B1(new_n263), .B2(new_n232), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n257), .A2(new_n264), .A3(KEYINPUT4), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n259), .A2(new_n202), .A3(new_n261), .A4(new_n265), .ZN(new_n266));
  OAI211_X1 g065(.A(KEYINPUT79), .B(new_n203), .C1(new_n238), .C2(new_n246), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n249), .A2(KEYINPUT5), .A3(new_n266), .A4(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT80), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT5), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n270), .B1(new_n247), .B2(new_n248), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT80), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n271), .A2(new_n272), .A3(new_n266), .A4(new_n267), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  OR2_X1    g073(.A1(new_n266), .A2(KEYINPUT5), .ZN(new_n275));
  XOR2_X1   g074(.A(G1gat), .B(G29gat), .Z(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(KEYINPUT0), .ZN(new_n277));
  XNOR2_X1  g076(.A(G57gat), .B(G85gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n274), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n274), .A2(new_n275), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n279), .B1(new_n285), .B2(KEYINPUT87), .ZN(new_n286));
  INV_X1    g085(.A(new_n275), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n287), .B1(new_n269), .B2(new_n273), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT87), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n284), .B1(new_n286), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n279), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n285), .A2(KEYINPUT6), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT22), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G211gat), .A2(G218gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(KEYINPUT72), .A2(KEYINPUT22), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G197gat), .B(G204gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AND2_X1   g100(.A1(G211gat), .A2(G218gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(G211gat), .A2(G218gat), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT73), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OR2_X1    g103(.A1(G211gat), .A2(G218gat), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT73), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n305), .A2(new_n306), .A3(new_n297), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n301), .A2(new_n304), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT74), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n305), .A2(new_n297), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n299), .A2(new_n310), .A3(new_n300), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT74), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n301), .A2(new_n312), .A3(new_n304), .A4(new_n307), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n309), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(G226gat), .A2(G233gat), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT66), .ZN(new_n318));
  INV_X1    g117(.A(G190gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT64), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT64), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(G190gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT28), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n320), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT27), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT27), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n327), .A2(KEYINPUT65), .A3(G183gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n324), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT64), .B(G190gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(KEYINPUT27), .B(G183gat), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n323), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n318), .B1(new_n330), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G183gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT27), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n327), .A2(G183gat), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n320), .A2(new_n322), .A3(new_n336), .A4(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT28), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n331), .A2(new_n323), .A3(new_n326), .A4(new_n328), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n339), .A2(KEYINPUT66), .A3(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT67), .ZN(new_n343));
  NAND2_X1  g142(.A1(G169gat), .A2(G176gat), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT67), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n345), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT26), .ZN(new_n347));
  INV_X1    g146(.A(G169gat), .ZN(new_n348));
  INV_X1    g147(.A(G176gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n343), .A2(new_n344), .A3(new_n346), .A4(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(G183gat), .A2(G190gat), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n334), .A2(new_n341), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT25), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n352), .A2(KEYINPUT24), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT24), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n357), .A2(G183gat), .A3(G190gat), .ZN(new_n358));
  AOI22_X1  g157(.A1(new_n356), .A2(new_n358), .B1(new_n335), .B2(new_n319), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n348), .A2(new_n349), .A3(KEYINPUT23), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT23), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n361), .B1(G169gat), .B2(G176gat), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n360), .A2(new_n362), .A3(new_n344), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n355), .B1(new_n359), .B2(new_n363), .ZN(new_n364));
  OR2_X1    g163(.A1(new_n363), .A2(new_n355), .ZN(new_n365));
  AOI22_X1  g164(.A1(new_n331), .A2(new_n335), .B1(new_n356), .B2(new_n358), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n354), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT29), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n317), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n316), .B1(new_n354), .B2(new_n367), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n315), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n368), .A2(new_n317), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT29), .B1(new_n354), .B2(new_n367), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n373), .B(new_n314), .C1(new_n317), .C2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(G8gat), .B(G36gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(G64gat), .B(G92gat), .ZN(new_n377));
  XOR2_X1   g176(.A(new_n376), .B(new_n377), .Z(new_n378));
  NAND3_X1  g177(.A1(new_n372), .A2(new_n375), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT38), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n372), .A2(new_n380), .A3(new_n375), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n380), .B1(new_n372), .B2(new_n375), .ZN(new_n382));
  OAI22_X1  g181(.A1(new_n381), .A2(new_n382), .B1(KEYINPUT37), .B2(new_n378), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n372), .A2(new_n375), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT38), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n378), .A2(KEYINPUT37), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n372), .A2(new_n380), .A3(new_n375), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n293), .A2(new_n379), .A3(new_n383), .A4(new_n388), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n291), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(G78gat), .B(G106gat), .ZN(new_n391));
  XOR2_X1   g190(.A(new_n391), .B(KEYINPUT83), .Z(new_n392));
  NAND2_X1  g191(.A1(G228gat), .A2(G233gat), .ZN(new_n393));
  XOR2_X1   g192(.A(new_n393), .B(KEYINPUT84), .Z(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT29), .B1(new_n257), .B2(new_n250), .ZN(new_n396));
  OR2_X1    g195(.A1(new_n314), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n310), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n301), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n399), .A2(KEYINPUT85), .A3(new_n311), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n310), .B1(new_n299), .B2(new_n300), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT85), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT29), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n250), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(new_n219), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n395), .B1(new_n397), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n313), .A2(new_n311), .ZN(new_n408));
  AND2_X1   g207(.A1(new_n307), .A2(new_n304), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n312), .B1(new_n409), .B2(new_n301), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n369), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n257), .B1(new_n411), .B2(new_n258), .ZN(new_n412));
  INV_X1    g211(.A(new_n393), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n413), .B1(new_n314), .B2(new_n396), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n407), .A2(new_n415), .A3(G22gat), .ZN(new_n416));
  INV_X1    g215(.A(G22gat), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT3), .B1(new_n314), .B2(new_n369), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n397), .B(new_n413), .C1(new_n418), .C2(new_n257), .ZN(new_n419));
  INV_X1    g218(.A(new_n250), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n420), .B1(new_n400), .B2(new_n403), .ZN(new_n421));
  OAI22_X1  g220(.A1(new_n421), .A2(new_n257), .B1(new_n314), .B2(new_n396), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(new_n394), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n417), .B1(new_n419), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n392), .B1(new_n416), .B2(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT31), .B(G50gat), .ZN(new_n426));
  OAI21_X1  g225(.A(G22gat), .B1(new_n407), .B2(new_n415), .ZN(new_n427));
  INV_X1    g226(.A(new_n392), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n419), .A2(new_n417), .A3(new_n423), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n425), .A2(new_n426), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n426), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n428), .B1(new_n427), .B2(new_n429), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n292), .B1(new_n288), .B2(new_n289), .ZN(new_n436));
  AOI211_X1 g235(.A(KEYINPUT87), .B(new_n287), .C1(new_n269), .C2(new_n273), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  XNOR2_X1  g237(.A(KEYINPUT76), .B(KEYINPUT30), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n379), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n378), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n384), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n372), .A2(KEYINPUT30), .A3(new_n375), .A4(new_n378), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n440), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n259), .A2(new_n261), .A3(new_n265), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n203), .ZN(new_n446));
  OR3_X1    g245(.A1(new_n238), .A2(new_n246), .A3(new_n203), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n446), .A2(KEYINPUT39), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n279), .B1(new_n446), .B2(KEYINPUT39), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT40), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OR2_X1    g250(.A1(new_n446), .A2(KEYINPUT39), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT40), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n452), .A2(new_n453), .A3(new_n279), .A4(new_n448), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n444), .A2(new_n455), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n431), .B(new_n435), .C1(new_n438), .C2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT88), .B1(new_n390), .B2(new_n457), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n383), .A2(new_n388), .A3(new_n379), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT6), .B1(new_n274), .B2(new_n281), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n460), .B1(new_n436), .B2(new_n437), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n459), .A2(new_n461), .A3(new_n293), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n435), .A2(new_n431), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT88), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n444), .B(new_n455), .C1(new_n436), .C2(new_n437), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n462), .A2(new_n464), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n458), .A2(new_n467), .ZN(new_n468));
  XOR2_X1   g267(.A(G15gat), .B(G43gat), .Z(new_n469));
  XNOR2_X1  g268(.A(G71gat), .B(G99gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n469), .B(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n368), .A2(new_n264), .ZN(new_n473));
  NAND2_X1  g272(.A1(G227gat), .A2(G233gat), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n354), .A2(new_n237), .A3(new_n367), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n473), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(KEYINPUT69), .B(KEYINPUT33), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n472), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n473), .A2(new_n476), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT34), .B1(new_n475), .B2(KEYINPUT70), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n481), .A2(new_n474), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n482), .B1(new_n481), .B2(new_n474), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n480), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n483), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n479), .B1(new_n487), .B2(new_n484), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n477), .A2(KEYINPUT32), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n490), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n486), .A2(new_n488), .A3(new_n492), .ZN(new_n493));
  NOR2_X1   g292(.A1(KEYINPUT71), .A2(KEYINPUT36), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT71), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT36), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n491), .B(new_n493), .C1(new_n494), .C2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n493), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n492), .B1(new_n486), .B2(new_n488), .ZN(new_n500));
  OAI22_X1  g299(.A1(new_n499), .A2(new_n500), .B1(new_n495), .B2(new_n496), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n435), .A2(KEYINPUT86), .A3(new_n431), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT86), .B1(new_n435), .B2(new_n431), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n442), .A2(KEYINPUT75), .A3(new_n443), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT75), .B1(new_n442), .B2(new_n443), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n440), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT81), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n460), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT82), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n285), .A2(new_n511), .A3(new_n292), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n280), .B1(new_n269), .B2(new_n273), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT81), .B1(new_n513), .B2(KEYINPUT6), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT82), .B1(new_n288), .B2(new_n279), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n510), .A2(new_n512), .A3(new_n514), .A4(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n508), .B1(new_n516), .B2(new_n293), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n502), .B1(new_n505), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT35), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n491), .A2(new_n435), .A3(new_n431), .A4(new_n493), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n519), .B1(new_n517), .B2(new_n521), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n461), .A2(new_n293), .ZN(new_n523));
  INV_X1    g322(.A(new_n444), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(new_n519), .ZN(new_n525));
  NOR3_X1   g324(.A1(new_n523), .A2(new_n520), .A3(new_n525), .ZN(new_n526));
  OAI22_X1  g325(.A1(new_n468), .A2(new_n518), .B1(new_n522), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(G113gat), .B(G141gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(G197gat), .ZN(new_n529));
  XOR2_X1   g328(.A(KEYINPUT11), .B(G169gat), .Z(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  XOR2_X1   g330(.A(new_n531), .B(KEYINPUT12), .Z(new_n532));
  XNOR2_X1  g331(.A(G43gat), .B(G50gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT15), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(G29gat), .A2(G36gat), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NOR3_X1   g337(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n536), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  XOR2_X1   g340(.A(G43gat), .B(G50gat), .Z(new_n542));
  INV_X1    g341(.A(KEYINPUT15), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n536), .B(KEYINPUT90), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(new_n534), .A3(new_n545), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n539), .A2(KEYINPUT89), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n539), .A2(KEYINPUT89), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n538), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n541), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT17), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT91), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n550), .A2(KEYINPUT91), .A3(new_n551), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT94), .ZN(new_n557));
  INV_X1    g356(.A(new_n550), .ZN(new_n558));
  XNOR2_X1  g357(.A(G15gat), .B(G22gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT92), .ZN(new_n560));
  INV_X1    g359(.A(G1gat), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT16), .ZN(new_n562));
  AOI22_X1  g361(.A1(new_n560), .A2(new_n561), .B1(new_n562), .B2(new_n559), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n559), .A2(KEYINPUT92), .A3(G1gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT93), .ZN(new_n566));
  OR2_X1    g365(.A1(new_n566), .A2(G8gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(G8gat), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n565), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n563), .A2(new_n566), .A3(G8gat), .A4(new_n564), .ZN(new_n570));
  AOI22_X1  g369(.A1(new_n558), .A2(KEYINPUT17), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n556), .A2(new_n557), .A3(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n569), .A2(new_n550), .A3(new_n570), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(G229gat), .A2(G233gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n556), .A2(new_n571), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT94), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n574), .A2(KEYINPUT18), .A3(new_n575), .A4(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n569), .A2(new_n570), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(new_n558), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n573), .A2(KEYINPUT96), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n575), .B(KEYINPUT13), .Z(new_n585));
  NAND2_X1  g384(.A1(new_n581), .A2(new_n582), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n578), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n577), .A2(new_n575), .A3(new_n573), .A4(new_n572), .ZN(new_n589));
  XNOR2_X1  g388(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n532), .B1(new_n588), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n532), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n591), .A2(new_n578), .A3(new_n594), .A4(new_n587), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n527), .A2(new_n596), .ZN(new_n597));
  OR2_X1    g396(.A1(G57gat), .A2(G64gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(G57gat), .A2(G64gat), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n598), .A2(KEYINPUT97), .A3(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G71gat), .B(G78gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(G71gat), .ZN(new_n603));
  INV_X1    g402(.A(G78gat), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n605), .A2(KEYINPUT9), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n602), .A2(new_n606), .A3(new_n598), .A4(new_n599), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n598), .B(new_n599), .C1(new_n605), .C2(KEYINPUT9), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n608), .A2(new_n601), .A3(new_n600), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n610), .A2(KEYINPUT21), .ZN(new_n611));
  NAND2_X1  g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(G127gat), .B(G155gat), .Z(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT20), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n613), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT21), .ZN(new_n619));
  INV_X1    g418(.A(new_n610), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n579), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(new_n621), .B(KEYINPUT99), .Z(new_n622));
  NAND2_X1  g421(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n621), .B(KEYINPUT99), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n624), .A2(new_n617), .A3(new_n616), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G183gat), .B(G211gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT98), .B(KEYINPUT19), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n627), .B(new_n628), .Z(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n623), .A2(new_n625), .A3(new_n629), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(G232gat), .A2(G233gat), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(KEYINPUT41), .ZN(new_n636));
  NAND2_X1  g435(.A1(G99gat), .A2(G106gat), .ZN(new_n637));
  INV_X1    g436(.A(G85gat), .ZN(new_n638));
  INV_X1    g437(.A(G92gat), .ZN(new_n639));
  AOI22_X1  g438(.A1(KEYINPUT8), .A2(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT7), .ZN(new_n641));
  OAI22_X1  g440(.A1(new_n638), .A2(new_n639), .B1(new_n641), .B2(KEYINPUT101), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT101), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n643), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n640), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g444(.A(G99gat), .B(G106gat), .Z(new_n646));
  OR2_X1    g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n636), .B1(new_n558), .B2(new_n649), .ZN(new_n650));
  AOI22_X1  g449(.A1(new_n558), .A2(KEYINPUT17), .B1(new_n647), .B2(new_n648), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n650), .B1(new_n556), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(G190gat), .B(G218gat), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n652), .A2(new_n654), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g457(.A(G134gat), .B(G162gat), .Z(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT100), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n635), .A2(KEYINPUT41), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n662), .B1(new_n655), .B2(KEYINPUT102), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n658), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n656), .A2(new_n657), .A3(KEYINPUT102), .A4(new_n662), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(G230gat), .A2(G233gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT104), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n646), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n645), .A2(new_n670), .A3(KEYINPUT103), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n645), .A2(KEYINPUT103), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(new_n646), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n610), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n647), .A2(new_n607), .A3(new_n609), .A4(new_n648), .ZN(new_n675));
  AOI21_X1  g474(.A(KEYINPUT10), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n610), .A2(KEYINPUT10), .A3(new_n647), .A4(new_n648), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n669), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n674), .A2(new_n675), .ZN(new_n680));
  INV_X1    g479(.A(new_n667), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(G120gat), .B(G148gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(G176gat), .B(G204gat), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n684), .B(new_n685), .Z(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n687), .B1(new_n680), .B2(new_n681), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n667), .B1(new_n676), .B2(new_n678), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n633), .A2(new_n666), .A3(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n597), .A2(new_n694), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n516), .A2(new_n293), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g497(.A1(new_n695), .A2(new_n444), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT16), .B(G8gat), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT105), .ZN(new_n702));
  AND3_X1   g501(.A1(new_n701), .A2(new_n702), .A3(KEYINPUT42), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n699), .A2(G8gat), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT42), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n705), .B1(new_n699), .B2(new_n700), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n702), .B1(new_n701), .B2(KEYINPUT42), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n703), .B1(new_n706), .B2(new_n707), .ZN(G1325gat));
  INV_X1    g507(.A(new_n695), .ZN(new_n709));
  OAI21_X1  g508(.A(G15gat), .B1(new_n709), .B2(new_n502), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n499), .A2(new_n500), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  OR2_X1    g511(.A1(new_n712), .A2(G15gat), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n710), .B1(new_n709), .B2(new_n713), .ZN(G1326gat));
  INV_X1    g513(.A(KEYINPUT86), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n463), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n435), .A2(KEYINPUT86), .A3(new_n431), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n695), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(KEYINPUT43), .B(G22gat), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(G1327gat));
  INV_X1    g520(.A(new_n586), .ZN(new_n722));
  INV_X1    g521(.A(new_n585), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n722), .A2(new_n583), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n572), .A2(new_n573), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n557), .B1(new_n556), .B2(new_n571), .ZN(new_n726));
  INV_X1    g525(.A(new_n575), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n724), .B1(new_n728), .B2(KEYINPUT18), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n594), .B1(new_n729), .B2(new_n591), .ZN(new_n730));
  INV_X1    g529(.A(new_n595), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n718), .B1(new_n696), .B2(new_n508), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n733), .A2(new_n502), .A3(new_n458), .A4(new_n467), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n517), .A2(new_n521), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(KEYINPUT35), .ZN(new_n736));
  OR3_X1    g535(.A1(new_n523), .A2(new_n520), .A3(new_n525), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n732), .B1(new_n734), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n633), .A2(new_n692), .ZN(new_n740));
  INV_X1    g539(.A(new_n666), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n740), .A2(KEYINPUT106), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT106), .B1(new_n740), .B2(new_n741), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n739), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n696), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n745), .A2(G29gat), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT44), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n750), .B1(new_n527), .B2(new_n741), .ZN(new_n751));
  AND3_X1   g550(.A1(new_n664), .A2(KEYINPUT108), .A3(new_n665), .ZN(new_n752));
  AOI21_X1  g551(.A(KEYINPUT108), .B1(new_n664), .B2(new_n665), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n750), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n755), .B1(new_n734), .B2(new_n738), .ZN(new_n756));
  OR2_X1    g555(.A1(new_n751), .A2(new_n756), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n732), .A2(new_n633), .A3(new_n692), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n757), .A2(new_n696), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G29gat), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n749), .A2(new_n760), .ZN(G1328gat));
  NOR3_X1   g560(.A1(new_n745), .A2(G36gat), .A3(new_n524), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT46), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n757), .A2(new_n444), .A3(new_n758), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(G36gat), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(G1329gat));
  INV_X1    g565(.A(new_n502), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n767), .B(new_n758), .C1(new_n751), .C2(new_n756), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(G43gat), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n712), .A2(G43gat), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n527), .A2(new_n596), .A3(new_n744), .A4(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n769), .A2(KEYINPUT47), .A3(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT109), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n739), .A2(KEYINPUT109), .A3(new_n744), .A4(new_n770), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n769), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT47), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT110), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT110), .ZN(new_n780));
  AOI211_X1 g579(.A(new_n780), .B(KEYINPUT47), .C1(new_n769), .C2(new_n776), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n772), .B1(new_n779), .B2(new_n781), .ZN(G1330gat));
  OR2_X1    g581(.A1(new_n505), .A2(G50gat), .ZN(new_n783));
  OAI21_X1  g582(.A(KEYINPUT48), .B1(new_n745), .B2(new_n783), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n463), .B(new_n758), .C1(new_n751), .C2(new_n756), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n784), .B1(G50gat), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT111), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AOI211_X1 g587(.A(KEYINPUT111), .B(new_n784), .C1(new_n785), .C2(G50gat), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n745), .A2(new_n783), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n757), .A2(new_n718), .A3(new_n758), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n790), .B1(new_n791), .B2(G50gat), .ZN(new_n792));
  OAI22_X1  g591(.A1(new_n788), .A2(new_n789), .B1(new_n792), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g592(.A(new_n633), .ZN(new_n794));
  NOR4_X1   g593(.A1(new_n794), .A2(new_n596), .A3(new_n741), .A4(new_n693), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n527), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n696), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g598(.A1(new_n797), .A2(KEYINPUT112), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT112), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n796), .A2(new_n801), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n804));
  AND2_X1   g603(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n803), .B(new_n444), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n803), .A2(new_n444), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n806), .B1(new_n807), .B2(new_n804), .ZN(G1333gat));
  AND3_X1   g607(.A1(new_n797), .A2(KEYINPUT113), .A3(new_n711), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT113), .B1(new_n797), .B2(new_n711), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n603), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n800), .A2(new_n767), .A3(new_n802), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(G71gat), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT50), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n811), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n814), .B1(new_n811), .B2(new_n813), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n815), .A2(new_n816), .ZN(G1334gat));
  NAND2_X1  g616(.A1(new_n803), .A2(new_n718), .ZN(new_n818));
  XNOR2_X1  g617(.A(KEYINPUT114), .B(G78gat), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n818), .B(new_n819), .ZN(G1335gat));
  AOI21_X1  g619(.A(new_n666), .B1(new_n734), .B2(new_n738), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n596), .A2(new_n633), .ZN(new_n822));
  AND3_X1   g621(.A1(new_n821), .A2(KEYINPUT51), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT51), .B1(new_n821), .B2(new_n822), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n826), .A2(new_n638), .A3(new_n696), .A4(new_n692), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT115), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n596), .A2(new_n633), .A3(new_n693), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n757), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n828), .B1(new_n830), .B2(new_n746), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(G85gat), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n830), .A2(new_n828), .A3(new_n746), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n827), .B1(new_n832), .B2(new_n833), .ZN(G1336gat));
  OAI211_X1 g633(.A(new_n444), .B(new_n829), .C1(new_n751), .C2(new_n756), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(G92gat), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n524), .A2(G92gat), .A3(new_n693), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n836), .B1(new_n825), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(KEYINPUT52), .ZN(G1337gat));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n841), .B1(new_n830), .B2(new_n502), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(G99gat), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n830), .A2(new_n841), .A3(new_n502), .ZN(new_n844));
  OR3_X1    g643(.A1(new_n712), .A2(G99gat), .A3(new_n693), .ZN(new_n845));
  OAI22_X1  g644(.A1(new_n843), .A2(new_n844), .B1(new_n825), .B2(new_n845), .ZN(G1338gat));
  OAI21_X1  g645(.A(G106gat), .B1(new_n830), .B2(new_n464), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT53), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n464), .A2(G106gat), .A3(new_n693), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n849), .B1(new_n823), .B2(new_n824), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n847), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n849), .B(KEYINPUT117), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n757), .A2(new_n718), .A3(new_n829), .ZN(new_n853));
  AOI22_X1  g652(.A1(new_n826), .A2(new_n852), .B1(new_n853), .B2(G106gat), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n851), .B1(new_n854), .B2(new_n848), .ZN(G1339gat));
  NOR2_X1   g654(.A1(new_n694), .A2(new_n596), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n857), .B(new_n669), .C1(new_n676), .C2(new_n678), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n687), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n668), .B(new_n677), .C1(new_n680), .C2(KEYINPUT10), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(KEYINPUT54), .A3(new_n690), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(KEYINPUT118), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT118), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n860), .A2(new_n863), .A3(new_n690), .A4(KEYINPUT54), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n859), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n691), .B1(new_n865), .B2(KEYINPUT55), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n862), .A2(new_n864), .ZN(new_n867));
  INV_X1    g666(.A(new_n859), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(KEYINPUT55), .A3(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT119), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n865), .A2(KEYINPUT119), .A3(KEYINPUT55), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n866), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n575), .B1(new_n574), .B2(new_n577), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n585), .B1(new_n584), .B2(new_n586), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n531), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n595), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n754), .A2(new_n873), .A3(new_n877), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n595), .A2(new_n876), .A3(new_n692), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n879), .B1(new_n873), .B2(new_n596), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n878), .B1(new_n880), .B2(new_n754), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n856), .B1(new_n881), .B2(new_n794), .ZN(new_n882));
  NOR4_X1   g681(.A1(new_n882), .A2(new_n746), .A3(new_n520), .A4(new_n444), .ZN(new_n883));
  AOI21_X1  g682(.A(G113gat), .B1(new_n883), .B2(new_n596), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n696), .A2(new_n524), .ZN(new_n885));
  NOR4_X1   g684(.A1(new_n882), .A2(new_n712), .A3(new_n718), .A4(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n732), .A2(new_n223), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n884), .B1(new_n886), .B2(new_n887), .ZN(G1340gat));
  NOR2_X1   g687(.A1(new_n220), .A2(new_n221), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n883), .A2(new_n889), .A3(new_n692), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n886), .A2(new_n692), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n890), .B1(new_n891), .B2(new_n224), .ZN(G1341gat));
  NAND3_X1  g691(.A1(new_n883), .A2(new_n230), .A3(new_n633), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n886), .A2(new_n633), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n893), .B1(new_n894), .B2(new_n230), .ZN(G1342gat));
  NAND3_X1  g694(.A1(new_n883), .A2(new_n228), .A3(new_n741), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n896), .A2(KEYINPUT56), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(KEYINPUT56), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n886), .A2(new_n741), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n897), .B(new_n898), .C1(new_n228), .C2(new_n899), .ZN(G1343gat));
  INV_X1    g699(.A(KEYINPUT57), .ZN(new_n901));
  INV_X1    g700(.A(new_n879), .ZN(new_n902));
  INV_X1    g701(.A(new_n866), .ZN(new_n903));
  INV_X1    g702(.A(new_n872), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT119), .B1(new_n865), .B2(KEYINPUT55), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n902), .B1(new_n906), .B2(new_n732), .ZN(new_n907));
  INV_X1    g706(.A(new_n754), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n633), .B1(new_n909), .B2(new_n878), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n901), .B(new_n463), .C1(new_n910), .C2(new_n856), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n878), .B1(new_n880), .B2(new_n741), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n856), .B1(new_n912), .B2(new_n794), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT57), .B1(new_n913), .B2(new_n505), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n767), .A2(new_n885), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n911), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(G141gat), .B1(new_n916), .B2(new_n732), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n882), .A2(new_n746), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n767), .A2(new_n464), .A3(new_n444), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n596), .A2(new_n204), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n917), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(KEYINPUT58), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT58), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n917), .B(new_n924), .C1(new_n920), .C2(new_n921), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(G1344gat));
  INV_X1    g725(.A(KEYINPUT122), .ZN(new_n927));
  OAI21_X1  g726(.A(KEYINPUT57), .B1(new_n882), .B2(new_n464), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n505), .A2(KEYINPUT57), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n907), .A2(new_n666), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n873), .A2(new_n741), .A3(new_n877), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n633), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n929), .B1(new_n932), .B2(new_n856), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT121), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n915), .A2(new_n934), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n767), .A2(new_n885), .A3(KEYINPUT121), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n935), .A2(new_n693), .A3(new_n936), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n928), .A2(new_n933), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(G148gat), .ZN(new_n939));
  XNOR2_X1  g738(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n911), .A2(new_n914), .A3(new_n692), .A4(new_n915), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n205), .A2(KEYINPUT59), .ZN(new_n942));
  AOI22_X1  g741(.A1(new_n939), .A2(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n920), .A2(G148gat), .A3(new_n693), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n927), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(new_n944), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n941), .A2(new_n942), .ZN(new_n947));
  INV_X1    g746(.A(new_n940), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n948), .B1(new_n938), .B2(G148gat), .ZN(new_n949));
  OAI211_X1 g748(.A(KEYINPUT122), .B(new_n946), .C1(new_n947), .C2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n945), .A2(new_n950), .ZN(G1345gat));
  OAI21_X1  g750(.A(G155gat), .B1(new_n916), .B2(new_n794), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n633), .A2(new_n212), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n952), .B1(new_n920), .B2(new_n953), .ZN(G1346gat));
  OAI21_X1  g753(.A(new_n216), .B1(new_n916), .B2(new_n908), .ZN(new_n955));
  OR2_X1    g754(.A1(new_n666), .A2(new_n216), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n955), .B1(new_n920), .B2(new_n956), .ZN(G1347gat));
  NOR2_X1   g756(.A1(new_n882), .A2(new_n696), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n520), .A2(new_n524), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g760(.A(G169gat), .B1(new_n961), .B2(new_n596), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n746), .A2(new_n444), .ZN(new_n963));
  NOR4_X1   g762(.A1(new_n882), .A2(new_n712), .A3(new_n718), .A4(new_n963), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n732), .A2(new_n348), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n962), .B1(new_n964), .B2(new_n965), .ZN(G1348gat));
  NAND3_X1  g765(.A1(new_n961), .A2(new_n349), .A3(new_n692), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n964), .A2(new_n692), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n967), .B1(new_n968), .B2(new_n349), .ZN(G1349gat));
  INV_X1    g768(.A(KEYINPUT123), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(KEYINPUT60), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n633), .A2(new_n332), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n971), .B1(new_n960), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n335), .B1(new_n964), .B2(new_n633), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n970), .A2(KEYINPUT60), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n975), .B(new_n976), .ZN(G1350gat));
  NAND3_X1  g776(.A1(new_n961), .A2(new_n331), .A3(new_n754), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT61), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n741), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n979), .B1(new_n980), .B2(G190gat), .ZN(new_n981));
  AOI211_X1 g780(.A(KEYINPUT61), .B(new_n319), .C1(new_n964), .C2(new_n741), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n978), .B1(new_n981), .B2(new_n982), .ZN(G1351gat));
  INV_X1    g782(.A(KEYINPUT125), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n502), .A2(new_n463), .A3(new_n444), .ZN(new_n985));
  XOR2_X1   g784(.A(new_n985), .B(KEYINPUT124), .Z(new_n986));
  AND3_X1   g785(.A1(new_n958), .A2(new_n984), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n984), .B1(new_n958), .B2(new_n986), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g788(.A(G197gat), .B1(new_n989), .B2(new_n596), .ZN(new_n990));
  AND2_X1   g789(.A1(new_n928), .A2(new_n933), .ZN(new_n991));
  NOR2_X1   g790(.A1(new_n963), .A2(new_n767), .ZN(new_n992));
  AND2_X1   g791(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AND2_X1   g792(.A1(new_n596), .A2(G197gat), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n990), .B1(new_n993), .B2(new_n994), .ZN(G1352gat));
  NAND3_X1  g794(.A1(new_n991), .A2(new_n692), .A3(new_n992), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n996), .A2(G204gat), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n958), .A2(new_n986), .ZN(new_n998));
  NOR2_X1   g797(.A1(new_n693), .A2(G204gat), .ZN(new_n999));
  INV_X1    g798(.A(new_n999), .ZN(new_n1000));
  OR3_X1    g799(.A1(new_n998), .A2(KEYINPUT126), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g800(.A(KEYINPUT62), .ZN(new_n1002));
  OAI21_X1  g801(.A(KEYINPUT126), .B1(new_n998), .B2(new_n1000), .ZN(new_n1003));
  AND3_X1   g802(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g803(.A(new_n1002), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1005));
  OAI21_X1  g804(.A(new_n997), .B1(new_n1004), .B2(new_n1005), .ZN(G1353gat));
  NAND4_X1  g805(.A1(new_n928), .A2(new_n933), .A3(new_n633), .A4(new_n992), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1007), .A2(G211gat), .ZN(new_n1008));
  OR2_X1    g807(.A1(new_n1008), .A2(KEYINPUT63), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1008), .A2(KEYINPUT63), .ZN(new_n1010));
  INV_X1    g809(.A(KEYINPUT127), .ZN(new_n1011));
  NOR2_X1   g810(.A1(new_n794), .A2(G211gat), .ZN(new_n1012));
  AND3_X1   g811(.A1(new_n989), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g812(.A(new_n1011), .B1(new_n989), .B2(new_n1012), .ZN(new_n1014));
  OAI211_X1 g813(.A(new_n1009), .B(new_n1010), .C1(new_n1013), .C2(new_n1014), .ZN(G1354gat));
  NAND3_X1  g814(.A1(new_n991), .A2(new_n741), .A3(new_n992), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1016), .A2(G218gat), .ZN(new_n1017));
  INV_X1    g816(.A(new_n989), .ZN(new_n1018));
  OR2_X1    g817(.A1(new_n908), .A2(G218gat), .ZN(new_n1019));
  OAI21_X1  g818(.A(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(G1355gat));
endmodule


