//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 1 0 1 0 0 0 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 1 1 1 1 0 0 0 0 0 1 1 0 1 1 0 1 0 0 0 1 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1214, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1276, new_n1277, new_n1278;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  AOI22_X1  g0005(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT65), .ZN(new_n207));
  INV_X1    g0007(.A(G50), .ZN(new_n208));
  INV_X1    g0008(.A(G226), .ZN(new_n209));
  INV_X1    g0009(.A(G68), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  OAI22_X1  g0011(.A1(new_n208), .A2(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI21_X1  g0012(.A(new_n212), .B1(G77), .B2(G244), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n207), .B(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n216), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n217), .B1(new_n202), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G20), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT66), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n220), .A2(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT0), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n223), .B(new_n226), .C1(KEYINPUT1), .C2(new_n221), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(G58), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(new_n210), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G50), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT64), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n227), .B1(new_n230), .B2(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT67), .ZN(G361));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G264), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n238), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n239), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT68), .ZN(new_n246));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G107), .B(G116), .Z(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  INV_X1    g0052(.A(KEYINPUT70), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n253), .B1(new_n220), .B2(new_n254), .ZN(new_n255));
  NAND4_X1  g0055(.A1(KEYINPUT70), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n255), .A2(new_n228), .A3(new_n256), .ZN(new_n257));
  AND2_X1   g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n229), .B(G87), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT22), .ZN(new_n261));
  OR2_X1    g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT22), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n264), .A2(new_n265), .A3(new_n229), .A4(G87), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G33), .A2(G116), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n261), .A2(new_n266), .B1(new_n229), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT24), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n229), .A2(G107), .ZN(new_n271));
  XNOR2_X1  g0071(.A(new_n271), .B(KEYINPUT23), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n269), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n270), .B1(new_n269), .B2(new_n272), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n257), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n215), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n218), .A2(G1698), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n278), .B(new_n279), .C1(new_n258), .C2(new_n259), .ZN(new_n280));
  XOR2_X1   g0080(.A(KEYINPUT85), .B(G294), .Z(new_n281));
  OAI21_X1  g0081(.A(new_n280), .B1(new_n281), .B2(new_n254), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G45), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n285), .A2(G1), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT5), .B(G41), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n283), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G264), .ZN(new_n289));
  INV_X1    g0089(.A(G190), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n287), .A2(G274), .A3(new_n286), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n284), .A2(new_n289), .A3(new_n290), .A4(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT86), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n282), .A2(new_n283), .B1(new_n288), .B2(G264), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT86), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n294), .A2(new_n295), .A3(new_n290), .A4(new_n291), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n284), .A2(new_n291), .A3(new_n289), .ZN(new_n297));
  INV_X1    g0097(.A(G200), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n293), .A2(new_n296), .A3(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n257), .ZN(new_n301));
  INV_X1    g0101(.A(G13), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(G1), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G20), .ZN(new_n304));
  INV_X1    g0104(.A(G1), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G33), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n301), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n307), .A2(new_n203), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n303), .A2(new_n271), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n309), .B(KEYINPUT25), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n276), .A2(new_n300), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(G169), .B1(new_n294), .B2(new_n291), .ZN(new_n313));
  INV_X1    g0113(.A(G179), .ZN(new_n314));
  AND4_X1   g0114(.A1(new_n314), .A2(new_n284), .A3(new_n291), .A4(new_n289), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n261), .A2(new_n266), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n268), .A2(new_n229), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n317), .A2(new_n272), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT24), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n301), .B1(new_n320), .B2(new_n273), .ZN(new_n321));
  INV_X1    g0121(.A(new_n311), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n316), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n312), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT87), .ZN(new_n325));
  INV_X1    g0125(.A(new_n303), .ZN(new_n326));
  INV_X1    g0126(.A(G116), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G20), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(G33), .A2(G283), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n330), .B(new_n229), .C1(G33), .C2(new_n202), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT83), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(G20), .B1(new_n254), .B2(G97), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n334), .A2(KEYINPUT83), .A3(new_n330), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n257), .A2(new_n333), .A3(new_n328), .A4(new_n335), .ZN(new_n336));
  XNOR2_X1  g0136(.A(KEYINPUT84), .B(KEYINPUT20), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n329), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AND2_X1   g0138(.A1(new_n333), .A2(new_n335), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT84), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n340), .A2(KEYINPUT20), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n339), .A2(new_n257), .A3(new_n341), .A4(new_n328), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n301), .A2(G116), .A3(new_n304), .A4(new_n306), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n338), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G264), .A2(G1698), .ZN(new_n345));
  OAI221_X1 g0145(.A(new_n345), .B1(new_n218), .B2(G1698), .C1(new_n258), .C2(new_n259), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n258), .A2(new_n259), .ZN(new_n347));
  INV_X1    g0147(.A(G303), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n346), .A2(new_n349), .A3(new_n283), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n287), .A2(new_n286), .ZN(new_n351));
  INV_X1    g0151(.A(G41), .ZN(new_n352));
  OAI211_X1 g0152(.A(G1), .B(G13), .C1(new_n254), .C2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n351), .A2(G270), .A3(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n350), .A2(new_n291), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n344), .A2(G179), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(G200), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(new_n290), .B2(new_n355), .ZN(new_n359));
  OR2_X1    g0159(.A1(new_n359), .A2(new_n344), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n344), .A2(G169), .A3(new_n355), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT21), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n344), .A2(KEYINPUT21), .A3(G169), .A4(new_n355), .ZN(new_n364));
  AND4_X1   g0164(.A1(new_n357), .A2(new_n360), .A3(new_n363), .A4(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(G274), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n286), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n215), .B1(new_n285), .B2(G1), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n367), .A2(new_n353), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n211), .A2(new_n277), .ZN(new_n370));
  INV_X1    g0170(.A(G244), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(G1698), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n370), .B(new_n372), .C1(new_n258), .C2(new_n259), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n373), .A2(new_n267), .ZN(new_n374));
  OAI211_X1 g0174(.A(G190), .B(new_n369), .C1(new_n374), .C2(new_n353), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n229), .B1(new_n254), .B2(new_n202), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n214), .A2(new_n202), .A3(new_n203), .ZN(new_n377));
  OR2_X1    g0177(.A1(KEYINPUT82), .A2(KEYINPUT19), .ZN(new_n378));
  NAND2_X1  g0178(.A1(KEYINPUT82), .A2(KEYINPUT19), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n376), .A2(new_n377), .A3(new_n378), .A4(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n378), .A2(new_n379), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n229), .A2(G33), .A3(G97), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n229), .B(G68), .C1(new_n258), .C2(new_n259), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n380), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n304), .ZN(new_n386));
  XOR2_X1   g0186(.A(KEYINPUT15), .B(G87), .Z(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n385), .A2(new_n257), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n353), .B1(new_n373), .B2(new_n267), .ZN(new_n390));
  AND3_X1   g0190(.A1(new_n367), .A2(new_n353), .A3(new_n368), .ZN(new_n391));
  OAI21_X1  g0191(.A(G200), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n301), .A2(G87), .A3(new_n304), .A4(new_n306), .ZN(new_n393));
  AND4_X1   g0193(.A1(new_n375), .A2(new_n389), .A3(new_n392), .A4(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n385), .A2(new_n257), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n301), .A2(new_n304), .A3(new_n387), .A4(new_n306), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n388), .A2(new_n386), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n390), .A2(new_n391), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT81), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(new_n400), .A3(new_n314), .ZN(new_n401));
  INV_X1    g0201(.A(G169), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(new_n390), .B2(new_n391), .ZN(new_n403));
  AND3_X1   g0203(.A1(new_n398), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n399), .A2(new_n314), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT81), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n394), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n264), .A2(G250), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n277), .B1(new_n408), .B2(KEYINPUT4), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT4), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n410), .A2(G1698), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n411), .B(G244), .C1(new_n259), .C2(new_n258), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n371), .B1(new_n262), .B2(new_n263), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n412), .B(new_n330), .C1(new_n413), .C2(KEYINPUT4), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n283), .B1(new_n409), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n288), .A2(G257), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n415), .A2(new_n291), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(G200), .ZN(new_n418));
  AOI21_X1  g0218(.A(KEYINPUT7), .B1(new_n347), .B2(new_n229), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT7), .ZN(new_n420));
  NOR4_X1   g0220(.A1(new_n258), .A2(new_n259), .A3(new_n420), .A4(G20), .ZN(new_n421));
  OAI21_X1  g0221(.A(G107), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n203), .A2(KEYINPUT6), .A3(G97), .ZN(new_n423));
  XOR2_X1   g0223(.A(G97), .B(G107), .Z(new_n424));
  OAI21_X1  g0224(.A(new_n423), .B1(new_n424), .B2(KEYINPUT6), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(G20), .ZN(new_n426));
  NOR3_X1   g0226(.A1(KEYINPUT71), .A2(G20), .A3(G33), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(KEYINPUT71), .B1(G20), .B2(G33), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(G77), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n422), .A2(new_n426), .A3(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n307), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n432), .A2(new_n257), .B1(new_n433), .B2(G97), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n386), .A2(new_n202), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n415), .A2(G190), .A3(new_n291), .A4(new_n416), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n418), .A2(new_n434), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n432), .A2(new_n257), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n433), .A2(G97), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(new_n435), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n417), .A2(new_n402), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n415), .A2(new_n314), .A3(new_n291), .A4(new_n416), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  AND3_X1   g0243(.A1(new_n407), .A2(new_n437), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT87), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n312), .A2(new_n323), .A3(new_n445), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n325), .A2(new_n365), .A3(new_n444), .A4(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n429), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n448), .A2(new_n427), .ZN(new_n449));
  INV_X1    g0249(.A(G150), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(G20), .B1(new_n232), .B2(G50), .ZN(new_n452));
  XNOR2_X1  g0252(.A(KEYINPUT8), .B(G58), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n254), .A2(G20), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n452), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n257), .B1(new_n451), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n386), .A2(new_n208), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n208), .B1(new_n305), .B2(G20), .ZN(new_n460));
  OR2_X1    g0260(.A1(new_n460), .A2(KEYINPUT72), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(KEYINPUT72), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n301), .A2(new_n461), .A3(new_n304), .A4(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT9), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n457), .A2(KEYINPUT9), .A3(new_n463), .A4(new_n458), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n277), .A2(G222), .ZN(new_n468));
  INV_X1    g0268(.A(G223), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n264), .B(new_n468), .C1(new_n469), .C2(new_n277), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n470), .B(new_n283), .C1(G77), .C2(new_n264), .ZN(new_n471));
  NOR2_X1   g0271(.A1(G41), .A2(G45), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n473), .A2(KEYINPUT69), .A3(new_n305), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT69), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n475), .B1(new_n472), .B2(G1), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n283), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G226), .ZN(new_n478));
  NOR3_X1   g0278(.A1(new_n472), .A2(G1), .A3(new_n366), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n471), .A2(new_n478), .A3(G190), .A4(new_n480), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n467), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT10), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n471), .A2(new_n480), .A3(new_n478), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G200), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n466), .A2(new_n482), .A3(new_n483), .A4(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n485), .A2(new_n467), .A3(new_n481), .ZN(new_n487));
  AOI21_X1  g0287(.A(KEYINPUT9), .B1(new_n459), .B2(new_n463), .ZN(new_n488));
  OAI21_X1  g0288(.A(KEYINPUT10), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(G238), .A2(G1698), .ZN(new_n491));
  INV_X1    g0291(.A(G232), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n264), .B(new_n491), .C1(new_n492), .C2(G1698), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n493), .B(new_n283), .C1(G107), .C2(new_n264), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n477), .A2(G244), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n494), .A2(new_n480), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n314), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n387), .A2(new_n454), .B1(G20), .B2(G77), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(new_n449), .B2(new_n453), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n257), .B1(new_n305), .B2(G20), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n500), .A2(new_n257), .B1(G77), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(G77), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n386), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n496), .A2(new_n402), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n498), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n494), .A2(G190), .A3(new_n495), .A4(new_n480), .ZN(new_n508));
  XNOR2_X1  g0308(.A(new_n508), .B(KEYINPUT73), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n504), .B(new_n502), .C1(new_n497), .C2(new_n298), .ZN(new_n510));
  OR2_X1    g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OR2_X1    g0311(.A1(new_n484), .A2(G179), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n484), .A2(new_n402), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n512), .A2(new_n464), .A3(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n490), .A2(new_n507), .A3(new_n511), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(KEYINPUT74), .ZN(new_n516));
  INV_X1    g0316(.A(new_n514), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n517), .B1(new_n486), .B2(new_n489), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT74), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n518), .A2(new_n519), .A3(new_n507), .A4(new_n511), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT16), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n262), .A2(new_n229), .A3(new_n263), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n420), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n347), .A2(KEYINPUT7), .A3(new_n229), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n210), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  XNOR2_X1  g0326(.A(G58), .B(G68), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G20), .ZN(new_n528));
  INV_X1    g0328(.A(G159), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n528), .B1(new_n449), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n522), .B1(new_n526), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(G68), .B1(new_n419), .B2(new_n421), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n430), .A2(G159), .B1(new_n527), .B2(G20), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n532), .A2(KEYINPUT16), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n531), .A2(new_n534), .A3(new_n257), .ZN(new_n535));
  INV_X1    g0335(.A(new_n453), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n536), .A2(new_n304), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n537), .B1(new_n501), .B2(new_n536), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n469), .A2(new_n277), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n209), .A2(G1698), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n540), .B(new_n541), .C1(new_n258), .C2(new_n259), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G87), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n283), .ZN(new_n545));
  INV_X1    g0345(.A(new_n476), .ZN(new_n546));
  NOR3_X1   g0346(.A1(new_n472), .A2(new_n475), .A3(G1), .ZN(new_n547));
  OAI211_X1 g0347(.A(G232), .B(new_n353), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  AND4_X1   g0348(.A1(G179), .A2(new_n545), .A3(new_n548), .A4(new_n480), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n479), .B1(new_n544), .B2(new_n283), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n402), .B1(new_n550), .B2(new_n548), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT78), .ZN(new_n552));
  NOR3_X1   g0352(.A1(new_n549), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n545), .A2(new_n548), .A3(new_n480), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(G169), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n550), .A2(G179), .A3(new_n548), .ZN(new_n556));
  AOI21_X1  g0356(.A(KEYINPUT78), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n539), .B1(new_n553), .B2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT18), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n552), .B1(new_n549), .B2(new_n551), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n555), .A2(KEYINPUT78), .A3(new_n556), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n563), .A2(KEYINPUT18), .A3(new_n539), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n550), .A2(G190), .A3(new_n548), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n554), .A2(G200), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n535), .A2(new_n566), .A3(new_n538), .A4(new_n567), .ZN(new_n568));
  XNOR2_X1  g0368(.A(new_n568), .B(KEYINPUT17), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  OR2_X1    g0370(.A1(new_n570), .A2(KEYINPUT79), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n209), .A2(new_n277), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n492), .A2(G1698), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI22_X1  g0374(.A1(new_n574), .A2(new_n347), .B1(new_n254), .B2(new_n202), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n479), .B1(new_n575), .B2(new_n283), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT13), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n477), .A2(G238), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n577), .B1(new_n576), .B2(new_n578), .ZN(new_n580));
  OAI21_X1  g0380(.A(G169), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(KEYINPUT77), .A2(KEYINPUT14), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n580), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n585), .A2(G179), .A3(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(G169), .B(new_n582), .C1(new_n579), .C2(new_n580), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n584), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n303), .A2(G20), .A3(new_n210), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT12), .ZN(new_n591));
  OR2_X1    g0391(.A1(new_n591), .A2(KEYINPUT75), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(KEYINPUT75), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n590), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT76), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n590), .A2(KEYINPUT76), .A3(new_n592), .A4(new_n593), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n596), .B(new_n597), .C1(KEYINPUT12), .C2(new_n590), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n501), .A2(G68), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n454), .A2(G77), .ZN(new_n601));
  OAI221_X1 g0401(.A(new_n601), .B1(new_n229), .B2(G68), .C1(new_n449), .C2(new_n208), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n257), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(KEYINPUT11), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT11), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n602), .A2(new_n605), .A3(new_n257), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n600), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n589), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n585), .A2(G190), .A3(new_n586), .ZN(new_n610));
  OAI21_X1  g0410(.A(G200), .B1(new_n579), .B2(new_n580), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n607), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n613), .B1(new_n570), .B2(KEYINPUT79), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n521), .A2(new_n571), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(KEYINPUT80), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT80), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n521), .A2(new_n571), .A3(new_n617), .A4(new_n614), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n447), .B1(new_n616), .B2(new_n618), .ZN(G372));
  NAND2_X1  g0419(.A1(new_n616), .A2(new_n618), .ZN(new_n620));
  AND4_X1   g0420(.A1(new_n323), .A2(new_n357), .A3(new_n363), .A4(new_n364), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n398), .A2(new_n405), .A3(new_n403), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n389), .A2(new_n375), .A3(new_n392), .A4(new_n393), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n312), .A2(new_n437), .A3(new_n443), .A4(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n406), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n398), .A2(new_n401), .A3(new_n403), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n623), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(KEYINPUT26), .B1(new_n443), .B2(new_n630), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n441), .A2(new_n442), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT26), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n632), .A2(new_n625), .A3(new_n633), .A4(new_n440), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n631), .A2(new_n634), .A3(new_n622), .ZN(new_n635));
  OR2_X1    g0435(.A1(new_n627), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n620), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n555), .A2(new_n556), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n539), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n559), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n539), .A2(KEYINPUT18), .A3(new_n638), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n612), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n609), .B1(new_n507), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n643), .B1(new_n645), .B2(new_n569), .ZN(new_n646));
  INV_X1    g0446(.A(new_n490), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n514), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n637), .A2(new_n649), .ZN(G369));
  OR3_X1    g0450(.A1(new_n326), .A2(KEYINPUT27), .A3(G20), .ZN(new_n651));
  OAI21_X1  g0451(.A(KEYINPUT27), .B1(new_n326), .B2(G20), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(G213), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(G343), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n344), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g0456(.A(new_n656), .B(KEYINPUT88), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n363), .A2(new_n357), .A3(new_n364), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n365), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(new_n657), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n661), .A2(G330), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n325), .A2(new_n446), .ZN(new_n663));
  INV_X1    g0463(.A(new_n655), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n664), .B1(new_n276), .B2(new_n311), .ZN(new_n665));
  OAI22_X1  g0465(.A1(new_n663), .A2(new_n665), .B1(new_n323), .B2(new_n664), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n621), .B1(new_n663), .B2(new_n323), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n664), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n667), .A2(new_n669), .ZN(G399));
  INV_X1    g0470(.A(new_n224), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(G41), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n377), .A2(G116), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G1), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n234), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n675), .B1(new_n676), .B2(new_n673), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT28), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n415), .A2(new_n291), .A3(new_n416), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n350), .A2(new_n354), .A3(G179), .A4(new_n291), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n680), .A2(new_n390), .A3(new_n391), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n679), .A2(KEYINPUT30), .A3(new_n294), .A4(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT30), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n356), .A2(G179), .A3(new_n399), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n415), .A2(new_n291), .A3(new_n416), .A4(new_n294), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n683), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n417), .A2(new_n314), .A3(new_n297), .A4(new_n355), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n682), .B(new_n686), .C1(new_n399), .C2(new_n687), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n688), .A2(KEYINPUT31), .A3(new_n655), .ZN(new_n689));
  AOI21_X1  g0489(.A(KEYINPUT31), .B1(new_n688), .B2(new_n655), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n689), .A2(new_n690), .A3(KEYINPUT89), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n688), .A2(new_n655), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT31), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT89), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(KEYINPUT90), .B1(new_n691), .B2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT90), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n690), .A2(KEYINPUT89), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n688), .A2(KEYINPUT31), .A3(new_n655), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n694), .A2(new_n700), .ZN(new_n701));
  OAI211_X1 g0501(.A(new_n698), .B(new_n699), .C1(new_n701), .C2(KEYINPUT89), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n325), .A2(new_n446), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n703), .A2(new_n444), .A3(new_n365), .A4(new_n664), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n697), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n705), .A2(G330), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n636), .A2(new_n664), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n707), .A2(KEYINPUT29), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n407), .A2(new_n632), .A3(new_n633), .A4(new_n440), .ZN(new_n709));
  OAI21_X1  g0509(.A(KEYINPUT26), .B1(new_n443), .B2(new_n624), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(new_n622), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT91), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n621), .A2(new_n626), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT91), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n709), .A2(new_n710), .A3(new_n714), .A4(new_n622), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n712), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n664), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(KEYINPUT29), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n708), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n706), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n678), .B1(new_n720), .B2(G1), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT92), .ZN(G364));
  INV_X1    g0522(.A(new_n662), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n302), .A2(G20), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G45), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n673), .A2(G1), .A3(new_n725), .ZN(new_n726));
  OR2_X1    g0526(.A1(new_n661), .A2(G330), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n723), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(G13), .A2(G33), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(G20), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n661), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n228), .B1(G20), .B2(new_n402), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g0535(.A(G355), .B(KEYINPUT93), .Z(new_n736));
  NAND2_X1  g0536(.A1(new_n264), .A2(new_n224), .ZN(new_n737));
  OAI22_X1  g0537(.A1(new_n736), .A2(new_n737), .B1(G116), .B2(new_n224), .ZN(new_n738));
  XOR2_X1   g0538(.A(new_n738), .B(KEYINPUT94), .Z(new_n739));
  NOR2_X1   g0539(.A1(new_n671), .A2(new_n264), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(new_n676), .B2(G45), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n741), .B1(new_n248), .B2(G45), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n735), .B1(new_n739), .B2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n726), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n229), .A2(G179), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n745), .A2(G190), .A3(G200), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n348), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n745), .A2(new_n290), .A3(G200), .ZN(new_n748));
  INV_X1    g0548(.A(G283), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n347), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n298), .A2(G190), .ZN(new_n751));
  OAI21_X1  g0551(.A(G20), .B1(new_n751), .B2(G179), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n281), .ZN(new_n754));
  NAND2_X1  g0554(.A1(G20), .A2(G179), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n756), .A2(KEYINPUT95), .A3(G200), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT95), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n758), .B1(new_n755), .B2(new_n298), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(G190), .ZN(new_n761));
  XNOR2_X1  g0561(.A(KEYINPUT33), .B(G317), .ZN(new_n762));
  AOI211_X1 g0562(.A(new_n750), .B(new_n754), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G190), .A2(G200), .ZN(new_n764));
  AND2_X1   g0564(.A1(new_n745), .A2(new_n764), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n765), .A2(KEYINPUT97), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(KEYINPUT97), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G329), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n756), .A2(new_n764), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G311), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT96), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(new_n760), .B2(new_n290), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n757), .A2(KEYINPUT96), .A3(G190), .A4(new_n759), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G326), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n763), .A2(new_n770), .A3(new_n773), .A4(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n751), .A2(new_n755), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n747), .B(new_n779), .C1(G322), .C2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n761), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n782), .A2(new_n210), .B1(new_n503), .B2(new_n771), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT32), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n768), .A2(new_n529), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n783), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n746), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G87), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n777), .A2(G50), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n786), .A2(new_n264), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n752), .B(KEYINPUT98), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n202), .ZN(new_n792));
  INV_X1    g0592(.A(new_n748), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G107), .ZN(new_n794));
  INV_X1    g0594(.A(new_n780), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n794), .B1(new_n231), .B2(new_n795), .C1(new_n785), .C2(new_n784), .ZN(new_n796));
  NOR3_X1   g0596(.A1(new_n790), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n734), .B1(new_n781), .B2(new_n797), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n733), .A2(new_n743), .A3(new_n744), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n728), .A2(new_n799), .ZN(G396));
  NOR2_X1   g0600(.A1(new_n507), .A2(new_n655), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n505), .A2(new_n655), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(new_n509), .B2(new_n510), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n801), .B1(new_n803), .B2(new_n507), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n707), .A2(new_n805), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n664), .B(new_n804), .C1(new_n627), .C2(new_n635), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n706), .B(new_n808), .Z(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(new_n744), .ZN(new_n810));
  INV_X1    g0610(.A(new_n734), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n777), .A2(G137), .B1(G143), .B2(new_n780), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n812), .B1(new_n450), .B2(new_n782), .C1(new_n529), .C2(new_n771), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT34), .Z(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(G50), .B2(new_n787), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n347), .B1(new_n752), .B2(G58), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n769), .A2(G132), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n793), .A2(G68), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n815), .A2(new_n816), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n347), .B1(new_n771), .B2(new_n327), .C1(new_n748), .C2(new_n214), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n792), .B1(G303), .B2(new_n777), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n203), .B2(new_n746), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n820), .B(new_n822), .C1(G311), .C2(new_n769), .ZN(new_n823));
  INV_X1    g0623(.A(G294), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n823), .B1(new_n749), .B2(new_n782), .C1(new_n824), .C2(new_n795), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n811), .B1(new_n819), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n734), .A2(new_n729), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT99), .Z(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(G77), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n804), .A2(new_n730), .ZN(new_n830));
  NOR4_X1   g0630(.A1(new_n826), .A2(new_n726), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n810), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(G384));
  NOR2_X1   g0633(.A1(new_n689), .A2(new_n690), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n447), .B2(new_n655), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n620), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n608), .A2(new_n655), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n609), .A2(new_n612), .A3(new_n837), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n608), .B(new_n655), .C1(new_n644), .C2(new_n589), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n805), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n653), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n539), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(new_n565), .B2(new_n569), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n558), .A2(new_n568), .A3(new_n842), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT37), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n568), .A2(KEYINPUT37), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n539), .B1(new_n638), .B2(new_n841), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT38), .ZN(new_n851));
  NOR3_X1   g0651(.A1(new_n843), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n842), .ZN(new_n853));
  AOI221_X4 g0653(.A(new_n559), .B1(new_n535), .B2(new_n538), .C1(new_n561), .C2(new_n562), .ZN(new_n854));
  AOI21_X1  g0654(.A(KEYINPUT18), .B1(new_n563), .B2(new_n539), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT17), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n568), .B(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n853), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n844), .A2(new_n845), .B1(new_n847), .B2(new_n848), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT38), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n835), .B(new_n840), .C1(new_n852), .C2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT40), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n838), .A2(new_n839), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n804), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(new_n834), .B2(new_n704), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n859), .A2(KEYINPUT38), .A3(new_n860), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n842), .B1(new_n569), .B2(new_n642), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n851), .B1(new_n850), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n863), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n862), .A2(new_n863), .B1(new_n866), .B2(new_n870), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n836), .B(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(G330), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n648), .B1(new_n719), .B2(new_n620), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n874), .B(KEYINPUT102), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n873), .B(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n864), .ZN(new_n877));
  INV_X1    g0677(.A(new_n801), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n807), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT101), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT101), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n807), .A2(new_n881), .A3(new_n878), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n877), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n852), .B2(new_n861), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n643), .A2(new_n653), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n867), .A2(new_n869), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT39), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n609), .A2(new_n655), .ZN(new_n889));
  INV_X1    g0689(.A(new_n861), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n890), .A2(new_n867), .A3(KEYINPUT39), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n884), .A2(new_n885), .A3(new_n892), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n876), .B(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n305), .B2(new_n724), .ZN(new_n895));
  OAI211_X1 g0695(.A(G116), .B(new_n230), .C1(new_n425), .C2(KEYINPUT35), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n896), .B(KEYINPUT100), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n425), .A2(KEYINPUT35), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n899), .B(KEYINPUT36), .ZN(new_n900));
  OAI21_X1  g0700(.A(G77), .B1(new_n231), .B2(new_n210), .ZN(new_n901));
  OAI22_X1  g0701(.A1(new_n676), .A2(new_n901), .B1(G50), .B2(new_n210), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n902), .A2(G1), .A3(new_n302), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n895), .A2(new_n900), .A3(new_n903), .ZN(G367));
  AND2_X1   g0704(.A1(new_n437), .A2(new_n443), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n440), .A2(new_n655), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n658), .A2(new_n664), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n666), .A2(new_n905), .A3(new_n906), .A4(new_n907), .ZN(new_n908));
  OR2_X1    g0708(.A1(new_n908), .A2(KEYINPUT42), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n905), .A2(new_n906), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n443), .B1(new_n910), .B2(new_n323), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n664), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n908), .A2(KEYINPUT42), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n909), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n664), .B1(new_n389), .B2(new_n393), .ZN(new_n915));
  INV_X1    g0715(.A(new_n622), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n624), .B2(new_n915), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT43), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n914), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n667), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n910), .B1(new_n443), .B2(new_n664), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n920), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n918), .A2(KEYINPUT43), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n920), .A2(new_n924), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n928), .ZN(new_n930));
  OAI22_X1  g0730(.A1(new_n930), .A2(new_n925), .B1(KEYINPUT43), .B2(new_n918), .ZN(new_n931));
  XOR2_X1   g0731(.A(KEYINPUT103), .B(KEYINPUT41), .Z(new_n932));
  XNOR2_X1  g0732(.A(new_n672), .B(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n669), .A2(new_n922), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT45), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT104), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT44), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n937), .B(new_n938), .C1(new_n669), .C2(new_n905), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n938), .B1(new_n669), .B2(new_n905), .ZN(new_n940));
  INV_X1    g0740(.A(new_n905), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n668), .A2(KEYINPUT44), .A3(new_n941), .A4(new_n664), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n940), .A2(KEYINPUT104), .A3(new_n942), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n936), .A2(new_n667), .A3(new_n939), .A4(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n939), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n921), .B1(new_n945), .B2(new_n935), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n662), .B(new_n666), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(new_n907), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n944), .A2(new_n720), .A3(new_n946), .A4(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n933), .B1(new_n949), .B2(new_n720), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n725), .A2(G1), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n929), .B(new_n931), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n264), .B1(new_n795), .B2(new_n450), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n787), .A2(G58), .B1(new_n772), .B2(G50), .ZN(new_n954));
  INV_X1    g0754(.A(G137), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n954), .B1(new_n503), .B2(new_n748), .C1(new_n768), .C2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n791), .ZN(new_n957));
  AOI211_X1 g0757(.A(new_n953), .B(new_n956), .C1(G68), .C2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(G143), .ZN(new_n959));
  INV_X1    g0759(.A(new_n777), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n958), .B1(new_n959), .B2(new_n960), .C1(new_n529), .C2(new_n782), .ZN(new_n961));
  INV_X1    g0761(.A(G311), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n793), .A2(G97), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n769), .A2(G317), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n746), .A2(new_n327), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n966), .A2(KEYINPUT46), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n966), .A2(KEYINPUT46), .B1(G303), .B2(new_n780), .ZN(new_n968));
  AND4_X1   g0768(.A1(new_n964), .A2(new_n965), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n752), .A2(G107), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n264), .B1(new_n772), .B2(G283), .ZN(new_n971));
  INV_X1    g0771(.A(new_n281), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n761), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n969), .A2(new_n970), .A3(new_n971), .A4(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n961), .B1(new_n963), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT47), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n734), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n918), .A2(new_n732), .ZN(new_n978));
  INV_X1    g0778(.A(new_n740), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n735), .B1(new_n224), .B2(new_n388), .C1(new_n239), .C2(new_n979), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n977), .A2(new_n744), .A3(new_n978), .A4(new_n980), .ZN(new_n981));
  AND3_X1   g0781(.A1(new_n952), .A2(KEYINPUT105), .A3(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(KEYINPUT105), .B1(new_n952), .B2(new_n981), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n985), .ZN(G387));
  NOR2_X1   g0786(.A1(new_n948), .A2(new_n720), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT114), .Z(new_n988));
  NAND2_X1  g0788(.A1(new_n948), .A2(new_n720), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n672), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(KEYINPUT113), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n990), .A2(KEYINPUT113), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n988), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n674), .B(new_n285), .C1(new_n210), .C2(new_n503), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT107), .Z(new_n995));
  NAND2_X1  g0795(.A1(new_n536), .A2(new_n208), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT50), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n740), .B1(new_n243), .B2(new_n285), .C1(new_n995), .C2(new_n997), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n998), .B1(G107), .B2(new_n224), .C1(new_n674), .C2(new_n737), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n726), .B1(new_n999), .B2(new_n735), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT108), .Z(new_n1001));
  AOI21_X1  g0801(.A(new_n347), .B1(new_n787), .B2(G77), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n1002), .B(new_n964), .C1(new_n768), .C2(new_n450), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT109), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n957), .A2(new_n387), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n780), .A2(G50), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n777), .A2(G159), .B1(new_n536), .B2(new_n761), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(G68), .B2(new_n772), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n777), .A2(G322), .B1(G317), .B2(new_n780), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1010), .B1(new_n348), .B2(new_n771), .C1(new_n962), .C2(new_n782), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT48), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT110), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n972), .A2(new_n787), .B1(G283), .B2(new_n752), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1013), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT111), .Z(new_n1018));
  NAND2_X1  g0818(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g0820(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n1021));
  XNOR2_X1  g0821(.A(new_n1020), .B(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n347), .B1(new_n748), .B2(new_n327), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(new_n769), .B2(G326), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1009), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1001), .B1(new_n666), .B2(new_n732), .C1(new_n1025), .C2(new_n811), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n948), .A2(new_n951), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT106), .Z(new_n1028));
  NAND3_X1  g0828(.A1(new_n993), .A2(new_n1026), .A3(new_n1028), .ZN(G393));
  NAND2_X1  g0829(.A1(new_n944), .A2(new_n946), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n989), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1031), .A2(new_n672), .A3(new_n949), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n944), .A2(new_n951), .A3(new_n946), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n768), .A2(new_n959), .B1(new_n210), .B2(new_n746), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT115), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n208), .B2(new_n782), .C1(new_n214), .C2(new_n748), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n777), .A2(G150), .B1(G159), .B2(new_n780), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT51), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n957), .A2(G77), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n453), .B2(new_n771), .ZN(new_n1040));
  NOR4_X1   g0840(.A1(new_n1036), .A2(new_n1038), .A3(new_n347), .A4(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT116), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n777), .A2(G317), .B1(G311), .B2(new_n780), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT52), .Z(new_n1044));
  NAND2_X1  g0844(.A1(new_n772), .A2(G294), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n769), .A2(G322), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1044), .A2(new_n347), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n746), .A2(new_n749), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n753), .A2(new_n327), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n794), .B1(new_n782), .B2(new_n348), .ZN(new_n1050));
  NOR4_X1   g0850(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n734), .B1(new_n1042), .B2(new_n1051), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n922), .A2(new_n732), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n735), .B1(new_n202), .B2(new_n224), .C1(new_n251), .C2(new_n979), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1052), .A2(new_n1053), .A3(new_n744), .A4(new_n1054), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1032), .A2(new_n1033), .A3(new_n1055), .ZN(G390));
  AND3_X1   g0856(.A1(new_n807), .A2(new_n881), .A3(new_n878), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n881), .B1(new_n807), .B2(new_n878), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n864), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n889), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n1059), .A2(new_n1060), .B1(new_n888), .B2(new_n891), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n803), .A2(new_n507), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n716), .A2(new_n664), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n877), .B1(new_n1063), .B2(new_n878), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n886), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n889), .B(KEYINPUT117), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  NOR3_X1   g0867(.A1(new_n1064), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n705), .A2(G330), .A3(new_n804), .A4(new_n864), .ZN(new_n1069));
  NOR3_X1   g0869(.A1(new_n1061), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  AND3_X1   g0870(.A1(new_n835), .A2(G330), .A3(new_n840), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n891), .A2(new_n888), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n883), .B2(new_n889), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n1063), .A2(new_n878), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n886), .B(new_n1066), .C1(new_n1074), .C2(new_n877), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1071), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1070), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n835), .A2(G330), .A3(new_n804), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n877), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1069), .A2(new_n1074), .A3(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n705), .A2(G330), .A3(new_n804), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1071), .B1(new_n1082), .B2(new_n877), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1081), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n719), .A2(new_n620), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n620), .A2(G330), .A3(new_n835), .ZN(new_n1087));
  AND3_X1   g0887(.A1(new_n1086), .A2(new_n1087), .A3(new_n649), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1078), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1077), .A2(new_n1089), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1091), .A2(new_n672), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1078), .A2(new_n951), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1072), .A2(new_n729), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n828), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n453), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n960), .A2(new_n749), .B1(new_n202), .B2(new_n771), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(G107), .B2(new_n761), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(KEYINPUT118), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n347), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n818), .B1(new_n1099), .B2(KEYINPUT118), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1039), .B1(new_n824), .B2(new_n768), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n788), .B1(new_n327), .B2(new_n795), .ZN(new_n1104));
  NOR4_X1   g0904(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n769), .A2(G125), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n761), .A2(G137), .ZN(new_n1107));
  OR3_X1    g0907(.A1(new_n746), .A2(KEYINPUT53), .A3(new_n450), .ZN(new_n1108));
  OAI21_X1  g0908(.A(KEYINPUT53), .B1(new_n746), .B2(new_n450), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(G128), .B2(new_n777), .ZN(new_n1111));
  XOR2_X1   g0911(.A(KEYINPUT54), .B(G143), .Z(new_n1112));
  NAND2_X1  g0912(.A1(new_n772), .A2(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n957), .A2(G159), .B1(G50), .B2(new_n793), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1111), .A2(new_n264), .A3(new_n1113), .A4(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(G132), .B2(new_n780), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n734), .B1(new_n1105), .B2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1095), .A2(new_n744), .A3(new_n1097), .A4(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1093), .A2(new_n1094), .A3(new_n1118), .ZN(G378));
  INV_X1    g0919(.A(new_n893), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n852), .A2(new_n861), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n447), .A2(new_n655), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n840), .B1(new_n1122), .B2(new_n701), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n863), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT120), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n886), .A2(KEYINPUT40), .A3(new_n835), .A4(new_n840), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1124), .A2(new_n1125), .A3(G330), .A4(new_n1126), .ZN(new_n1127));
  XOR2_X1   g0927(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1128));
  XNOR2_X1  g0928(.A(new_n518), .B(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n464), .A2(new_n841), .ZN(new_n1130));
  XOR2_X1   g0930(.A(new_n1129), .B(new_n1130), .Z(new_n1131));
  NAND2_X1  g0931(.A1(new_n1127), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1125), .B1(new_n871), .B2(G330), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n1125), .B(new_n1131), .C1(new_n871), .C2(G330), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1120), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1124), .A2(G330), .A3(new_n1126), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(KEYINPUT120), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1138), .A2(new_n1127), .A3(new_n1131), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1139), .A2(new_n1140), .A3(new_n893), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1136), .A2(KEYINPUT121), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT121), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1143), .B(new_n1120), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1142), .A2(new_n951), .A3(new_n1144), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n782), .A2(new_n202), .B1(new_n791), .B2(new_n210), .ZN(new_n1146));
  AOI211_X1 g0946(.A(G41), .B(new_n264), .C1(new_n769), .C2(G283), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n1147), .B1(new_n231), .B2(new_n748), .C1(new_n503), .C2(new_n746), .ZN(new_n1148));
  XOR2_X1   g0948(.A(new_n1148), .B(KEYINPUT119), .Z(new_n1149));
  AOI211_X1 g0949(.A(new_n1146), .B(new_n1149), .C1(new_n387), .C2(new_n772), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1150), .B1(new_n203), .B2(new_n795), .C1(new_n327), .C2(new_n960), .ZN(new_n1151));
  XOR2_X1   g0951(.A(new_n1151), .B(KEYINPUT58), .Z(new_n1152));
  OAI21_X1  g0952(.A(new_n208), .B1(new_n258), .B2(G41), .ZN(new_n1153));
  AND2_X1   g0953(.A1(new_n761), .A2(G132), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n787), .A2(new_n1112), .B1(G128), .B2(new_n780), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n1155), .B1(new_n955), .B2(new_n771), .C1(new_n791), .C2(new_n450), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n1154), .B(new_n1156), .C1(G125), .C2(new_n777), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT59), .ZN(new_n1158));
  AOI21_X1  g0958(.A(G33), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(G41), .B1(new_n769), .B2(G124), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1159), .B(new_n1160), .C1(new_n529), .C2(new_n748), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1153), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n734), .B1(new_n1152), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1096), .A2(new_n208), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1131), .A2(new_n729), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1164), .A2(new_n744), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n1145), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1085), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1088), .B1(new_n1077), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1142), .A2(new_n1170), .A3(new_n1144), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT57), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1136), .A2(KEYINPUT122), .A3(new_n1141), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT122), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1139), .A2(new_n1140), .A3(new_n1175), .A4(new_n893), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1174), .A2(new_n1170), .A3(KEYINPUT57), .A4(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n672), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1168), .B1(new_n1173), .B2(new_n1178), .ZN(G375));
  NAND2_X1  g0979(.A1(new_n777), .A2(G132), .ZN(new_n1180));
  XOR2_X1   g0980(.A(new_n1180), .B(KEYINPUT124), .Z(new_n1181));
  AOI22_X1  g0981(.A1(new_n761), .A2(new_n1112), .B1(G137), .B2(new_n780), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT125), .Z(new_n1184));
  NAND2_X1  g0984(.A1(new_n769), .A2(G128), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1184), .A2(new_n264), .A3(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n771), .A2(new_n450), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n791), .A2(new_n208), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n748), .A2(new_n231), .B1(new_n746), .B2(new_n529), .ZN(new_n1189));
  NOR4_X1   g0989(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n769), .A2(G303), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n793), .A2(G77), .B1(new_n772), .B2(G107), .ZN(new_n1192));
  AND3_X1   g0992(.A1(new_n1191), .A2(new_n1005), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n780), .A2(G283), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n264), .B1(new_n761), .B2(G116), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n777), .A2(G294), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .A4(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G97), .B2(new_n787), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n734), .B1(new_n1190), .B2(new_n1198), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1199), .B(new_n744), .C1(new_n730), .C2(new_n864), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n210), .B2(new_n1096), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n951), .B2(new_n1085), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n933), .B(KEYINPUT123), .Z(new_n1204));
  NAND2_X1  g1004(.A1(new_n1089), .A2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1202), .B1(new_n1203), .B2(new_n1205), .ZN(G381));
  NOR3_X1   g1006(.A1(new_n982), .A2(new_n984), .A3(G390), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(G396), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n993), .A2(new_n1209), .A3(new_n1026), .A4(new_n1028), .ZN(new_n1210));
  NOR4_X1   g1010(.A1(new_n1208), .A2(G384), .A3(G381), .A4(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(G375), .A2(G378), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(G407));
  OAI21_X1  g1013(.A(new_n1212), .B1(new_n1211), .B2(new_n654), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(G213), .ZN(G409));
  NAND2_X1  g1015(.A1(G393), .A2(G396), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n1210), .ZN(new_n1217));
  INV_X1    g1017(.A(G390), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n952), .B2(new_n981), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1217), .B1(new_n1207), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1219), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1218), .A2(new_n952), .A3(new_n981), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1221), .A2(new_n1210), .A3(new_n1216), .A4(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1220), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  OAI211_X1 g1025(.A(G378), .B(new_n1168), .C1(new_n1173), .C2(new_n1178), .ZN(new_n1226));
  INV_X1    g1026(.A(G378), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1174), .A2(new_n951), .A3(new_n1176), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1204), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1167), .B(new_n1228), .C1(new_n1171), .C2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1227), .A2(new_n1230), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1226), .A2(KEYINPUT126), .A3(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(KEYINPUT126), .B1(new_n1226), .B2(new_n1231), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n654), .A2(G213), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NOR3_X1   g1035(.A1(new_n1232), .A2(new_n1233), .A3(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1203), .A2(KEYINPUT60), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1237), .A2(new_n672), .A3(new_n1089), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1203), .A2(KEYINPUT60), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1202), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n832), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1240), .A2(new_n832), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1236), .A2(new_n1244), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1245), .A2(KEYINPUT62), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1226), .A2(new_n1231), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1234), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1244), .ZN(new_n1249));
  OAI21_X1  g1049(.A(KEYINPUT62), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(G2897), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1234), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1244), .A2(new_n1252), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n1242), .A2(new_n1243), .B1(new_n1251), .B2(new_n1234), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1248), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT61), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1250), .A2(new_n1256), .A3(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1225), .B1(new_n1246), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1255), .ZN(new_n1260));
  OAI21_X1  g1060(.A(KEYINPUT63), .B1(new_n1236), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1245), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1247), .A2(KEYINPUT63), .A3(new_n1244), .A4(new_n1234), .ZN(new_n1263));
  AND3_X1   g1063(.A1(new_n1224), .A2(new_n1263), .A3(new_n1257), .ZN(new_n1264));
  AOI21_X1  g1064(.A(KEYINPUT127), .B1(new_n1262), .B2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT63), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT126), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1247), .A2(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1226), .A2(KEYINPUT126), .A3(new_n1231), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1268), .A2(new_n1234), .A3(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1266), .B1(new_n1270), .B2(new_n1255), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1270), .A2(new_n1249), .ZN(new_n1272));
  OAI211_X1 g1072(.A(KEYINPUT127), .B(new_n1264), .C1(new_n1271), .C2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1259), .B1(new_n1265), .B2(new_n1274), .ZN(G405));
  NAND2_X1  g1075(.A1(G375), .A2(new_n1227), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1226), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(new_n1277), .B(new_n1244), .ZN(new_n1278));
  XNOR2_X1  g1078(.A(new_n1278), .B(new_n1225), .ZN(G402));
endmodule


