

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590;

  NOR2_X1 U324 ( .A1(n547), .A2(n473), .ZN(n575) );
  NOR2_X1 U325 ( .A1(n557), .A2(n486), .ZN(n405) );
  XNOR2_X1 U326 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U327 ( .A(n438), .B(n318), .ZN(n322) );
  XNOR2_X1 U328 ( .A(n469), .B(n468), .ZN(n546) );
  XNOR2_X1 U329 ( .A(n450), .B(n449), .ZN(n501) );
  XOR2_X1 U330 ( .A(KEYINPUT21), .B(G211GAT), .Z(n292) );
  XNOR2_X1 U331 ( .A(n430), .B(n429), .ZN(n454) );
  XNOR2_X1 U332 ( .A(KEYINPUT45), .B(KEYINPUT66), .ZN(n461) );
  XNOR2_X1 U333 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U334 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U335 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U336 ( .A(n413), .B(n381), .ZN(n382) );
  XNOR2_X1 U337 ( .A(n317), .B(G134GAT), .ZN(n318) );
  XNOR2_X1 U338 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U339 ( .A(n470), .B(KEYINPUT118), .ZN(n471) );
  INV_X1 U340 ( .A(KEYINPUT27), .ZN(n395) );
  XNOR2_X1 U341 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n468) );
  XNOR2_X1 U342 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U343 ( .A(n520), .B(n395), .ZN(n401) );
  XOR2_X1 U344 ( .A(KEYINPUT36), .B(n542), .Z(n586) );
  NAND2_X1 U345 ( .A1(n401), .A2(n574), .ZN(n549) );
  XNOR2_X1 U346 ( .A(KEYINPUT37), .B(n406), .ZN(n516) );
  XOR2_X1 U347 ( .A(n329), .B(n328), .Z(n542) );
  XOR2_X1 U348 ( .A(n392), .B(n391), .Z(n507) );
  XNOR2_X1 U349 ( .A(n478), .B(G190GAT), .ZN(n479) );
  XNOR2_X1 U350 ( .A(n451), .B(G29GAT), .ZN(n452) );
  XNOR2_X1 U351 ( .A(n480), .B(n479), .ZN(G1351GAT) );
  XNOR2_X1 U352 ( .A(n453), .B(n452), .ZN(G1328GAT) );
  XOR2_X1 U353 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n294) );
  XNOR2_X1 U354 ( .A(KEYINPUT91), .B(KEYINPUT6), .ZN(n293) );
  XNOR2_X1 U355 ( .A(n294), .B(n293), .ZN(n312) );
  XOR2_X1 U356 ( .A(G148GAT), .B(G85GAT), .Z(n296) );
  XNOR2_X1 U357 ( .A(G29GAT), .B(G162GAT), .ZN(n295) );
  XNOR2_X1 U358 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U359 ( .A(G155GAT), .B(G57GAT), .Z(n298) );
  XNOR2_X1 U360 ( .A(G120GAT), .B(G127GAT), .ZN(n297) );
  XNOR2_X1 U361 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U362 ( .A(n300), .B(n299), .Z(n305) );
  XOR2_X1 U363 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n302) );
  NAND2_X1 U364 ( .A1(G225GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U365 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U366 ( .A(KEYINPUT1), .B(n303), .ZN(n304) );
  XNOR2_X1 U367 ( .A(n305), .B(n304), .ZN(n308) );
  XOR2_X1 U368 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n307) );
  XNOR2_X1 U369 ( .A(G141GAT), .B(KEYINPUT88), .ZN(n306) );
  XNOR2_X1 U370 ( .A(n307), .B(n306), .ZN(n355) );
  XOR2_X1 U371 ( .A(n308), .B(n355), .Z(n310) );
  XOR2_X1 U372 ( .A(G113GAT), .B(G1GAT), .Z(n434) );
  XOR2_X1 U373 ( .A(G134GAT), .B(KEYINPUT0), .Z(n376) );
  XNOR2_X1 U374 ( .A(n434), .B(n376), .ZN(n309) );
  XNOR2_X1 U375 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U376 ( .A(n312), .B(n311), .ZN(n517) );
  INV_X1 U377 ( .A(n517), .ZN(n547) );
  XOR2_X1 U378 ( .A(KEYINPUT79), .B(KEYINPUT67), .Z(n314) );
  XNOR2_X1 U379 ( .A(KEYINPUT9), .B(G92GAT), .ZN(n313) );
  XNOR2_X1 U380 ( .A(n314), .B(n313), .ZN(n329) );
  XOR2_X1 U381 ( .A(G29GAT), .B(G43GAT), .Z(n316) );
  XNOR2_X1 U382 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n315) );
  XNOR2_X1 U383 ( .A(n316), .B(n315), .ZN(n438) );
  AND2_X1 U384 ( .A1(G232GAT), .A2(G233GAT), .ZN(n317) );
  XOR2_X1 U385 ( .A(KEYINPUT78), .B(G106GAT), .Z(n320) );
  XNOR2_X1 U386 ( .A(KEYINPUT11), .B(KEYINPUT65), .ZN(n319) );
  XNOR2_X1 U387 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U388 ( .A(n322), .B(n321), .ZN(n327) );
  XOR2_X1 U389 ( .A(KEYINPUT10), .B(G218GAT), .Z(n324) );
  XOR2_X1 U390 ( .A(G36GAT), .B(G190GAT), .Z(n385) );
  XOR2_X1 U391 ( .A(G99GAT), .B(G85GAT), .Z(n414) );
  XNOR2_X1 U392 ( .A(n385), .B(n414), .ZN(n323) );
  XNOR2_X1 U393 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U394 ( .A(G50GAT), .B(G162GAT), .Z(n358) );
  XOR2_X1 U395 ( .A(n325), .B(n358), .Z(n326) );
  XNOR2_X1 U396 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U397 ( .A(KEYINPUT84), .B(KEYINPUT15), .Z(n331) );
  XNOR2_X1 U398 ( .A(G211GAT), .B(KEYINPUT82), .ZN(n330) );
  XNOR2_X1 U399 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U400 ( .A(KEYINPUT83), .B(KEYINPUT12), .Z(n333) );
  XNOR2_X1 U401 ( .A(KEYINPUT81), .B(KEYINPUT14), .ZN(n332) );
  XNOR2_X1 U402 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U403 ( .A(n335), .B(n334), .ZN(n346) );
  XOR2_X1 U404 ( .A(G22GAT), .B(G155GAT), .Z(n357) );
  XOR2_X1 U405 ( .A(n357), .B(G78GAT), .Z(n337) );
  XOR2_X1 U406 ( .A(G15GAT), .B(G127GAT), .Z(n363) );
  XNOR2_X1 U407 ( .A(G71GAT), .B(n363), .ZN(n336) );
  XNOR2_X1 U408 ( .A(n337), .B(n336), .ZN(n342) );
  XNOR2_X1 U409 ( .A(G8GAT), .B(G183GAT), .ZN(n338) );
  XOR2_X1 U410 ( .A(n338), .B(KEYINPUT80), .Z(n390) );
  XOR2_X1 U411 ( .A(KEYINPUT13), .B(G57GAT), .Z(n409) );
  XNOR2_X1 U412 ( .A(n390), .B(n409), .ZN(n340) );
  NAND2_X1 U413 ( .A1(G231GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U414 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U415 ( .A(n342), .B(n341), .Z(n344) );
  XNOR2_X1 U416 ( .A(G1GAT), .B(G64GAT), .ZN(n343) );
  XNOR2_X1 U417 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U418 ( .A(n346), .B(n345), .Z(n557) );
  XNOR2_X1 U419 ( .A(G218GAT), .B(G204GAT), .ZN(n347) );
  XNOR2_X1 U420 ( .A(n292), .B(n347), .ZN(n348) );
  XOR2_X1 U421 ( .A(G197GAT), .B(n348), .Z(n383) );
  XOR2_X1 U422 ( .A(KEYINPUT90), .B(KEYINPUT23), .Z(n350) );
  XNOR2_X1 U423 ( .A(KEYINPUT24), .B(KEYINPUT22), .ZN(n349) );
  XNOR2_X1 U424 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U425 ( .A(n383), .B(n351), .ZN(n362) );
  XNOR2_X1 U426 ( .A(G106GAT), .B(G78GAT), .ZN(n352) );
  XNOR2_X1 U427 ( .A(n352), .B(G148GAT), .ZN(n423) );
  XOR2_X1 U428 ( .A(n423), .B(KEYINPUT89), .Z(n354) );
  NAND2_X1 U429 ( .A1(G228GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U430 ( .A(n354), .B(n353), .ZN(n356) );
  XOR2_X1 U431 ( .A(n356), .B(n355), .Z(n360) );
  XNOR2_X1 U432 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U433 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U434 ( .A(n362), .B(n361), .ZN(n474) );
  XOR2_X1 U435 ( .A(G120GAT), .B(G71GAT), .Z(n418) );
  XNOR2_X1 U436 ( .A(n418), .B(n363), .ZN(n366) );
  XOR2_X1 U437 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n365) );
  XNOR2_X1 U438 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n364) );
  XNOR2_X1 U439 ( .A(n365), .B(n364), .ZN(n389) );
  XNOR2_X1 U440 ( .A(n366), .B(n389), .ZN(n370) );
  XOR2_X1 U441 ( .A(KEYINPUT20), .B(KEYINPUT86), .Z(n368) );
  NAND2_X1 U442 ( .A1(G227GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U443 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U444 ( .A(n370), .B(n369), .Z(n375) );
  XOR2_X1 U445 ( .A(G183GAT), .B(G176GAT), .Z(n372) );
  XNOR2_X1 U446 ( .A(G113GAT), .B(G99GAT), .ZN(n371) );
  XNOR2_X1 U447 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U448 ( .A(n373), .B(KEYINPUT87), .ZN(n374) );
  XNOR2_X1 U449 ( .A(n375), .B(n374), .ZN(n377) );
  XOR2_X1 U450 ( .A(n377), .B(n376), .Z(n379) );
  XNOR2_X1 U451 ( .A(G43GAT), .B(G190GAT), .ZN(n378) );
  XOR2_X1 U452 ( .A(n379), .B(n378), .Z(n524) );
  INV_X1 U453 ( .A(n524), .ZN(n532) );
  XNOR2_X1 U454 ( .A(G176GAT), .B(G92GAT), .ZN(n380) );
  XNOR2_X1 U455 ( .A(n380), .B(G64GAT), .ZN(n413) );
  XOR2_X1 U456 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n381) );
  XOR2_X1 U457 ( .A(n385), .B(n384), .Z(n387) );
  NAND2_X1 U458 ( .A1(G226GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U459 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U460 ( .A(n389), .B(n388), .ZN(n392) );
  INV_X1 U461 ( .A(n390), .ZN(n391) );
  NAND2_X1 U462 ( .A1(n532), .A2(n507), .ZN(n393) );
  NAND2_X1 U463 ( .A1(n474), .A2(n393), .ZN(n394) );
  XOR2_X1 U464 ( .A(KEYINPUT25), .B(n394), .Z(n398) );
  INV_X1 U465 ( .A(n507), .ZN(n520) );
  XNOR2_X1 U466 ( .A(KEYINPUT26), .B(KEYINPUT96), .ZN(n397) );
  NOR2_X1 U467 ( .A1(n532), .A2(n474), .ZN(n396) );
  XNOR2_X1 U468 ( .A(n397), .B(n396), .ZN(n574) );
  NAND2_X1 U469 ( .A1(n398), .A2(n549), .ZN(n399) );
  XNOR2_X1 U470 ( .A(KEYINPUT97), .B(n399), .ZN(n400) );
  NOR2_X1 U471 ( .A1(n547), .A2(n400), .ZN(n404) );
  XNOR2_X1 U472 ( .A(n474), .B(KEYINPUT28), .ZN(n529) );
  AND2_X1 U473 ( .A1(n529), .A2(n401), .ZN(n402) );
  NAND2_X1 U474 ( .A1(n547), .A2(n402), .ZN(n534) );
  NOR2_X1 U475 ( .A1(n532), .A2(n534), .ZN(n403) );
  NOR2_X1 U476 ( .A1(n404), .A2(n403), .ZN(n486) );
  NAND2_X1 U477 ( .A1(n586), .A2(n405), .ZN(n406) );
  XOR2_X1 U478 ( .A(KEYINPUT73), .B(KEYINPUT72), .Z(n408) );
  XNOR2_X1 U479 ( .A(KEYINPUT76), .B(KEYINPUT33), .ZN(n407) );
  XNOR2_X1 U480 ( .A(n408), .B(n407), .ZN(n410) );
  XNOR2_X1 U481 ( .A(n410), .B(n409), .ZN(n422) );
  INV_X1 U482 ( .A(n413), .ZN(n412) );
  INV_X1 U483 ( .A(n414), .ZN(n411) );
  NAND2_X1 U484 ( .A1(n412), .A2(n411), .ZN(n416) );
  NAND2_X1 U485 ( .A1(n414), .A2(n413), .ZN(n415) );
  NAND2_X1 U486 ( .A1(n416), .A2(n415), .ZN(n420) );
  AND2_X1 U487 ( .A1(G230GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U488 ( .A(n422), .B(n421), .ZN(n424) );
  XNOR2_X1 U489 ( .A(n424), .B(n423), .ZN(n430) );
  XOR2_X1 U490 ( .A(G204GAT), .B(KEYINPUT75), .Z(n426) );
  XNOR2_X1 U491 ( .A(KEYINPUT31), .B(KEYINPUT32), .ZN(n425) );
  XOR2_X1 U492 ( .A(n426), .B(n425), .Z(n428) );
  XNOR2_X1 U493 ( .A(KEYINPUT77), .B(KEYINPUT74), .ZN(n427) );
  XOR2_X1 U494 ( .A(G8GAT), .B(KEYINPUT69), .Z(n432) );
  XNOR2_X1 U495 ( .A(G50GAT), .B(G36GAT), .ZN(n431) );
  XNOR2_X1 U496 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U497 ( .A(n434), .B(n433), .Z(n436) );
  NAND2_X1 U498 ( .A1(G229GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U499 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U500 ( .A(n437), .B(G141GAT), .Z(n440) );
  XNOR2_X1 U501 ( .A(G169GAT), .B(n438), .ZN(n439) );
  XNOR2_X1 U502 ( .A(n440), .B(n439), .ZN(n448) );
  XOR2_X1 U503 ( .A(KEYINPUT71), .B(KEYINPUT68), .Z(n442) );
  XNOR2_X1 U504 ( .A(G22GAT), .B(G15GAT), .ZN(n441) );
  XNOR2_X1 U505 ( .A(n442), .B(n441), .ZN(n446) );
  XOR2_X1 U506 ( .A(G197GAT), .B(KEYINPUT70), .Z(n444) );
  XNOR2_X1 U507 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n443) );
  XNOR2_X1 U508 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U509 ( .A(n446), .B(n445), .Z(n447) );
  XOR2_X1 U510 ( .A(n448), .B(n447), .Z(n550) );
  INV_X1 U511 ( .A(n550), .ZN(n576) );
  NOR2_X1 U512 ( .A1(n454), .A2(n576), .ZN(n487) );
  NAND2_X1 U513 ( .A1(n516), .A2(n487), .ZN(n450) );
  XNOR2_X1 U514 ( .A(KEYINPUT38), .B(KEYINPUT101), .ZN(n449) );
  NAND2_X1 U515 ( .A1(n547), .A2(n501), .ZN(n453) );
  XOR2_X1 U516 ( .A(KEYINPUT102), .B(KEYINPUT39), .Z(n451) );
  XOR2_X1 U517 ( .A(KEYINPUT41), .B(n454), .Z(n552) );
  NAND2_X1 U518 ( .A1(n552), .A2(n550), .ZN(n456) );
  XNOR2_X1 U519 ( .A(KEYINPUT46), .B(KEYINPUT110), .ZN(n455) );
  XNOR2_X1 U520 ( .A(n456), .B(n455), .ZN(n458) );
  INV_X1 U521 ( .A(n557), .ZN(n584) );
  AND2_X1 U522 ( .A1(n542), .A2(n584), .ZN(n457) );
  NAND2_X1 U523 ( .A1(n458), .A2(n457), .ZN(n459) );
  XNOR2_X1 U524 ( .A(n459), .B(KEYINPUT47), .ZN(n460) );
  XNOR2_X1 U525 ( .A(n460), .B(KEYINPUT111), .ZN(n467) );
  NAND2_X1 U526 ( .A1(n557), .A2(n586), .ZN(n462) );
  NOR2_X1 U527 ( .A1(n463), .A2(n454), .ZN(n464) );
  XNOR2_X1 U528 ( .A(n464), .B(KEYINPUT112), .ZN(n465) );
  NAND2_X1 U529 ( .A1(n465), .A2(n576), .ZN(n466) );
  NAND2_X1 U530 ( .A1(n467), .A2(n466), .ZN(n469) );
  NAND2_X1 U531 ( .A1(n507), .A2(n546), .ZN(n472) );
  XOR2_X1 U532 ( .A(KEYINPUT119), .B(KEYINPUT54), .Z(n470) );
  NAND2_X1 U533 ( .A1(n575), .A2(n474), .ZN(n475) );
  XNOR2_X1 U534 ( .A(n475), .B(KEYINPUT120), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n476), .B(KEYINPUT55), .ZN(n477) );
  NAND2_X1 U536 ( .A1(n477), .A2(n532), .ZN(n570) );
  NOR2_X1 U537 ( .A1(n570), .A2(n542), .ZN(n480) );
  INV_X1 U538 ( .A(KEYINPUT58), .ZN(n478) );
  NOR2_X1 U539 ( .A1(n576), .A2(n570), .ZN(n482) );
  XNOR2_X1 U540 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n481) );
  XNOR2_X1 U541 ( .A(n482), .B(n481), .ZN(G1348GAT) );
  XOR2_X1 U542 ( .A(KEYINPUT85), .B(KEYINPUT16), .Z(n484) );
  NAND2_X1 U543 ( .A1(n542), .A2(n557), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n484), .B(n483), .ZN(n485) );
  NOR2_X1 U545 ( .A1(n486), .A2(n485), .ZN(n503) );
  NAND2_X1 U546 ( .A1(n487), .A2(n503), .ZN(n496) );
  NOR2_X1 U547 ( .A1(n517), .A2(n496), .ZN(n489) );
  XNOR2_X1 U548 ( .A(KEYINPUT34), .B(KEYINPUT98), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U550 ( .A(G1GAT), .B(n490), .Z(G1324GAT) );
  NOR2_X1 U551 ( .A1(n520), .A2(n496), .ZN(n491) );
  XOR2_X1 U552 ( .A(G8GAT), .B(n491), .Z(G1325GAT) );
  NOR2_X1 U553 ( .A1(n496), .A2(n524), .ZN(n495) );
  XOR2_X1 U554 ( .A(KEYINPUT99), .B(KEYINPUT35), .Z(n493) );
  XNOR2_X1 U555 ( .A(G15GAT), .B(KEYINPUT100), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n495), .B(n494), .ZN(G1326GAT) );
  NOR2_X1 U558 ( .A1(n529), .A2(n496), .ZN(n497) );
  XOR2_X1 U559 ( .A(G22GAT), .B(n497), .Z(G1327GAT) );
  NAND2_X1 U560 ( .A1(n501), .A2(n507), .ZN(n498) );
  XNOR2_X1 U561 ( .A(n498), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U562 ( .A1(n501), .A2(n532), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n499), .B(KEYINPUT40), .ZN(n500) );
  XNOR2_X1 U564 ( .A(G43GAT), .B(n500), .ZN(G1330GAT) );
  INV_X1 U565 ( .A(n529), .ZN(n511) );
  NAND2_X1 U566 ( .A1(n501), .A2(n511), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n502), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n506) );
  INV_X1 U569 ( .A(n552), .ZN(n564) );
  NOR2_X1 U570 ( .A1(n550), .A2(n564), .ZN(n515) );
  NAND2_X1 U571 ( .A1(n503), .A2(n515), .ZN(n504) );
  XNOR2_X1 U572 ( .A(n504), .B(KEYINPUT103), .ZN(n512) );
  NAND2_X1 U573 ( .A1(n547), .A2(n512), .ZN(n505) );
  XNOR2_X1 U574 ( .A(n506), .B(n505), .ZN(G1332GAT) );
  NAND2_X1 U575 ( .A1(n507), .A2(n512), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n508), .B(KEYINPUT104), .ZN(n509) );
  XNOR2_X1 U577 ( .A(G64GAT), .B(n509), .ZN(G1333GAT) );
  NAND2_X1 U578 ( .A1(n512), .A2(n532), .ZN(n510) );
  XNOR2_X1 U579 ( .A(n510), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U580 ( .A(G78GAT), .B(KEYINPUT43), .Z(n514) );
  NAND2_X1 U581 ( .A1(n512), .A2(n511), .ZN(n513) );
  XNOR2_X1 U582 ( .A(n514), .B(n513), .ZN(G1335GAT) );
  NAND2_X1 U583 ( .A1(n516), .A2(n515), .ZN(n528) );
  NOR2_X1 U584 ( .A1(n517), .A2(n528), .ZN(n519) );
  XNOR2_X1 U585 ( .A(G85GAT), .B(KEYINPUT105), .ZN(n518) );
  XNOR2_X1 U586 ( .A(n519), .B(n518), .ZN(G1336GAT) );
  NOR2_X1 U587 ( .A1(n520), .A2(n528), .ZN(n522) );
  XNOR2_X1 U588 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n521) );
  XNOR2_X1 U589 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U590 ( .A(G92GAT), .B(n523), .ZN(G1337GAT) );
  NOR2_X1 U591 ( .A1(n524), .A2(n528), .ZN(n525) );
  XOR2_X1 U592 ( .A(G99GAT), .B(n525), .Z(G1338GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT108), .B(KEYINPUT44), .Z(n527) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(KEYINPUT109), .ZN(n526) );
  XNOR2_X1 U595 ( .A(n527), .B(n526), .ZN(n531) );
  NOR2_X1 U596 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U597 ( .A(n531), .B(n530), .Z(G1339GAT) );
  NAND2_X1 U598 ( .A1(n532), .A2(n546), .ZN(n533) );
  NOR2_X1 U599 ( .A1(n534), .A2(n533), .ZN(n543) );
  NAND2_X1 U600 ( .A1(n543), .A2(n550), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n535), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT113), .B(KEYINPUT49), .Z(n537) );
  NAND2_X1 U603 ( .A1(n543), .A2(n552), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U605 ( .A(G120GAT), .B(n538), .Z(G1341GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT114), .B(KEYINPUT50), .Z(n540) );
  NAND2_X1 U607 ( .A1(n543), .A2(n557), .ZN(n539) );
  XNOR2_X1 U608 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U609 ( .A(G127GAT), .B(n541), .Z(G1342GAT) );
  XOR2_X1 U610 ( .A(G134GAT), .B(KEYINPUT51), .Z(n545) );
  INV_X1 U611 ( .A(n542), .ZN(n560) );
  NAND2_X1 U612 ( .A1(n543), .A2(n560), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(G1343GAT) );
  NAND2_X1 U614 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U615 ( .A1(n549), .A2(n548), .ZN(n561) );
  NAND2_X1 U616 ( .A1(n561), .A2(n550), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n551), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT115), .B(KEYINPUT53), .Z(n554) );
  NAND2_X1 U619 ( .A1(n561), .A2(n552), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(n556) );
  XOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT52), .Z(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1345GAT) );
  NAND2_X1 U623 ( .A1(n557), .A2(n561), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(KEYINPUT116), .ZN(n559) );
  XNOR2_X1 U625 ( .A(G155GAT), .B(n559), .ZN(G1346GAT) );
  XOR2_X1 U626 ( .A(G162GAT), .B(KEYINPUT117), .Z(n563) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(G1347GAT) );
  NOR2_X1 U629 ( .A1(n564), .A2(n570), .ZN(n569) );
  XOR2_X1 U630 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n566) );
  XNOR2_X1 U631 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(KEYINPUT56), .B(n567), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(G1349GAT) );
  NOR2_X1 U635 ( .A1(n584), .A2(n570), .ZN(n571) );
  XOR2_X1 U636 ( .A(G183GAT), .B(n571), .Z(G1350GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT124), .B(KEYINPUT59), .Z(n573) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n578) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n583) );
  NOR2_X1 U641 ( .A1(n576), .A2(n583), .ZN(n577) );
  XOR2_X1 U642 ( .A(n578), .B(n577), .Z(G1352GAT) );
  INV_X1 U643 ( .A(n583), .ZN(n587) );
  AND2_X1 U644 ( .A1(n587), .A2(n454), .ZN(n582) );
  XOR2_X1 U645 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n580) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n579) );
  XNOR2_X1 U647 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  NOR2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U650 ( .A(G211GAT), .B(n585), .Z(G1354GAT) );
  XOR2_X1 U651 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n589) );
  NAND2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

