//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 1 0 1 0 0 0 1 1 0 0 1 1 1 1 0 0 1 1 0 0 0 1 0 1 1 1 0 0 0 0 1 0 0 0 0 1 0 0 0 0 0 0 0 1 0 1 0 0 1 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n804, new_n805, new_n807,
    new_n808, new_n809, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n873, new_n874, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n923, new_n924;
  XOR2_X1   g000(.A(G211gat), .B(G218gat), .Z(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT76), .ZN(new_n203));
  XNOR2_X1  g002(.A(G197gat), .B(G204gat), .ZN(new_n204));
  INV_X1    g003(.A(G211gat), .ZN(new_n205));
  INV_X1    g004(.A(G218gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI211_X1 g006(.A(new_n203), .B(new_n204), .C1(KEYINPUT22), .C2(new_n207), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n202), .A2(KEYINPUT76), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT29), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n208), .A2(new_n209), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT3), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216));
  INV_X1    g015(.A(G155gat), .ZN(new_n217));
  INV_X1    g016(.A(G162gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G141gat), .B(G148gat), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n216), .B(new_n219), .C1(new_n220), .C2(KEYINPUT2), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n221), .B(KEYINPUT81), .ZN(new_n222));
  INV_X1    g021(.A(G148gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(G141gat), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT82), .B(G141gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n224), .B1(new_n225), .B2(new_n223), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n216), .B1(new_n219), .B2(KEYINPUT2), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n222), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n215), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n210), .A2(new_n212), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n229), .A2(KEYINPUT3), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n231), .B1(new_n232), .B2(KEYINPUT29), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT85), .B1(new_n230), .B2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n234), .A2(G228gat), .A3(G233gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n230), .A2(new_n233), .A3(KEYINPUT85), .ZN(new_n236));
  INV_X1    g035(.A(G228gat), .ZN(new_n237));
  INV_X1    g036(.A(G233gat), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n235), .B1(new_n239), .B2(new_n234), .ZN(new_n240));
  XNOR2_X1  g039(.A(G78gat), .B(G106gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT31), .B(G50gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n241), .B(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n240), .A2(new_n244), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n235), .B(new_n243), .C1(new_n239), .C2(new_n234), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT86), .ZN(new_n247));
  INV_X1    g046(.A(G22gat), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n248), .B1(new_n246), .B2(new_n247), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n245), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n246), .A2(new_n247), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(G22gat), .ZN(new_n253));
  INV_X1    g052(.A(new_n245), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n253), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  AND2_X1   g055(.A1(new_n251), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G15gat), .B(G43gat), .ZN(new_n258));
  INV_X1    g057(.A(G99gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT71), .B(G71gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT33), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT66), .ZN(new_n265));
  INV_X1    g064(.A(G183gat), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n265), .B1(new_n266), .B2(KEYINPUT27), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT27), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n268), .A2(KEYINPUT66), .A3(G183gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n266), .A2(KEYINPUT27), .ZN(new_n270));
  NOR2_X1   g069(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n267), .A2(new_n269), .A3(new_n270), .A4(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(G183gat), .A2(G190gat), .ZN(new_n273));
  AND2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(G169gat), .A2(G176gat), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT26), .ZN(new_n276));
  OR3_X1    g075(.A1(new_n275), .A2(KEYINPUT68), .A3(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(KEYINPUT68), .B1(new_n275), .B2(new_n276), .ZN(new_n278));
  AND2_X1   g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n279), .B1(new_n276), .B2(new_n275), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n277), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n268), .A2(G183gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n266), .A2(KEYINPUT27), .ZN(new_n283));
  OAI21_X1  g082(.A(KEYINPUT67), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n268), .A2(G183gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT67), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n270), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(G190gat), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT28), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n274), .B(new_n281), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT25), .ZN(new_n291));
  AND3_X1   g090(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n292));
  OAI21_X1  g091(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n292), .B1(new_n273), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(G169gat), .ZN(new_n295));
  INV_X1    g094(.A(G176gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n295), .A2(new_n296), .A3(KEYINPUT23), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT23), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n298), .B1(G169gat), .B2(G176gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(G169gat), .A2(G176gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n297), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n291), .B1(new_n294), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT64), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT24), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n273), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(G190gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n266), .A2(new_n306), .ZN(new_n307));
  OAI211_X1 g106(.A(G183gat), .B(G190gat), .C1(KEYINPUT64), .C2(KEYINPUT24), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n305), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n279), .B1(KEYINPUT23), .B2(new_n275), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n309), .A2(new_n310), .A3(KEYINPUT25), .A4(new_n299), .ZN(new_n311));
  AND3_X1   g110(.A1(new_n302), .A2(new_n311), .A3(KEYINPUT65), .ZN(new_n312));
  AOI21_X1  g111(.A(KEYINPUT65), .B1(new_n302), .B2(new_n311), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n290), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G113gat), .B(G120gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n315), .A2(KEYINPUT1), .ZN(new_n316));
  XOR2_X1   g115(.A(G127gat), .B(G134gat), .Z(new_n317));
  XNOR2_X1  g116(.A(new_n316), .B(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n318), .B(new_n290), .C1(new_n312), .C2(new_n313), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(G227gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n323), .A2(new_n238), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n264), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n324), .ZN(new_n326));
  AOI211_X1 g125(.A(KEYINPUT69), .B(new_n326), .C1(new_n320), .C2(new_n321), .ZN(new_n327));
  OAI211_X1 g126(.A(KEYINPUT32), .B(new_n263), .C1(new_n325), .C2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT73), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT72), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT33), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n332), .B1(new_n325), .B2(new_n327), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT32), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n302), .A2(new_n311), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT65), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n302), .A2(new_n311), .A3(KEYINPUT65), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n318), .B1(new_n339), .B2(new_n290), .ZN(new_n340));
  INV_X1    g139(.A(new_n321), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n324), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT69), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n322), .A2(new_n264), .A3(new_n324), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n334), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT70), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n262), .B(new_n333), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT32), .B1(new_n325), .B2(new_n327), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n348), .A2(KEYINPUT70), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n331), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n333), .A2(new_n262), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n345), .A2(new_n346), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n348), .A2(KEYINPUT70), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n351), .A2(KEYINPUT72), .A3(new_n352), .A4(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n330), .B1(new_n350), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n320), .A2(new_n326), .A3(new_n321), .ZN(new_n356));
  XOR2_X1   g155(.A(new_n356), .B(KEYINPUT34), .Z(new_n357));
  OR2_X1    g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n350), .A2(new_n354), .ZN(new_n359));
  INV_X1    g158(.A(new_n330), .ZN(new_n360));
  AND4_X1   g159(.A1(KEYINPUT74), .A2(new_n359), .A3(new_n357), .A4(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT74), .B1(new_n355), .B2(new_n357), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n257), .B(new_n358), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  AND2_X1   g162(.A1(new_n222), .A2(new_n228), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(new_n318), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n229), .A2(new_n319), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(G225gat), .A2(G233gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(KEYINPUT84), .B(KEYINPUT5), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NOR3_X1   g169(.A1(new_n367), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n365), .B(KEYINPUT4), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n232), .A2(new_n318), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n373), .B1(new_n214), .B2(new_n364), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n372), .A2(new_n368), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n375), .A2(KEYINPUT83), .A3(new_n369), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n369), .A2(KEYINPUT83), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n372), .A2(new_n368), .A3(new_n374), .A4(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n371), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(G1gat), .B(G29gat), .ZN(new_n380));
  INV_X1    g179(.A(G85gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n380), .B(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(KEYINPUT0), .B(G57gat), .ZN(new_n383));
  XOR2_X1   g182(.A(new_n382), .B(new_n383), .Z(new_n384));
  AND2_X1   g183(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT6), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT6), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n387), .B1(new_n379), .B2(new_n384), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n386), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n314), .B(KEYINPUT78), .ZN(new_n390));
  NAND2_X1  g189(.A1(G226gat), .A2(G233gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n391), .B(KEYINPUT77), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  AND2_X1   g192(.A1(new_n290), .A2(new_n335), .ZN(new_n394));
  OR2_X1    g193(.A1(new_n394), .A2(KEYINPUT29), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n390), .A2(new_n393), .B1(new_n391), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n231), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n394), .A2(new_n391), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n390), .A2(new_n211), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n399), .B1(new_n400), .B2(new_n392), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n398), .B1(new_n401), .B2(new_n397), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(G8gat), .B(G36gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(G64gat), .B(G92gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n404), .B(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT80), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OR2_X1    g209(.A1(new_n410), .A2(KEYINPUT30), .ZN(new_n411));
  XOR2_X1   g210(.A(new_n402), .B(KEYINPUT79), .Z(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(new_n406), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n410), .A2(KEYINPUT30), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n389), .A2(new_n411), .A3(new_n413), .A4(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(KEYINPUT35), .B1(new_n363), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT75), .B1(new_n361), .B2(new_n362), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n359), .A2(new_n357), .A3(new_n360), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT74), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT75), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n355), .A2(KEYINPUT74), .A3(new_n357), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n411), .A2(new_n413), .A3(new_n414), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n417), .A2(new_n423), .A3(new_n424), .A4(new_n358), .ZN(new_n425));
  INV_X1    g224(.A(new_n388), .ZN(new_n426));
  XOR2_X1   g225(.A(new_n384), .B(KEYINPUT88), .Z(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n379), .A2(new_n428), .ZN(new_n429));
  AOI22_X1  g228(.A1(new_n426), .A2(new_n429), .B1(new_n385), .B2(KEYINPUT6), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n251), .A2(new_n256), .ZN(new_n431));
  OR3_X1    g230(.A1(new_n430), .A2(new_n431), .A3(KEYINPUT35), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n416), .B1(new_n425), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n257), .A2(KEYINPUT87), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT87), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n415), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT37), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n407), .B1(new_n403), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT38), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n438), .B1(new_n396), .B2(new_n231), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n441), .B1(new_n401), .B2(new_n231), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n439), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n430), .A2(new_n443), .A3(new_n408), .ZN(new_n444));
  AND2_X1   g243(.A1(new_n412), .A2(KEYINPUT37), .ZN(new_n445));
  INV_X1    g244(.A(new_n439), .ZN(new_n446));
  OAI211_X1 g245(.A(KEYINPUT90), .B(KEYINPUT38), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT90), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n446), .B1(new_n412), .B2(KEYINPUT37), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n448), .B1(new_n449), .B2(new_n440), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n444), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n368), .B1(new_n372), .B2(new_n374), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT39), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n428), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n367), .A2(new_n368), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT39), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n454), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT89), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT40), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n460), .B(new_n429), .C1(new_n459), .C2(new_n457), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n458), .B1(new_n457), .B2(new_n459), .ZN(new_n462));
  OR2_X1    g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n257), .B1(new_n424), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n437), .B1(new_n451), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT36), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n355), .A2(new_n357), .ZN(new_n467));
  AOI211_X1 g266(.A(new_n466), .B(new_n467), .C1(new_n420), .C2(new_n422), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n417), .A2(new_n423), .A3(new_n358), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n468), .B1(new_n469), .B2(new_n466), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n433), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(G15gat), .B(G22gat), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT16), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n472), .B1(new_n473), .B2(G1gat), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n474), .B1(G1gat), .B2(new_n472), .ZN(new_n475));
  INV_X1    g274(.A(G8gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n475), .B(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT95), .ZN(new_n479));
  INV_X1    g278(.A(G71gat), .ZN(new_n480));
  INV_X1    g279(.A(G78gat), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OR2_X1    g281(.A1(G57gat), .A2(G64gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(G57gat), .A2(G64gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n482), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(G71gat), .B(G78gat), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n488), .B(new_n482), .C1(new_n485), .C2(new_n486), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n478), .B1(KEYINPUT21), .B2(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n492), .B(KEYINPUT21), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(new_n477), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(G183gat), .B(G211gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n497), .B(KEYINPUT96), .ZN(new_n498));
  NAND2_X1  g297(.A1(G231gat), .A2(G233gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n498), .B(new_n499), .ZN(new_n500));
  OR2_X1    g299(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(G127gat), .B(G155gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n502), .B(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n496), .A2(new_n500), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n501), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n504), .B1(new_n501), .B2(new_n505), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XOR2_X1   g307(.A(G190gat), .B(G218gat), .Z(new_n509));
  OR2_X1    g308(.A1(G99gat), .A2(G106gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(G99gat), .A2(G106gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT100), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT100), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n510), .A2(new_n514), .A3(new_n511), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT98), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT7), .ZN(new_n518));
  NAND2_X1  g317(.A1(G85gat), .A2(G92gat), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n517), .B(new_n518), .C1(new_n519), .C2(KEYINPUT99), .ZN(new_n520));
  INV_X1    g319(.A(G92gat), .ZN(new_n521));
  AOI22_X1  g320(.A1(KEYINPUT8), .A2(new_n511), .B1(new_n381), .B2(new_n521), .ZN(new_n522));
  AND2_X1   g321(.A1(G85gat), .A2(G92gat), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT99), .ZN(new_n524));
  AOI21_X1  g323(.A(KEYINPUT98), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT7), .B1(new_n519), .B2(new_n517), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n520), .B(new_n522), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n516), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n516), .A2(new_n527), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT14), .ZN(new_n531));
  INV_X1    g330(.A(G29gat), .ZN(new_n532));
  INV_X1    g331(.A(G36gat), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n535));
  AOI22_X1  g334(.A1(new_n534), .A2(new_n535), .B1(G29gat), .B2(G36gat), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT15), .ZN(new_n537));
  INV_X1    g336(.A(G50gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(G43gat), .ZN(new_n539));
  INV_X1    g338(.A(G43gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(G50gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT91), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n537), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G43gat), .B(G50gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT91), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n536), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n542), .A2(KEYINPUT92), .A3(new_n537), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT92), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n549), .B1(new_n545), .B2(KEYINPUT15), .ZN(new_n550));
  OAI21_X1  g349(.A(KEYINPUT15), .B1(new_n545), .B2(KEYINPUT91), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n542), .A2(new_n543), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n548), .B(new_n550), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n547), .B1(new_n553), .B2(new_n536), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT93), .ZN(new_n555));
  AOI21_X1  g354(.A(KEYINPUT17), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n554), .A2(new_n555), .A3(KEYINPUT17), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n530), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(G232gat), .A2(G233gat), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  AOI22_X1  g360(.A1(new_n530), .A2(new_n554), .B1(KEYINPUT41), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n509), .B1(new_n559), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n530), .ZN(new_n565));
  INV_X1    g364(.A(new_n558), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n565), .B1(new_n566), .B2(new_n556), .ZN(new_n567));
  INV_X1    g366(.A(new_n509), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n567), .A2(new_n568), .A3(new_n562), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n561), .A2(KEYINPUT41), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT97), .ZN(new_n572));
  XNOR2_X1  g371(.A(G134gat), .B(G162gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n564), .A2(new_n574), .A3(new_n569), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n508), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(G230gat), .A2(G233gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT102), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  OAI211_X1 g381(.A(new_n490), .B(new_n491), .C1(new_n528), .C2(new_n529), .ZN(new_n583));
  OR2_X1    g382(.A1(new_n516), .A2(new_n527), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n516), .A2(new_n527), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n584), .A2(new_n492), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n583), .A2(KEYINPUT101), .A3(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT101), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n530), .A2(new_n588), .A3(new_n492), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT10), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT10), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n586), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n582), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n587), .A2(new_n581), .A3(new_n589), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G120gat), .B(G148gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(G176gat), .B(G204gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n595), .A2(new_n598), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n477), .B1(new_n566), .B2(new_n556), .ZN(new_n604));
  NAND2_X1  g403(.A1(G229gat), .A2(G233gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n478), .A2(new_n554), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT18), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n604), .A2(KEYINPUT18), .A3(new_n605), .A4(new_n606), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n477), .B(new_n554), .ZN(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT94), .B(KEYINPUT13), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(new_n605), .ZN(new_n613));
  OR2_X1    g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n609), .A2(new_n610), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G113gat), .B(G141gat), .ZN(new_n616));
  INV_X1    g415(.A(G197gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(KEYINPUT11), .B(G169gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n615), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n609), .A2(new_n610), .A3(new_n614), .A4(new_n621), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AND4_X1   g424(.A1(new_n471), .A2(new_n579), .A3(new_n603), .A4(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n389), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(KEYINPUT103), .B(G1gat), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(G1324gat));
  INV_X1    g429(.A(new_n424), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n626), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(KEYINPUT42), .B1(new_n632), .B2(new_n476), .ZN(new_n633));
  NAND2_X1  g432(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n473), .A2(new_n476), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n632), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  MUX2_X1   g435(.A(KEYINPUT42), .B(new_n633), .S(new_n636), .Z(G1325gat));
  INV_X1    g436(.A(new_n469), .ZN(new_n638));
  AOI21_X1  g437(.A(G15gat), .B1(new_n626), .B2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n361), .A2(new_n362), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n467), .B1(new_n640), .B2(new_n421), .ZN(new_n641));
  AOI21_X1  g440(.A(KEYINPUT36), .B1(new_n641), .B2(new_n417), .ZN(new_n642));
  OAI21_X1  g441(.A(KEYINPUT104), .B1(new_n642), .B2(new_n468), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT104), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n470), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n646), .A2(G15gat), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n639), .B1(new_n626), .B2(new_n647), .ZN(G1326gat));
  AND2_X1   g447(.A1(new_n434), .A2(new_n436), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n626), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT43), .B(G22gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(G1327gat));
  NAND3_X1  g451(.A1(new_n603), .A2(new_n508), .A3(new_n625), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n471), .A2(new_n578), .A3(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n656), .A2(new_n532), .A3(new_n627), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT45), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n471), .A2(new_n578), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(KEYINPUT44), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT44), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n471), .A2(new_n661), .A3(new_n578), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n653), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(G29gat), .B1(new_n664), .B2(new_n389), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n658), .A2(new_n665), .ZN(G1328gat));
  OAI21_X1  g465(.A(G36gat), .B1(new_n664), .B2(new_n424), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n655), .A2(G36gat), .A3(new_n424), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT46), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(G1329gat));
  NAND2_X1  g469(.A1(new_n663), .A2(new_n646), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n469), .A2(G43gat), .ZN(new_n672));
  AOI22_X1  g471(.A1(new_n671), .A2(G43gat), .B1(new_n656), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n540), .B1(new_n663), .B2(new_n470), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n656), .A2(new_n672), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(KEYINPUT47), .ZN(new_n676));
  OAI22_X1  g475(.A1(new_n673), .A2(KEYINPUT47), .B1(new_n674), .B2(new_n676), .ZN(G1330gat));
  INV_X1    g476(.A(new_n649), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n655), .A2(G50gat), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n649), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n679), .B1(new_n680), .B2(G50gat), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n538), .B1(new_n663), .B2(new_n431), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT48), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  OAI22_X1  g483(.A1(new_n681), .A2(KEYINPUT48), .B1(new_n682), .B2(new_n684), .ZN(G1331gat));
  INV_X1    g484(.A(new_n625), .ZN(new_n686));
  AND3_X1   g485(.A1(new_n686), .A2(new_n579), .A3(new_n602), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n471), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT105), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n471), .A2(KEYINPUT105), .A3(new_n687), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n389), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n693), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g493(.A1(new_n692), .A2(new_n424), .ZN(new_n695));
  NOR2_X1   g494(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n696));
  AND2_X1   g495(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n695), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n698), .B1(new_n695), .B2(new_n696), .ZN(G1333gat));
  AND2_X1   g498(.A1(new_n643), .A2(new_n645), .ZN(new_n700));
  OAI21_X1  g499(.A(G71gat), .B1(new_n692), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n638), .A2(new_n480), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n701), .B1(new_n692), .B2(new_n702), .ZN(new_n703));
  XOR2_X1   g502(.A(KEYINPUT106), .B(KEYINPUT50), .Z(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n704), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n701), .B(new_n706), .C1(new_n692), .C2(new_n702), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(G1334gat));
  NOR2_X1   g507(.A1(new_n692), .A2(new_n678), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(new_n481), .ZN(G1335gat));
  INV_X1    g509(.A(new_n508), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n711), .A2(new_n625), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n471), .A2(new_n578), .A3(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT51), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n714), .A2(KEYINPUT108), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n715), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n471), .A2(new_n578), .A3(new_n712), .A4(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n714), .A2(KEYINPUT108), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n603), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n721), .A2(new_n381), .A3(new_n627), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n660), .A2(new_n662), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n712), .A2(new_n602), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT107), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(G85gat), .B1(new_n726), .B2(new_n389), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n722), .A2(new_n727), .ZN(G1336gat));
  NOR2_X1   g527(.A1(new_n424), .A2(G92gat), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  AOI211_X1 g529(.A(new_n603), .B(new_n730), .C1(new_n719), .C2(new_n720), .ZN(new_n731));
  INV_X1    g530(.A(new_n725), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n732), .B1(new_n660), .B2(new_n662), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n521), .B1(new_n733), .B2(new_n631), .ZN(new_n734));
  OAI21_X1  g533(.A(KEYINPUT52), .B1(new_n731), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n721), .A2(new_n729), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT52), .ZN(new_n737));
  OAI21_X1  g536(.A(G92gat), .B1(new_n726), .B2(new_n424), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n735), .A2(new_n739), .ZN(G1337gat));
  NAND3_X1  g539(.A1(new_n721), .A2(new_n259), .A3(new_n638), .ZN(new_n741));
  OAI21_X1  g540(.A(G99gat), .B1(new_n726), .B2(new_n700), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(G1338gat));
  NOR2_X1   g542(.A1(new_n257), .A2(G106gat), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n721), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n662), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n661), .B1(new_n471), .B2(new_n578), .ZN(new_n747));
  OAI211_X1 g546(.A(new_n431), .B(new_n725), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT53), .B1(new_n748), .B2(G106gat), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n733), .A2(new_n649), .ZN(new_n751));
  AOI22_X1  g550(.A1(new_n721), .A2(new_n744), .B1(new_n751), .B2(G106gat), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT53), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n750), .B1(new_n752), .B2(new_n753), .ZN(G1339gat));
  INV_X1    g553(.A(KEYINPUT54), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n755), .B(new_n582), .C1(new_n590), .C2(new_n592), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n756), .A2(new_n598), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n587), .A2(new_n589), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n591), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT110), .ZN(new_n760));
  INV_X1    g559(.A(new_n592), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n759), .A2(new_n760), .A3(new_n581), .A4(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n762), .A2(KEYINPUT54), .A3(new_n593), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n590), .A2(new_n592), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n760), .B1(new_n764), .B2(new_n581), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n757), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT55), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n757), .B(KEYINPUT55), .C1(new_n763), .C2(new_n765), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n768), .A2(new_n600), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n605), .B1(new_n604), .B2(new_n606), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n611), .A2(new_n613), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n620), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(KEYINPUT111), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT111), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n775), .B(new_n620), .C1(new_n771), .C2(new_n772), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n578), .A2(new_n774), .A3(new_n624), .A4(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(KEYINPUT112), .B1(new_n770), .B2(new_n777), .ZN(new_n778));
  AND4_X1   g577(.A1(new_n578), .A2(new_n774), .A3(new_n624), .A4(new_n776), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT112), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n599), .B1(new_n766), .B2(new_n767), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n779), .A2(new_n780), .A3(new_n781), .A4(new_n769), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n778), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n781), .A2(new_n625), .A3(new_n769), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n602), .A2(new_n774), .A3(new_n624), .A4(new_n776), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n578), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n508), .B1(new_n783), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n686), .A2(new_n603), .A3(new_n579), .ZN(new_n788));
  XOR2_X1   g587(.A(new_n788), .B(KEYINPUT109), .Z(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT113), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n787), .A2(new_n789), .A3(new_n792), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n425), .A2(new_n649), .A3(new_n389), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(G113gat), .B1(new_n796), .B2(new_n686), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n631), .A2(new_n389), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n794), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n363), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n686), .A2(G113gat), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n797), .B1(new_n801), .B2(new_n802), .ZN(G1340gat));
  OAI21_X1  g602(.A(G120gat), .B1(new_n796), .B2(new_n603), .ZN(new_n804));
  OR2_X1    g603(.A1(new_n603), .A2(G120gat), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n804), .B1(new_n801), .B2(new_n805), .ZN(G1341gat));
  INV_X1    g605(.A(G127gat), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n796), .A2(new_n807), .A3(new_n508), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n799), .A2(new_n800), .A3(new_n711), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n808), .B1(new_n809), .B2(new_n807), .ZN(G1342gat));
  INV_X1    g609(.A(new_n578), .ZN(new_n811));
  OR3_X1    g610(.A1(new_n801), .A2(G134gat), .A3(new_n811), .ZN(new_n812));
  OR2_X1    g611(.A1(new_n812), .A2(KEYINPUT56), .ZN(new_n813));
  OAI21_X1  g612(.A(G134gat), .B1(new_n796), .B2(new_n811), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(KEYINPUT56), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(G1343gat));
  NOR2_X1   g615(.A1(new_n646), .A2(new_n257), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n817), .A2(new_n799), .ZN(new_n818));
  INV_X1    g617(.A(G141gat), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n818), .A2(new_n819), .A3(new_n625), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n790), .A2(new_n649), .A3(KEYINPUT57), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n791), .A2(new_n431), .A3(new_n793), .ZN(new_n822));
  XOR2_X1   g621(.A(KEYINPUT115), .B(KEYINPUT57), .Z(new_n823));
  OAI21_X1  g622(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n798), .ZN(new_n825));
  OAI21_X1  g624(.A(KEYINPUT114), .B1(new_n470), .B2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT114), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n827), .B(new_n798), .C1(new_n642), .C2(new_n468), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n824), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n225), .B1(new_n829), .B2(new_n686), .ZN(new_n830));
  XNOR2_X1  g629(.A(KEYINPUT116), .B(KEYINPUT58), .ZN(new_n831));
  AND3_X1   g630(.A1(new_n820), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n831), .B1(new_n820), .B2(new_n830), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n832), .A2(new_n833), .ZN(G1344gat));
  NAND3_X1  g633(.A1(new_n818), .A2(new_n223), .A3(new_n602), .ZN(new_n835));
  XOR2_X1   g634(.A(KEYINPUT117), .B(KEYINPUT59), .Z(new_n836));
  NAND4_X1  g635(.A1(new_n791), .A2(new_n431), .A3(new_n793), .A4(new_n823), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT57), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n770), .A2(new_n777), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n508), .B1(new_n786), .B2(new_n839), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n840), .A2(new_n788), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n838), .B1(new_n678), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n837), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n843), .A2(new_n828), .A3(new_n602), .A4(new_n826), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(KEYINPUT118), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(G148gat), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n844), .A2(KEYINPUT118), .ZN(new_n847));
  OAI211_X1 g646(.A(KEYINPUT119), .B(new_n836), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n223), .A2(KEYINPUT59), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n849), .B1(new_n829), .B2(new_n603), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n223), .B1(new_n844), .B2(KEYINPUT118), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n852), .B1(KEYINPUT118), .B2(new_n844), .ZN(new_n853));
  AOI21_X1  g652(.A(KEYINPUT119), .B1(new_n853), .B2(new_n836), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n835), .B1(new_n851), .B2(new_n854), .ZN(G1345gat));
  NOR3_X1   g654(.A1(new_n829), .A2(new_n217), .A3(new_n508), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n818), .A2(new_n711), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n856), .B1(new_n857), .B2(new_n217), .ZN(G1346gat));
  NAND3_X1  g657(.A1(new_n818), .A2(new_n218), .A3(new_n578), .ZN(new_n859));
  OAI21_X1  g658(.A(G162gat), .B1(new_n829), .B2(new_n811), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(G1347gat));
  NOR2_X1   g660(.A1(new_n424), .A2(new_n627), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n638), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(KEYINPUT121), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n864), .A2(new_n678), .A3(new_n794), .ZN(new_n865));
  OAI21_X1  g664(.A(G169gat), .B1(new_n865), .B2(new_n686), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n794), .A2(new_n389), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n363), .A2(new_n424), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n868), .B(KEYINPUT120), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n870), .A2(new_n295), .A3(new_n625), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n866), .A2(new_n871), .ZN(G1348gat));
  NOR3_X1   g671(.A1(new_n865), .A2(new_n296), .A3(new_n603), .ZN(new_n873));
  AOI21_X1  g672(.A(G176gat), .B1(new_n870), .B2(new_n602), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n873), .A2(new_n874), .ZN(G1349gat));
  NAND2_X1  g674(.A1(new_n284), .A2(new_n287), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n711), .A2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT122), .B1(new_n870), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(G183gat), .B1(new_n865), .B2(new_n508), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g681(.A1(new_n870), .A2(new_n306), .A3(new_n578), .ZN(new_n883));
  OAI21_X1  g682(.A(G190gat), .B1(new_n865), .B2(new_n811), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(KEYINPUT61), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT123), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT61), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n887), .B(G190gat), .C1(new_n865), .C2(new_n811), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n885), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n888), .A2(new_n886), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n883), .B1(new_n889), .B2(new_n890), .ZN(G1351gat));
  NAND4_X1  g690(.A1(new_n700), .A2(new_n631), .A3(new_n867), .A4(new_n431), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n893), .A2(new_n617), .A3(new_n625), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n643), .A2(new_n645), .A3(new_n862), .ZN(new_n895));
  AOI22_X1  g694(.A1(new_n895), .A2(KEYINPUT124), .B1(new_n842), .B2(new_n837), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT124), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n643), .A2(new_n897), .A3(new_n645), .A4(new_n862), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n899), .A2(new_n625), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n894), .B1(new_n900), .B2(new_n617), .ZN(G1352gat));
  OR2_X1    g700(.A1(new_n603), .A2(G204gat), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n892), .A2(KEYINPUT62), .A3(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(KEYINPUT62), .B1(new_n892), .B2(new_n902), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT125), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI211_X1 g705(.A(KEYINPUT125), .B(KEYINPUT62), .C1(new_n892), .C2(new_n902), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n903), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n896), .A2(new_n602), .A3(new_n898), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n909), .A2(KEYINPUT126), .ZN(new_n910));
  OAI21_X1  g709(.A(G204gat), .B1(new_n909), .B2(KEYINPUT126), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(G1353gat));
  NAND3_X1  g711(.A1(new_n893), .A2(new_n205), .A3(new_n711), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n895), .A2(KEYINPUT124), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n914), .A2(new_n711), .A3(new_n843), .A4(new_n898), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT127), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n896), .A2(KEYINPUT127), .A3(new_n711), .A4(new_n898), .ZN(new_n918));
  AND4_X1   g717(.A1(KEYINPUT63), .A2(new_n917), .A3(G211gat), .A4(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n205), .B1(new_n915), .B2(new_n916), .ZN(new_n920));
  AOI21_X1  g719(.A(KEYINPUT63), .B1(new_n920), .B2(new_n918), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n913), .B1(new_n919), .B2(new_n921), .ZN(G1354gat));
  AOI21_X1  g721(.A(G218gat), .B1(new_n893), .B2(new_n578), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n811), .A2(new_n206), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n923), .B1(new_n899), .B2(new_n924), .ZN(G1355gat));
endmodule


