//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 0 0 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT82), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT78), .B1(new_n190), .B2(G104), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT78), .ZN(new_n192));
  INV_X1    g006(.A(G104), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G107), .ZN(new_n194));
  AND3_X1   g008(.A1(new_n190), .A2(KEYINPUT3), .A3(G104), .ZN(new_n195));
  AOI21_X1  g009(.A(KEYINPUT3), .B1(new_n190), .B2(G104), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n191), .B(new_n194), .C1(new_n195), .C2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G101), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(KEYINPUT4), .ZN(new_n199));
  AND3_X1   g013(.A1(new_n197), .A2(KEYINPUT79), .A3(new_n199), .ZN(new_n200));
  AOI21_X1  g014(.A(KEYINPUT79), .B1(new_n197), .B2(new_n199), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n202), .B1(new_n193), .B2(G107), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n190), .A2(KEYINPUT3), .A3(G104), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n205), .A2(new_n198), .A3(new_n191), .A4(new_n194), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT4), .ZN(new_n207));
  AND2_X1   g021(.A1(new_n191), .A2(new_n194), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n198), .B1(new_n208), .B2(new_n205), .ZN(new_n209));
  OAI22_X1  g023(.A1(new_n200), .A2(new_n201), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  XNOR2_X1  g024(.A(G116), .B(G119), .ZN(new_n211));
  INV_X1    g025(.A(G113), .ZN(new_n212));
  AND2_X1   g026(.A1(new_n212), .A2(KEYINPUT2), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n212), .A2(KEYINPUT2), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n211), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G119), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G116), .ZN(new_n217));
  INV_X1    g031(.A(G116), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G119), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT2), .B(G113), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n215), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n220), .A2(new_n221), .A3(KEYINPUT68), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n189), .B1(new_n210), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n211), .A2(KEYINPUT5), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n228), .B(G113), .C1(KEYINPUT5), .C2(new_n217), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n229), .A2(new_n215), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n193), .A2(G107), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n190), .A2(G104), .ZN(new_n232));
  OAI21_X1  g046(.A(G101), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n206), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n230), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n197), .A2(new_n199), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT79), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n197), .A2(KEYINPUT79), .A3(new_n199), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n226), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n197), .A2(G101), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(KEYINPUT4), .A3(new_n206), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n241), .A2(new_n242), .A3(KEYINPUT82), .A4(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n227), .A2(new_n236), .A3(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(G110), .B(G122), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n227), .A2(new_n247), .A3(new_n236), .A4(new_n245), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n249), .A2(KEYINPUT6), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT6), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n246), .A2(new_n252), .A3(new_n248), .ZN(new_n253));
  INV_X1    g067(.A(G146), .ZN(new_n254));
  AND2_X1   g068(.A1(KEYINPUT64), .A2(G143), .ZN(new_n255));
  NOR2_X1   g069(.A1(KEYINPUT64), .A2(G143), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G143), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G146), .ZN(new_n259));
  OAI21_X1  g073(.A(KEYINPUT1), .B1(new_n258), .B2(G146), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n257), .A2(new_n259), .B1(G128), .B2(new_n260), .ZN(new_n261));
  OR2_X1    g075(.A1(KEYINPUT64), .A2(G143), .ZN(new_n262));
  NAND2_X1  g076(.A1(KEYINPUT64), .A2(G143), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n262), .A2(KEYINPUT65), .A3(G146), .A4(new_n263), .ZN(new_n264));
  NOR3_X1   g078(.A1(new_n255), .A2(new_n256), .A3(new_n254), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT65), .B1(new_n254), .B2(G143), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n264), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT1), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G128), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n261), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G125), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n257), .A2(new_n259), .ZN(new_n275));
  AND2_X1   g089(.A1(KEYINPUT0), .A2(G128), .ZN(new_n276));
  NOR2_X1   g090(.A1(KEYINPUT0), .A2(G128), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n268), .A2(new_n276), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT66), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT66), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n268), .A2(new_n283), .A3(new_n276), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n280), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n274), .B1(new_n285), .B2(new_n273), .ZN(new_n286));
  INV_X1    g100(.A(G953), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G224), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n288), .B(KEYINPUT83), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n286), .B(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n251), .A2(new_n253), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n289), .A2(KEYINPUT7), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n286), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n293), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n274), .B(new_n295), .C1(new_n285), .C2(new_n273), .ZN(new_n296));
  XOR2_X1   g110(.A(KEYINPUT84), .B(KEYINPUT8), .Z(new_n297));
  XNOR2_X1  g111(.A(new_n297), .B(new_n247), .ZN(new_n298));
  INV_X1    g112(.A(new_n236), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n230), .A2(new_n235), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n294), .A2(new_n250), .A3(new_n296), .A4(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G902), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(KEYINPUT85), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n292), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(KEYINPUT85), .B1(new_n302), .B2(new_n303), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n188), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT86), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n302), .A2(new_n303), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT85), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n311), .A2(new_n187), .A3(new_n292), .A4(new_n304), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(new_n292), .A3(new_n304), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT86), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(new_n314), .A3(new_n188), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n308), .A2(new_n312), .A3(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(G214), .B1(G237), .B2(G902), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n317), .B(KEYINPUT81), .ZN(new_n318));
  AND2_X1   g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G469), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n285), .A2(new_n241), .A3(new_n244), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT11), .ZN(new_n322));
  INV_X1    g136(.A(G134), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n322), .B1(new_n323), .B2(G137), .ZN(new_n324));
  INV_X1    g138(.A(G137), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(KEYINPUT11), .A3(G134), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n323), .A2(G137), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n324), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G131), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n328), .B(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G128), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n331), .B1(new_n257), .B2(KEYINPUT1), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n268), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n262), .A2(new_n263), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n266), .B1(new_n334), .B2(new_n254), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n270), .B1(new_n335), .B2(new_n264), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n235), .B1(new_n333), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT10), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n268), .A2(new_n271), .ZN(new_n339));
  INV_X1    g153(.A(new_n261), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n234), .A2(new_n338), .ZN(new_n342));
  AOI22_X1  g156(.A1(new_n337), .A2(new_n338), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n321), .A2(new_n330), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n272), .A2(new_n234), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n337), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n330), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT12), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n287), .A2(G227), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n350), .B(KEYINPUT77), .ZN(new_n351));
  XNOR2_X1  g165(.A(G110), .B(G140), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n351), .B(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT12), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n346), .A2(new_n355), .A3(new_n347), .ZN(new_n356));
  AND4_X1   g170(.A1(new_n344), .A2(new_n349), .A3(new_n354), .A4(new_n356), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n268), .A2(new_n283), .A3(new_n276), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n283), .B1(new_n268), .B2(new_n276), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n279), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n360), .A2(new_n210), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n342), .A2(new_n341), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n269), .B1(new_n334), .B2(new_n254), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n335), .B(new_n264), .C1(new_n363), .C2(new_n331), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n234), .B1(new_n364), .B2(new_n339), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n362), .B1(new_n365), .B2(KEYINPUT10), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n347), .B1(new_n361), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n354), .B1(new_n367), .B2(new_n344), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n320), .B(new_n303), .C1(new_n357), .C2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(G469), .A2(G902), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n344), .A2(new_n349), .A3(new_n356), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n353), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n367), .A2(new_n344), .A3(new_n354), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(G469), .A3(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n369), .A2(new_n370), .A3(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT80), .ZN(new_n376));
  XNOR2_X1  g190(.A(KEYINPUT9), .B(G234), .ZN(new_n377));
  OAI21_X1  g191(.A(G221), .B1(new_n377), .B2(G902), .ZN(new_n378));
  AND3_X1   g192(.A1(new_n375), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n376), .B1(new_n375), .B2(new_n378), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G214), .ZN(new_n384));
  NOR3_X1   g198(.A1(new_n384), .A2(G237), .A3(G953), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G143), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n386), .B1(new_n334), .B2(new_n385), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G131), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT17), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n386), .B(new_n329), .C1(new_n334), .C2(new_n385), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT74), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(new_n273), .A3(G140), .ZN(new_n393));
  INV_X1    g207(.A(G140), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G125), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n273), .A2(G140), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI211_X1 g211(.A(KEYINPUT16), .B(new_n393), .C1(new_n397), .C2(new_n392), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT16), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G146), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n398), .A2(new_n254), .A3(new_n400), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n387), .A2(KEYINPUT17), .A3(G131), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n391), .A2(new_n402), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(G113), .B(G122), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n406), .B(new_n193), .ZN(new_n407));
  NAND2_X1  g221(.A1(KEYINPUT18), .A2(G131), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n387), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n408), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n386), .B(new_n410), .C1(new_n334), .C2(new_n385), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NOR3_X1   g226(.A1(new_n394), .A2(KEYINPUT74), .A3(G125), .ZN(new_n413));
  XNOR2_X1  g227(.A(G125), .B(G140), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n413), .B1(new_n414), .B2(KEYINPUT74), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G146), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n254), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n412), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n405), .A2(new_n407), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n407), .B1(new_n405), .B2(new_n419), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n303), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G475), .ZN(new_n424));
  AOI22_X1  g238(.A1(new_n388), .A2(new_n390), .B1(new_n401), .B2(G146), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT19), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n415), .A2(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n414), .A2(KEYINPUT19), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n254), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n425), .A2(new_n429), .B1(new_n418), .B2(new_n412), .ZN(new_n430));
  OAI21_X1  g244(.A(KEYINPUT87), .B1(new_n430), .B2(new_n407), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n388), .A2(new_n390), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n429), .A2(new_n402), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n419), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT87), .ZN(new_n435));
  INV_X1    g249(.A(new_n407), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n431), .A2(new_n420), .A3(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT20), .ZN(new_n439));
  NOR2_X1   g253(.A1(G475), .A2(G902), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n439), .B1(new_n438), .B2(new_n440), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n424), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n287), .A2(G952), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n445), .B1(G234), .B2(G237), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  XOR2_X1   g261(.A(KEYINPUT21), .B(G898), .Z(new_n448));
  NAND2_X1  g262(.A1(G234), .A2(G237), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(G902), .A3(G953), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n447), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  XOR2_X1   g265(.A(new_n451), .B(KEYINPUT93), .Z(new_n452));
  NAND2_X1  g266(.A1(new_n444), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(G478), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n454), .A2(KEYINPUT15), .ZN(new_n455));
  INV_X1    g269(.A(G217), .ZN(new_n456));
  NOR3_X1   g270(.A1(new_n377), .A2(new_n456), .A3(G953), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NOR3_X1   g272(.A1(new_n255), .A2(new_n256), .A3(new_n331), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n258), .A2(G128), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n323), .ZN(new_n462));
  XNOR2_X1  g276(.A(KEYINPUT88), .B(G122), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n463), .A2(new_n218), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n218), .A2(G122), .ZN(new_n465));
  OAI21_X1  g279(.A(G107), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NOR3_X1   g281(.A1(new_n464), .A2(G107), .A3(new_n465), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT89), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT13), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n460), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n470), .B1(new_n459), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n262), .A2(G128), .A3(new_n263), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n474), .B(KEYINPUT89), .C1(new_n471), .C2(new_n460), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT90), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n459), .A2(new_n476), .A3(KEYINPUT13), .ZN(new_n477));
  OAI21_X1  g291(.A(KEYINPUT90), .B1(new_n474), .B2(new_n471), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n473), .A2(new_n475), .A3(new_n477), .A4(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT91), .B1(new_n479), .B2(G134), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n479), .A2(KEYINPUT91), .A3(G134), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n469), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT14), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n464), .A2(new_n484), .ZN(new_n485));
  OR2_X1    g299(.A1(new_n466), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n461), .B(new_n323), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n464), .A2(new_n465), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n488), .B1(KEYINPUT14), .B2(new_n190), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n486), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n458), .B1(new_n483), .B2(new_n491), .ZN(new_n492));
  OR2_X1    g306(.A1(new_n467), .A2(new_n468), .ZN(new_n493));
  INV_X1    g307(.A(new_n482), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n493), .B(new_n462), .C1(new_n494), .C2(new_n480), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(new_n490), .A3(new_n457), .ZN(new_n496));
  AOI21_X1  g310(.A(G902), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n497), .A2(KEYINPUT92), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT92), .ZN(new_n499));
  AOI211_X1 g313(.A(new_n499), .B(G902), .C1(new_n492), .C2(new_n496), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n455), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  OAI22_X1  g315(.A1(new_n497), .A2(KEYINPUT92), .B1(KEYINPUT15), .B2(new_n454), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n453), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n319), .A2(new_n383), .A3(new_n504), .ZN(new_n505));
  OR2_X1    g319(.A1(new_n328), .A2(G131), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n325), .A2(KEYINPUT67), .A3(G134), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n327), .ZN(new_n508));
  AOI21_X1  g322(.A(KEYINPUT67), .B1(new_n325), .B2(G134), .ZN(new_n509));
  OAI21_X1  g323(.A(G131), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AND2_X1   g324(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n341), .A2(new_n511), .A3(KEYINPUT70), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT70), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n506), .A2(new_n510), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n513), .B1(new_n272), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n347), .B(new_n279), .C1(new_n358), .C2(new_n359), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT69), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n282), .A2(new_n284), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n520), .A2(KEYINPUT69), .A3(new_n279), .A4(new_n347), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n516), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n522), .A2(new_n226), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n522), .A2(new_n226), .ZN(new_n524));
  OAI21_X1  g338(.A(KEYINPUT28), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT28), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n517), .B1(new_n272), .B2(new_n514), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n526), .B1(new_n527), .B2(new_n242), .ZN(new_n528));
  XOR2_X1   g342(.A(KEYINPUT26), .B(G101), .Z(new_n529));
  INV_X1    g343(.A(G237), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n530), .A2(new_n287), .A3(G210), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n529), .B(new_n531), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n532), .B(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT29), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n525), .A2(new_n528), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n522), .A2(new_n226), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n527), .A2(new_n242), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n526), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n534), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n528), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n535), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT30), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n519), .A2(new_n521), .ZN(new_n545));
  INV_X1    g359(.A(new_n516), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n527), .A2(KEYINPUT30), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n242), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n541), .B1(new_n549), .B2(new_n538), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n537), .B(new_n303), .C1(new_n543), .C2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT72), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n551), .A2(new_n552), .A3(G472), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n552), .B1(new_n551), .B2(G472), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n534), .B1(new_n522), .B2(new_n226), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n549), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(KEYINPUT31), .ZN(new_n557));
  INV_X1    g371(.A(new_n528), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n534), .B1(new_n540), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT31), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n549), .A2(new_n560), .A3(new_n555), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n557), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT32), .ZN(new_n563));
  NOR2_X1   g377(.A1(G472), .A2(G902), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n563), .B1(new_n562), .B2(new_n564), .ZN(new_n566));
  OAI22_X1  g380(.A1(new_n553), .A2(new_n554), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n402), .A2(new_n403), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n216), .A2(G128), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT23), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n331), .A2(G119), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT73), .ZN(new_n572));
  XOR2_X1   g386(.A(new_n570), .B(new_n572), .Z(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(G110), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n569), .A2(new_n571), .ZN(new_n575));
  XNOR2_X1  g389(.A(KEYINPUT24), .B(G110), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n568), .B(new_n574), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n575), .A2(new_n576), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(KEYINPUT75), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n579), .B1(G110), .B2(new_n573), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n580), .A2(new_n402), .A3(new_n417), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n287), .A2(G221), .A3(G234), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(KEYINPUT76), .ZN(new_n583));
  XNOR2_X1  g397(.A(KEYINPUT22), .B(G137), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n583), .B(new_n584), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n577), .A2(new_n581), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n585), .B1(new_n577), .B2(new_n581), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n589), .A2(KEYINPUT25), .A3(new_n303), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT25), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n591), .B1(new_n588), .B2(G902), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n456), .B1(G234), .B2(new_n303), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n594), .A2(G902), .ZN(new_n595));
  AOI22_X1  g409(.A1(new_n593), .A2(new_n594), .B1(new_n589), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n567), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n505), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g412(.A(KEYINPUT94), .B(G101), .Z(new_n599));
  XNOR2_X1  g413(.A(new_n598), .B(new_n599), .ZN(G3));
  NOR3_X1   g414(.A1(new_n483), .A2(new_n491), .A3(new_n458), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n457), .B1(new_n495), .B2(new_n490), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n303), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n603), .A2(KEYINPUT96), .A3(new_n454), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT96), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n605), .B1(new_n497), .B2(G478), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(KEYINPUT33), .B1(new_n601), .B2(new_n602), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT33), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n492), .A2(new_n496), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n454), .A2(G902), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI211_X1 g427(.A(KEYINPUT97), .B(new_n443), .C1(new_n607), .C2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT97), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n604), .A2(new_n606), .B1(new_n611), .B2(new_n612), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n615), .B1(new_n616), .B2(new_n444), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT95), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n307), .A2(new_n619), .A3(new_n312), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n313), .A2(KEYINPUT95), .A3(new_n188), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n620), .A2(new_n317), .A3(new_n452), .A4(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n562), .A2(new_n564), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n549), .A2(new_n560), .A3(new_n555), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n560), .B1(new_n549), .B2(new_n555), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(G902), .B1(new_n627), .B2(new_n559), .ZN(new_n628));
  INV_X1    g442(.A(G472), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n624), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n596), .B1(new_n379), .B2(new_n381), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n623), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT34), .B(G104), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G6));
  INV_X1    g449(.A(new_n452), .ZN(new_n636));
  AOI211_X1 g450(.A(new_n636), .B(new_n443), .C1(new_n501), .C2(new_n502), .ZN(new_n637));
  AND4_X1   g451(.A1(new_n317), .A2(new_n637), .A3(new_n620), .A4(new_n621), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n632), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT35), .B(G107), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G9));
  AOI21_X1  g455(.A(new_n629), .B1(new_n562), .B2(new_n303), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n642), .B1(new_n564), .B2(new_n562), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n593), .A2(new_n594), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n577), .A2(new_n581), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n585), .A2(KEYINPUT36), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n595), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n650), .A2(new_n453), .A3(new_n503), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n319), .A2(new_n643), .A3(new_n383), .A4(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT37), .B(G110), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G12));
  OAI21_X1  g468(.A(new_n649), .B1(new_n379), .B2(new_n381), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n551), .A2(G472), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(KEYINPUT72), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n551), .A2(new_n552), .A3(G472), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n566), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n655), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  OR2_X1    g477(.A1(new_n450), .A2(G900), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n447), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n503), .A2(new_n444), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(KEYINPUT98), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT98), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n503), .A2(new_n668), .A3(new_n444), .A4(new_n665), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n620), .A2(new_n317), .A3(new_n621), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n663), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  NAND2_X1  g488(.A1(new_n503), .A2(new_n443), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n650), .A2(new_n317), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n665), .B(KEYINPUT39), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n383), .A2(new_n677), .ZN(new_n678));
  AOI211_X1 g492(.A(new_n675), .B(new_n676), .C1(new_n678), .C2(KEYINPUT40), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n316), .B(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  OR2_X1    g496(.A1(new_n678), .A2(KEYINPUT40), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n549), .A2(new_n538), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n684), .A2(new_n534), .ZN(new_n685));
  OR2_X1    g499(.A1(new_n523), .A2(new_n524), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n303), .B1(new_n686), .B2(new_n541), .ZN(new_n687));
  OAI21_X1  g501(.A(G472), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n662), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n679), .A2(new_n682), .A3(new_n683), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(new_n334), .ZN(G45));
  NOR2_X1   g505(.A1(new_n616), .A2(new_n444), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n665), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n671), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n663), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G146), .ZN(G48));
  OR2_X1    g511(.A1(new_n357), .A2(new_n368), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n320), .B1(new_n698), .B2(new_n303), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n369), .A2(KEYINPUT100), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AOI211_X1 g515(.A(KEYINPUT100), .B(new_n320), .C1(new_n698), .C2(new_n303), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n378), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n623), .A2(new_n567), .A3(new_n596), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT41), .B(G113), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G15));
  NAND4_X1  g521(.A1(new_n638), .A2(new_n567), .A3(new_n596), .A4(new_n704), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G116), .ZN(G18));
  NOR2_X1   g523(.A1(new_n671), .A2(new_n703), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n567), .A2(new_n710), .A3(new_n651), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G119), .ZN(G21));
  NOR3_X1   g526(.A1(new_n622), .A2(new_n703), .A3(new_n675), .ZN(new_n713));
  INV_X1    g527(.A(new_n564), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n525), .A2(new_n528), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n534), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n714), .B1(new_n627), .B2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n596), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n642), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n713), .A2(new_n719), .ZN(new_n720));
  XOR2_X1   g534(.A(KEYINPUT101), .B(G122), .Z(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G24));
  NOR3_X1   g536(.A1(new_n642), .A2(new_n650), .A3(new_n717), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n693), .A2(new_n694), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n710), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G125), .ZN(G27));
  AND2_X1   g540(.A1(new_n312), .A2(new_n317), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n308), .A2(new_n727), .A3(new_n315), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(KEYINPUT104), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT104), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n308), .A2(new_n727), .A3(new_n730), .A4(new_n315), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n373), .A2(KEYINPUT102), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT102), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n367), .A2(new_n344), .A3(new_n733), .A4(new_n354), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n732), .A2(new_n372), .A3(new_n734), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n369), .B(new_n370), .C1(new_n735), .C2(new_n320), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n736), .A2(KEYINPUT103), .A3(new_n378), .ZN(new_n737));
  AOI21_X1  g551(.A(KEYINPUT103), .B1(new_n736), .B2(new_n378), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n729), .A2(new_n731), .A3(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n718), .B1(new_n659), .B2(new_n662), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n741), .A2(new_n742), .A3(new_n724), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT42), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n741), .A2(new_n742), .A3(KEYINPUT42), .A4(new_n724), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G131), .ZN(G33));
  INV_X1    g562(.A(new_n670), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n741), .A2(new_n742), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G134), .ZN(G36));
  NAND2_X1  g565(.A1(new_n729), .A2(new_n731), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n616), .A2(new_n443), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(KEYINPUT43), .ZN(new_n754));
  XOR2_X1   g568(.A(new_n754), .B(KEYINPUT105), .Z(new_n755));
  NAND3_X1  g569(.A1(new_n755), .A2(new_n630), .A3(new_n649), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT44), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n752), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n758), .B1(new_n757), .B2(new_n756), .ZN(new_n759));
  OR2_X1    g573(.A1(new_n759), .A2(KEYINPUT106), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(KEYINPUT106), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT45), .ZN(new_n762));
  OR2_X1    g576(.A1(new_n735), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n372), .A2(new_n373), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n762), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n763), .A2(G469), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n370), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT46), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n369), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n767), .A2(new_n768), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n378), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n677), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n760), .A2(new_n761), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G137), .ZN(G39));
  XNOR2_X1  g590(.A(new_n772), .B(KEYINPUT47), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n724), .A2(new_n718), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n752), .A2(new_n779), .A3(new_n567), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n780), .A2(KEYINPUT107), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(KEYINPUT107), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n778), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G140), .ZN(G42));
  OAI21_X1  g598(.A(new_n663), .B1(new_n672), .B2(new_n695), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n671), .A2(new_n675), .ZN(new_n786));
  AND4_X1   g600(.A1(new_n378), .A2(new_n650), .A3(new_n665), .A4(new_n736), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n689), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n785), .A2(new_n725), .A3(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n785), .A2(KEYINPUT52), .A3(new_n725), .A4(new_n788), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n791), .A2(KEYINPUT112), .A3(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT112), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n789), .A2(new_n794), .A3(new_n790), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n655), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n503), .A2(new_n443), .A3(new_n694), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n567), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n723), .A2(new_n724), .ZN(new_n800));
  OAI22_X1  g614(.A1(new_n799), .A2(new_n752), .B1(new_n800), .B2(new_n740), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n597), .A2(new_n740), .A3(new_n670), .ZN(new_n802));
  OAI21_X1  g616(.A(KEYINPUT110), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n741), .A2(new_n724), .A3(new_n723), .ZN(new_n804));
  INV_X1    g618(.A(new_n752), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n663), .A2(new_n805), .A3(new_n798), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT110), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n750), .A2(new_n804), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n803), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n316), .A2(new_n318), .A3(new_n637), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT108), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT108), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n316), .A2(new_n637), .A3(new_n812), .A4(new_n318), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n811), .A2(new_n632), .A3(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT109), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n814), .A2(new_n815), .A3(new_n652), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n815), .B1(new_n814), .B2(new_n652), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n319), .A2(new_n383), .A3(new_n643), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n692), .A2(new_n596), .A3(new_n452), .ZN(new_n819));
  OAI22_X1  g633(.A1(new_n597), .A2(new_n505), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n816), .A2(new_n817), .A3(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n705), .A2(new_n708), .A3(new_n720), .A4(new_n711), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n822), .B1(new_n745), .B2(new_n746), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n809), .A2(new_n821), .A3(KEYINPUT53), .A4(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n796), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n809), .A2(new_n821), .A3(new_n823), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT111), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n809), .A2(new_n821), .A3(new_n823), .A4(KEYINPUT111), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n791), .A2(new_n792), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT53), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n825), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n834), .A2(KEYINPUT113), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n825), .ZN(new_n837));
  INV_X1    g651(.A(new_n831), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n838), .B1(new_n828), .B2(new_n829), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n835), .B(new_n837), .C1(new_n839), .C2(KEYINPUT53), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT113), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n832), .A2(KEYINPUT53), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n830), .A2(new_n833), .A3(new_n795), .A4(new_n793), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n843), .A2(KEYINPUT54), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n836), .A2(new_n842), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT114), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n846), .B(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n752), .A2(new_n703), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  NOR4_X1   g664(.A1(new_n850), .A2(new_n718), .A3(new_n447), .A4(new_n689), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT115), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n852), .A2(new_n444), .A3(new_n616), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n754), .A2(new_n719), .A3(new_n446), .ZN(new_n854));
  NOR4_X1   g668(.A1(new_n682), .A2(new_n854), .A3(new_n317), .A4(new_n703), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(KEYINPUT50), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n699), .B(new_n700), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n777), .B1(new_n378), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n854), .A2(new_n752), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n849), .A2(new_n446), .A3(new_n754), .ZN(new_n861));
  AOI22_X1  g675(.A1(new_n859), .A2(new_n860), .B1(new_n723), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n853), .A2(new_n856), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT51), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n863), .A2(new_n864), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n445), .B(KEYINPUT116), .ZN(new_n867));
  INV_X1    g681(.A(new_n710), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n867), .B1(new_n854), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n861), .A2(new_n742), .ZN(new_n870));
  XOR2_X1   g684(.A(new_n870), .B(KEYINPUT48), .Z(new_n871));
  INV_X1    g685(.A(new_n618), .ZN(new_n872));
  AOI211_X1 g686(.A(new_n869), .B(new_n871), .C1(new_n872), .C2(new_n852), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n865), .A2(new_n866), .A3(new_n873), .ZN(new_n874));
  OAI22_X1  g688(.A1(new_n848), .A2(new_n874), .B1(G952), .B2(G953), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n857), .B(KEYINPUT49), .Z(new_n876));
  NAND4_X1  g690(.A1(new_n753), .A2(new_n596), .A3(new_n318), .A4(new_n378), .ZN(new_n877));
  OR4_X1    g691(.A1(new_n682), .A2(new_n876), .A3(new_n689), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n875), .A2(new_n878), .ZN(G75));
  NOR2_X1   g693(.A1(new_n287), .A2(G952), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n251), .A2(new_n253), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(new_n291), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n882), .B(KEYINPUT55), .Z(new_n883));
  OAI21_X1  g697(.A(new_n837), .B1(new_n839), .B2(KEYINPUT53), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n884), .A2(G210), .A3(G902), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT56), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n883), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(KEYINPUT117), .B1(new_n834), .B2(new_n303), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT117), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n884), .A2(new_n889), .A3(G902), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n888), .A2(new_n188), .A3(new_n890), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n883), .A2(new_n886), .ZN(new_n892));
  AOI211_X1 g706(.A(new_n880), .B(new_n887), .C1(new_n891), .C2(new_n892), .ZN(G51));
  INV_X1    g707(.A(new_n766), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n888), .A2(new_n894), .A3(new_n890), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(KEYINPUT119), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT119), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n888), .A2(new_n897), .A3(new_n894), .A4(new_n890), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n884), .A2(KEYINPUT54), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n840), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n370), .B(KEYINPUT118), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT57), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n698), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n896), .A2(new_n898), .A3(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n880), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT120), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n905), .A2(KEYINPUT120), .A3(new_n906), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(G54));
  NAND4_X1  g725(.A1(new_n888), .A2(KEYINPUT58), .A3(G475), .A4(new_n890), .ZN(new_n912));
  INV_X1    g726(.A(new_n438), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n912), .A2(new_n913), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n914), .A2(new_n915), .A3(new_n880), .ZN(G60));
  NAND2_X1  g730(.A1(G478), .A2(G902), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT59), .Z(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n611), .B1(new_n848), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n900), .A2(new_n611), .A3(new_n919), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(new_n906), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n920), .A2(new_n922), .ZN(G63));
  XNOR2_X1  g737(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n924));
  NAND2_X1  g738(.A1(G217), .A2(G902), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT122), .Z(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT60), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n834), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n647), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n906), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n928), .A2(new_n589), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n924), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT123), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(KEYINPUT61), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n906), .B(new_n929), .C1(new_n931), .C2(new_n933), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n932), .B1(new_n935), .B2(new_n936), .ZN(G66));
  AOI21_X1  g751(.A(new_n287), .B1(new_n448), .B2(G224), .ZN(new_n938));
  INV_X1    g752(.A(new_n821), .ZN(new_n939));
  OR2_X1    g753(.A1(new_n939), .A2(new_n822), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n938), .B1(new_n940), .B2(new_n287), .ZN(new_n941));
  INV_X1    g755(.A(G898), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n881), .B1(new_n942), .B2(G953), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n941), .B(new_n943), .ZN(G69));
  NOR2_X1   g758(.A1(new_n547), .A2(new_n548), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n427), .A2(new_n428), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT124), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n945), .B(new_n947), .Z(new_n948));
  NAND2_X1  g762(.A1(new_n785), .A2(new_n725), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n690), .ZN(new_n951));
  OR2_X1    g765(.A1(new_n951), .A2(KEYINPUT62), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(KEYINPUT62), .ZN(new_n953));
  INV_X1    g767(.A(new_n783), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n692), .B1(new_n503), .B2(new_n444), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n597), .A2(new_n678), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n954), .B1(new_n805), .B2(new_n956), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n775), .A2(new_n952), .A3(new_n953), .A4(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n948), .B1(new_n958), .B2(new_n287), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n774), .A2(new_n742), .A3(new_n786), .ZN(new_n960));
  AND4_X1   g774(.A1(new_n750), .A2(new_n783), .A3(new_n950), .A4(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n775), .A2(new_n747), .A3(new_n961), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n962), .A2(G953), .ZN(new_n963));
  INV_X1    g777(.A(new_n948), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n964), .B1(G900), .B2(G953), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n959), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n287), .B1(G227), .B2(G900), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n966), .B(new_n967), .Z(G72));
  XNOR2_X1  g782(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n629), .A2(new_n303), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n969), .B(new_n970), .Z(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT126), .Z(new_n972));
  OAI21_X1  g786(.A(new_n972), .B1(new_n958), .B2(new_n940), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n880), .B1(new_n973), .B2(new_n685), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n972), .B1(new_n962), .B2(new_n940), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n975), .A2(KEYINPUT127), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n684), .A2(new_n534), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n977), .B1(new_n975), .B2(KEYINPUT127), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n974), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n843), .A2(new_n844), .ZN(new_n980));
  INV_X1    g794(.A(new_n971), .ZN(new_n981));
  NOR3_X1   g795(.A1(new_n977), .A2(new_n685), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n979), .B1(new_n980), .B2(new_n982), .ZN(G57));
endmodule


