

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785;

  XNOR2_X1 U361 ( .A(n647), .B(n442), .ZN(n339) );
  NAND2_X1 U362 ( .A1(n343), .A2(n430), .ZN(n429) );
  NOR2_X1 U363 ( .A1(n690), .A2(n344), .ZN(n343) );
  INV_X1 U364 ( .A(KEYINPUT84), .ZN(n344) );
  AND2_X1 U365 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U366 ( .A1(n625), .A2(n713), .ZN(n628) );
  XOR2_X1 U367 ( .A(KEYINPUT69), .B(KEYINPUT22), .Z(n619) );
  AND2_X1 U368 ( .A1(n463), .A2(n461), .ZN(n459) );
  XNOR2_X1 U369 ( .A(n444), .B(n391), .ZN(n674) );
  XNOR2_X2 U370 ( .A(n537), .B(n536), .ZN(n347) );
  NAND2_X1 U371 ( .A1(n418), .A2(n464), .ZN(n342) );
  NAND2_X1 U372 ( .A1(n725), .A2(n580), .ZN(n425) );
  XNOR2_X2 U373 ( .A(n586), .B(n540), .ZN(n725) );
  NAND2_X2 U374 ( .A1(n339), .A2(n338), .ZN(n396) );
  XNOR2_X2 U375 ( .A(n414), .B(KEYINPUT45), .ZN(n338) );
  XNOR2_X2 U376 ( .A(n390), .B(n584), .ZN(n658) );
  NOR2_X2 U377 ( .A1(n785), .A2(n658), .ZN(n585) );
  NAND2_X1 U378 ( .A1(n340), .A2(n465), .ZN(n418) );
  NAND2_X1 U379 ( .A1(n427), .A2(n429), .ZN(n340) );
  AND2_X2 U380 ( .A1(n396), .A2(n452), .ZN(n451) );
  AND2_X2 U381 ( .A1(n424), .A2(n423), .ZN(n389) );
  AND2_X2 U382 ( .A1(n490), .A2(n646), .ZN(n647) );
  NOR2_X2 U383 ( .A1(n396), .A2(n649), .ZN(n449) );
  AND2_X2 U384 ( .A1(n341), .A2(n622), .ZN(n690) );
  XNOR2_X1 U385 ( .A(n638), .B(n621), .ZN(n341) );
  NAND2_X2 U386 ( .A1(n433), .A2(n432), .ZN(n431) );
  NAND2_X2 U387 ( .A1(n342), .A2(n415), .ZN(n414) );
  XNOR2_X2 U388 ( .A(n620), .B(n619), .ZN(n625) );
  XNOR2_X2 U389 ( .A(n547), .B(n546), .ZN(n426) );
  XNOR2_X1 U390 ( .A(n530), .B(n529), .ZN(n393) );
  NOR2_X1 U391 ( .A1(n588), .A2(n643), .ZN(n575) );
  INV_X2 U392 ( .A(G953), .ZN(n779) );
  NOR2_X1 U393 ( .A1(n445), .A2(n449), .ZN(n443) );
  XNOR2_X1 U394 ( .A(n412), .B(n411), .ZN(n498) );
  NAND2_X1 U395 ( .A1(n486), .A2(n482), .ZN(n643) );
  OR2_X1 U396 ( .A1(n661), .A2(n483), .ZN(n482) );
  NOR2_X1 U397 ( .A1(n664), .A2(n757), .ZN(n667) );
  NOR2_X1 U398 ( .A1(n672), .A2(n757), .ZN(n673) );
  NOR2_X1 U399 ( .A1(n654), .A2(n757), .ZN(n656) );
  NOR2_X1 U400 ( .A1(n679), .A2(n757), .ZN(n680) );
  NAND2_X1 U401 ( .A1(n357), .A2(n455), .ZN(n453) );
  INV_X1 U402 ( .A(n498), .ZN(n345) );
  XNOR2_X1 U403 ( .A(n643), .B(n587), .ZN(n639) );
  XNOR2_X1 U404 ( .A(n676), .B(n675), .ZN(n677) );
  AND2_X1 U405 ( .A1(n488), .A2(n487), .ZN(n486) );
  XNOR2_X1 U406 ( .A(n559), .B(n495), .ZN(n624) );
  XNOR2_X1 U407 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U408 ( .A(n511), .B(n469), .ZN(n669) );
  XNOR2_X1 U409 ( .A(n470), .B(n553), .ZN(n469) );
  XNOR2_X1 U410 ( .A(n524), .B(n491), .ZN(n553) );
  XNOR2_X2 U411 ( .A(KEYINPUT3), .B(KEYINPUT67), .ZN(n528) );
  NOR2_X1 U412 ( .A1(G237), .A2(G953), .ZN(n508) );
  NAND2_X2 U413 ( .A1(n459), .A2(n458), .ZN(n631) );
  AND2_X1 U414 ( .A1(n439), .A2(n725), .ZN(n544) );
  NAND2_X1 U415 ( .A1(n400), .A2(n407), .ZN(n399) );
  NAND2_X1 U416 ( .A1(n367), .A2(n403), .ZN(n402) );
  NOR2_X1 U417 ( .A1(n695), .A2(n401), .ZN(n400) );
  XNOR2_X1 U418 ( .A(n474), .B(G134), .ZN(n772) );
  NAND2_X1 U419 ( .A1(n550), .A2(G217), .ZN(n365) );
  XOR2_X1 U420 ( .A(G137), .B(G140), .Z(n554) );
  XNOR2_X1 U421 ( .A(n772), .B(G146), .ZN(n572) );
  XNOR2_X1 U422 ( .A(n468), .B(G146), .ZN(n524) );
  INV_X1 U423 ( .A(G125), .ZN(n468) );
  NAND2_X1 U424 ( .A1(n582), .A2(n426), .ZN(n394) );
  NOR2_X1 U425 ( .A1(n480), .A2(n479), .ZN(n478) );
  AND2_X1 U426 ( .A1(n417), .A2(n416), .ZN(n415) );
  AND2_X1 U427 ( .A1(n681), .A2(n378), .ZN(n416) );
  XNOR2_X1 U428 ( .A(n426), .B(KEYINPUT1), .ZN(n633) );
  NAND2_X1 U429 ( .A1(n493), .A2(n492), .ZN(n604) );
  AND2_X1 U430 ( .A1(n699), .A2(n724), .ZN(n492) );
  XNOR2_X1 U431 ( .A(n410), .B(KEYINPUT106), .ZN(n493) );
  NOR2_X1 U432 ( .A1(n639), .A2(n588), .ZN(n410) );
  NOR2_X1 U433 ( .A1(n368), .A2(n728), .ZN(n594) );
  XNOR2_X1 U434 ( .A(n534), .B(G902), .ZN(n648) );
  INV_X1 U435 ( .A(KEYINPUT15), .ZN(n534) );
  INV_X1 U436 ( .A(G237), .ZN(n535) );
  NAND2_X1 U437 ( .A1(n569), .A2(G210), .ZN(n473) );
  XNOR2_X1 U438 ( .A(n528), .B(n527), .ZN(n530) );
  XNOR2_X1 U439 ( .A(KEYINPUT9), .B(KEYINPUT100), .ZN(n467) );
  XNOR2_X1 U440 ( .A(n516), .B(n515), .ZN(n364) );
  XNOR2_X1 U441 ( .A(G134), .B(G107), .ZN(n515) );
  XNOR2_X1 U442 ( .A(n533), .B(n500), .ZN(n499) );
  XNOR2_X1 U443 ( .A(n525), .B(n501), .ZN(n500) );
  INV_X1 U444 ( .A(KEYINPUT18), .ZN(n501) );
  NAND2_X1 U445 ( .A1(n498), .A2(n497), .ZN(n465) );
  NAND2_X1 U446 ( .A1(n457), .A2(n460), .ZN(n458) );
  OR2_X1 U447 ( .A1(n346), .A2(n462), .ZN(n461) );
  NAND2_X1 U448 ( .A1(n485), .A2(n484), .ZN(n483) );
  NAND2_X1 U449 ( .A1(n574), .A2(G902), .ZN(n487) );
  INV_X1 U450 ( .A(KEYINPUT80), .ZN(n420) );
  XNOR2_X1 U451 ( .A(n393), .B(n502), .ZN(n762) );
  XNOR2_X1 U452 ( .A(G122), .B(KEYINPUT16), .ZN(n502) );
  XNOR2_X1 U453 ( .A(n372), .B(n371), .ZN(n370) );
  XNOR2_X1 U454 ( .A(KEYINPUT94), .B(KEYINPUT92), .ZN(n371) );
  XNOR2_X1 U455 ( .A(n373), .B(G110), .ZN(n372) );
  INV_X1 U456 ( .A(KEYINPUT24), .ZN(n373) );
  XNOR2_X1 U457 ( .A(n548), .B(n549), .ZN(n374) );
  XNOR2_X1 U458 ( .A(n514), .B(n366), .ZN(n550) );
  INV_X1 U459 ( .A(KEYINPUT8), .ZN(n366) );
  INV_X1 U460 ( .A(KEYINPUT10), .ZN(n491) );
  XNOR2_X1 U461 ( .A(n545), .B(n572), .ZN(n489) );
  XNOR2_X1 U462 ( .A(n558), .B(n496), .ZN(n495) );
  INV_X1 U463 ( .A(KEYINPUT25), .ZN(n496) );
  INV_X1 U464 ( .A(KEYINPUT81), .ZN(n442) );
  INV_X1 U465 ( .A(n453), .ZN(n742) );
  INV_X1 U466 ( .A(n604), .ZN(n407) );
  NOR2_X1 U467 ( .A1(n607), .A2(n351), .ZN(n406) );
  NAND2_X1 U468 ( .A1(n397), .A2(n404), .ZN(n367) );
  AND2_X1 U469 ( .A1(n633), .A2(n405), .ZN(n404) );
  NAND2_X1 U470 ( .A1(n604), .A2(n351), .ZN(n397) );
  NAND2_X1 U471 ( .A1(n369), .A2(n457), .ZN(n368) );
  INV_X1 U472 ( .A(n591), .ZN(n369) );
  AND2_X1 U473 ( .A1(n593), .A2(n592), .ZN(n699) );
  INV_X1 U474 ( .A(n406), .ZN(n401) );
  INV_X1 U475 ( .A(n695), .ZN(n403) );
  NAND2_X1 U476 ( .A1(G224), .A2(n779), .ZN(n525) );
  AND2_X1 U477 ( .A1(n409), .A2(n408), .ZN(n600) );
  XNOR2_X1 U478 ( .A(n594), .B(KEYINPUT47), .ZN(n408) );
  AND2_X1 U479 ( .A1(n346), .A2(n462), .ZN(n460) );
  NOR2_X1 U480 ( .A1(n486), .A2(KEYINPUT30), .ZN(n479) );
  NOR2_X1 U481 ( .A1(n581), .A2(n481), .ZN(n477) );
  INV_X1 U482 ( .A(KEYINPUT30), .ZN(n481) );
  NAND2_X1 U483 ( .A1(n556), .A2(KEYINPUT65), .ZN(n446) );
  NOR2_X1 U484 ( .A1(n649), .A2(KEYINPUT2), .ZN(n448) );
  NAND2_X1 U485 ( .A1(n380), .A2(n379), .ZN(n378) );
  INV_X1 U486 ( .A(n728), .ZN(n379) );
  NAND2_X1 U487 ( .A1(n382), .A2(n381), .ZN(n380) );
  INV_X1 U488 ( .A(n687), .ZN(n381) );
  INV_X1 U489 ( .A(KEYINPUT19), .ZN(n589) );
  XNOR2_X1 U490 ( .A(n387), .B(n472), .ZN(n386) );
  XNOR2_X1 U491 ( .A(n393), .B(n572), .ZN(n387) );
  XNOR2_X1 U492 ( .A(n363), .B(n361), .ZN(n650) );
  XNOR2_X1 U493 ( .A(n365), .B(n364), .ZN(n363) );
  XNOR2_X1 U494 ( .A(n467), .B(KEYINPUT7), .ZN(n362) );
  XOR2_X1 U495 ( .A(KEYINPUT98), .B(G104), .Z(n507) );
  XNOR2_X1 U496 ( .A(G143), .B(G131), .ZN(n506) );
  XNOR2_X1 U497 ( .A(n505), .B(n471), .ZN(n470) );
  XNOR2_X1 U498 ( .A(KEYINPUT12), .B(KEYINPUT11), .ZN(n471) );
  INV_X1 U499 ( .A(G140), .ZN(n503) );
  XNOR2_X1 U500 ( .A(n762), .B(n392), .ZN(n391) );
  XNOR2_X1 U501 ( .A(n499), .B(n526), .ZN(n392) );
  XNOR2_X1 U502 ( .A(n542), .B(KEYINPUT41), .ZN(n543) );
  NOR2_X1 U503 ( .A1(n394), .A2(KEYINPUT39), .ZN(n421) );
  NAND2_X1 U504 ( .A1(n494), .A2(n712), .ZN(n709) );
  INV_X1 U505 ( .A(n624), .ZN(n494) );
  INV_X1 U506 ( .A(n778), .ZN(n419) );
  XNOR2_X1 U507 ( .A(n374), .B(n370), .ZN(n552) );
  XOR2_X1 U508 ( .A(KEYINPUT122), .B(n650), .Z(n651) );
  INV_X1 U509 ( .A(KEYINPUT35), .ZN(n411) );
  NAND2_X1 U510 ( .A1(n413), .A2(n637), .ZN(n412) );
  XNOR2_X1 U511 ( .A(n636), .B(KEYINPUT34), .ZN(n413) );
  NOR2_X1 U512 ( .A1(n710), .A2(n626), .ZN(n627) );
  XNOR2_X1 U513 ( .A(n435), .B(KEYINPUT31), .ZN(n703) );
  XNOR2_X1 U514 ( .A(n384), .B(KEYINPUT83), .ZN(n383) );
  XNOR2_X1 U515 ( .A(n751), .B(n353), .ZN(n752) );
  AND2_X1 U516 ( .A1(n396), .A2(n743), .ZN(n744) );
  AND2_X1 U517 ( .A1(n407), .A2(n406), .ZN(n398) );
  INV_X1 U518 ( .A(n699), .ZN(n697) );
  OR2_X1 U519 ( .A1(n614), .A2(n613), .ZN(n346) );
  XNOR2_X1 U520 ( .A(n590), .B(n589), .ZN(n615) );
  AND2_X1 U521 ( .A1(G227), .A2(n779), .ZN(n348) );
  AND2_X1 U522 ( .A1(n482), .A2(n724), .ZN(n349) );
  AND2_X1 U523 ( .A1(n385), .A2(n580), .ZN(n350) );
  INV_X1 U524 ( .A(G902), .ZN(n484) );
  XOR2_X1 U525 ( .A(KEYINPUT85), .B(KEYINPUT36), .Z(n351) );
  NOR2_X1 U526 ( .A1(n739), .A2(n358), .ZN(n352) );
  XOR2_X1 U527 ( .A(n750), .B(n749), .Z(n353) );
  XNOR2_X1 U528 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n354) );
  INV_X1 U529 ( .A(KEYINPUT2), .ZN(n455) );
  INV_X1 U530 ( .A(KEYINPUT44), .ZN(n497) );
  XNOR2_X2 U531 ( .A(n414), .B(KEYINPUT45), .ZN(n355) );
  BUF_X1 U532 ( .A(n725), .Z(n356) );
  XNOR2_X1 U533 ( .A(n456), .B(n419), .ZN(n780) );
  OR2_X2 U534 ( .A1(n377), .A2(n591), .ZN(n578) );
  XNOR2_X1 U535 ( .A(n544), .B(n543), .ZN(n377) );
  NOR2_X2 U536 ( .A1(n625), .A2(n633), .ZN(n638) );
  NAND2_X1 U537 ( .A1(n355), .A2(n456), .ZN(n357) );
  BUF_X1 U538 ( .A(n377), .Z(n358) );
  NAND2_X1 U539 ( .A1(n389), .A2(n388), .ZN(n359) );
  NAND2_X1 U540 ( .A1(n389), .A2(n388), .ZN(n438) );
  XNOR2_X1 U541 ( .A(n661), .B(n660), .ZN(n662) );
  INV_X1 U542 ( .A(n607), .ZN(n360) );
  BUF_X1 U543 ( .A(n747), .Z(n753) );
  NAND2_X1 U544 ( .A1(n438), .A2(n699), .ZN(n390) );
  XNOR2_X1 U545 ( .A(n521), .B(n362), .ZN(n361) );
  NOR2_X1 U546 ( .A1(n398), .A2(n367), .ZN(n706) );
  NAND2_X1 U547 ( .A1(n355), .A2(n779), .ZN(n761) );
  NOR2_X1 U548 ( .A1(n368), .A2(n697), .ZN(n698) );
  NOR2_X1 U549 ( .A1(n368), .A2(n692), .ZN(n694) );
  XNOR2_X2 U550 ( .A(n376), .B(n523), .ZN(n444) );
  XNOR2_X1 U551 ( .A(n376), .B(n386), .ZN(n661) );
  XNOR2_X2 U552 ( .A(n770), .B(G101), .ZN(n376) );
  NOR2_X1 U553 ( .A1(n723), .A2(n358), .ZN(n734) );
  INV_X1 U554 ( .A(n703), .ZN(n382) );
  NAND2_X1 U555 ( .A1(n383), .A2(n713), .ZN(n681) );
  NAND2_X1 U556 ( .A1(n638), .A2(n639), .ZN(n384) );
  INV_X1 U557 ( .A(n394), .ZN(n385) );
  NAND2_X1 U558 ( .A1(n422), .A2(n421), .ZN(n388) );
  NAND2_X1 U559 ( .A1(n674), .A2(n556), .ZN(n538) );
  NAND2_X1 U560 ( .A1(n402), .A2(n399), .ZN(n409) );
  XNOR2_X1 U561 ( .A(n611), .B(n610), .ZN(n490) );
  XNOR2_X2 U562 ( .A(n441), .B(n420), .ZN(n456) );
  NAND2_X1 U563 ( .A1(n394), .A2(KEYINPUT39), .ZN(n423) );
  NAND2_X1 U564 ( .A1(n607), .A2(n351), .ZN(n405) );
  NAND2_X1 U565 ( .A1(n345), .A2(KEYINPUT44), .ZN(n417) );
  INV_X1 U566 ( .A(n425), .ZN(n422) );
  NAND2_X1 U567 ( .A1(n425), .A2(KEYINPUT39), .ZN(n424) );
  NAND2_X1 U568 ( .A1(n640), .A2(n426), .ZN(n641) );
  NAND2_X1 U569 ( .A1(n576), .A2(n426), .ZN(n591) );
  INV_X1 U570 ( .A(n431), .ZN(n427) );
  NAND2_X1 U571 ( .A1(n429), .A2(n428), .ZN(n464) );
  NOR2_X1 U572 ( .A1(n431), .A2(KEYINPUT44), .ZN(n428) );
  INV_X1 U573 ( .A(n784), .ZN(n430) );
  NAND2_X1 U574 ( .A1(n784), .A2(n630), .ZN(n432) );
  NAND2_X1 U575 ( .A1(n690), .A2(n630), .ZN(n433) );
  NAND2_X1 U576 ( .A1(n631), .A2(n721), .ZN(n435) );
  XNOR2_X1 U577 ( .A(n437), .B(n436), .ZN(n721) );
  INV_X1 U578 ( .A(KEYINPUT97), .ZN(n436) );
  NOR2_X1 U579 ( .A1(n644), .A2(n643), .ZN(n437) );
  NAND2_X1 U580 ( .A1(n359), .A2(n702), .ZN(n657) );
  NAND2_X1 U581 ( .A1(n356), .A2(n724), .ZN(n440) );
  NOR2_X1 U582 ( .A1(n727), .A2(n581), .ZN(n439) );
  NOR2_X1 U583 ( .A1(n728), .A2(n440), .ZN(n729) );
  NOR2_X1 U584 ( .A1(n349), .A2(KEYINPUT30), .ZN(n480) );
  NAND2_X1 U585 ( .A1(n453), .A2(n451), .ZN(n450) );
  NAND2_X1 U586 ( .A1(n490), .A2(n657), .ZN(n441) );
  NAND2_X1 U587 ( .A1(n447), .A2(n446), .ZN(n445) );
  INV_X1 U588 ( .A(n598), .ZN(n586) );
  NAND2_X2 U589 ( .A1(n443), .A2(n450), .ZN(n747) );
  NAND2_X1 U590 ( .A1(n357), .A2(n448), .ZN(n447) );
  XNOR2_X1 U591 ( .A(n444), .B(n489), .ZN(n748) );
  AND2_X1 U592 ( .A1(n648), .A2(n649), .ZN(n452) );
  INV_X1 U593 ( .A(n615), .ZN(n457) );
  NAND2_X1 U594 ( .A1(n631), .A2(n618), .ZN(n620) );
  INV_X1 U595 ( .A(n616), .ZN(n462) );
  NAND2_X1 U596 ( .A1(n615), .A2(n616), .ZN(n463) );
  XNOR2_X2 U597 ( .A(n629), .B(KEYINPUT32), .ZN(n784) );
  XNOR2_X1 U598 ( .A(n473), .B(n571), .ZN(n472) );
  INV_X1 U599 ( .A(G131), .ZN(n474) );
  NAND2_X1 U600 ( .A1(n478), .A2(n475), .ZN(n582) );
  NAND2_X1 U601 ( .A1(n486), .A2(n476), .ZN(n475) );
  AND2_X1 U602 ( .A1(n482), .A2(n477), .ZN(n476) );
  INV_X1 U603 ( .A(n574), .ZN(n485) );
  NAND2_X1 U604 ( .A1(n661), .A2(n574), .ZN(n488) );
  BUF_X1 U605 ( .A(n586), .Z(n607) );
  XNOR2_X2 U606 ( .A(n578), .B(n577), .ZN(n785) );
  INV_X1 U607 ( .A(KEYINPUT84), .ZN(n630) );
  XNOR2_X1 U608 ( .A(KEYINPUT87), .B(KEYINPUT0), .ZN(n616) );
  XNOR2_X1 U609 ( .A(n504), .B(n503), .ZN(n505) );
  INV_X1 U610 ( .A(KEYINPUT109), .ZN(n542) );
  BUF_X1 U611 ( .A(n674), .Z(n676) );
  INV_X1 U612 ( .A(n639), .ZN(n626) );
  NOR2_X1 U613 ( .A1(n593), .A2(n592), .ZN(n702) );
  INV_X1 U614 ( .A(KEYINPUT123), .ZN(n655) );
  XNOR2_X1 U615 ( .A(KEYINPUT13), .B(G475), .ZN(n513) );
  XNOR2_X1 U616 ( .A(G113), .B(G122), .ZN(n504) );
  XNOR2_X1 U617 ( .A(n507), .B(n506), .ZN(n510) );
  XNOR2_X1 U618 ( .A(KEYINPUT72), .B(n508), .ZN(n569) );
  NAND2_X1 U619 ( .A1(n569), .A2(G214), .ZN(n509) );
  XOR2_X1 U620 ( .A(n510), .B(n509), .Z(n511) );
  NOR2_X1 U621 ( .A1(G902), .A2(n669), .ZN(n512) );
  XNOR2_X1 U622 ( .A(n513), .B(n512), .ZN(n596) );
  NAND2_X1 U623 ( .A1(G234), .A2(n779), .ZN(n514) );
  XNOR2_X1 U624 ( .A(G116), .B(G122), .ZN(n516) );
  XNOR2_X2 U625 ( .A(G143), .B(KEYINPUT76), .ZN(n518) );
  INV_X1 U626 ( .A(G128), .ZN(n517) );
  XNOR2_X2 U627 ( .A(n518), .B(n517), .ZN(n521) );
  NAND2_X1 U628 ( .A1(n650), .A2(n484), .ZN(n519) );
  XNOR2_X1 U629 ( .A(n519), .B(G478), .ZN(n595) );
  NOR2_X1 U630 ( .A1(n596), .A2(n595), .ZN(n520) );
  XNOR2_X1 U631 ( .A(n520), .B(KEYINPUT101), .ZN(n727) );
  XNOR2_X2 U632 ( .A(n521), .B(KEYINPUT4), .ZN(n770) );
  XOR2_X1 U633 ( .A(G104), .B(G107), .Z(n522) );
  XNOR2_X1 U634 ( .A(G110), .B(n522), .ZN(n763) );
  XNOR2_X1 U635 ( .A(n763), .B(KEYINPUT68), .ZN(n523) );
  XOR2_X1 U636 ( .A(n524), .B(KEYINPUT88), .Z(n526) );
  INV_X1 U637 ( .A(G119), .ZN(n527) );
  XOR2_X1 U638 ( .A(G116), .B(G113), .Z(n529) );
  XOR2_X1 U639 ( .A(KEYINPUT17), .B(KEYINPUT73), .Z(n532) );
  XNOR2_X1 U640 ( .A(KEYINPUT75), .B(KEYINPUT74), .ZN(n531) );
  XNOR2_X1 U641 ( .A(n532), .B(n531), .ZN(n533) );
  INV_X1 U642 ( .A(n648), .ZN(n556) );
  XOR2_X1 U643 ( .A(KEYINPUT91), .B(KEYINPUT77), .Z(n537) );
  NAND2_X1 U644 ( .A1(n484), .A2(n535), .ZN(n541) );
  NAND2_X1 U645 ( .A1(G210), .A2(n541), .ZN(n536) );
  XNOR2_X2 U646 ( .A(n538), .B(n347), .ZN(n598) );
  INV_X1 U647 ( .A(KEYINPUT71), .ZN(n539) );
  XNOR2_X1 U648 ( .A(n539), .B(KEYINPUT38), .ZN(n540) );
  NAND2_X1 U649 ( .A1(n541), .A2(G214), .ZN(n724) );
  XNOR2_X1 U650 ( .A(n554), .B(n348), .ZN(n545) );
  NOR2_X1 U651 ( .A1(n748), .A2(G902), .ZN(n547) );
  INV_X1 U652 ( .A(G469), .ZN(n546) );
  XNOR2_X1 U653 ( .A(G128), .B(G119), .ZN(n548) );
  XNOR2_X1 U654 ( .A(KEYINPUT93), .B(KEYINPUT23), .ZN(n549) );
  NAND2_X1 U655 ( .A1(G221), .A2(n550), .ZN(n551) );
  XNOR2_X1 U656 ( .A(n552), .B(n551), .ZN(n555) );
  XOR2_X1 U657 ( .A(n554), .B(n553), .Z(n771) );
  XNOR2_X1 U658 ( .A(n555), .B(n771), .ZN(n754) );
  NOR2_X1 U659 ( .A1(n754), .A2(G902), .ZN(n559) );
  NAND2_X1 U660 ( .A1(G234), .A2(n556), .ZN(n557) );
  XNOR2_X1 U661 ( .A(KEYINPUT20), .B(n557), .ZN(n566) );
  NAND2_X1 U662 ( .A1(n566), .A2(G217), .ZN(n558) );
  NAND2_X1 U663 ( .A1(G234), .A2(G237), .ZN(n560) );
  XNOR2_X1 U664 ( .A(n560), .B(KEYINPUT14), .ZN(n561) );
  XNOR2_X1 U665 ( .A(KEYINPUT70), .B(n561), .ZN(n563) );
  AND2_X1 U666 ( .A1(n563), .A2(G953), .ZN(n562) );
  NAND2_X1 U667 ( .A1(G902), .A2(n562), .ZN(n612) );
  OR2_X1 U668 ( .A1(n612), .A2(G900), .ZN(n565) );
  NAND2_X1 U669 ( .A1(G952), .A2(n563), .ZN(n737) );
  NOR2_X1 U670 ( .A1(n737), .A2(G953), .ZN(n614) );
  INV_X1 U671 ( .A(n614), .ZN(n564) );
  AND2_X1 U672 ( .A1(n565), .A2(n564), .ZN(n579) );
  NAND2_X1 U673 ( .A1(n566), .A2(G221), .ZN(n567) );
  XOR2_X1 U674 ( .A(KEYINPUT21), .B(n567), .Z(n712) );
  INV_X1 U675 ( .A(n712), .ZN(n617) );
  NOR2_X1 U676 ( .A1(n579), .A2(n617), .ZN(n568) );
  NAND2_X1 U677 ( .A1(n624), .A2(n568), .ZN(n588) );
  XNOR2_X1 U678 ( .A(KEYINPUT5), .B(G137), .ZN(n570) );
  XNOR2_X1 U679 ( .A(n570), .B(KEYINPUT95), .ZN(n571) );
  INV_X1 U680 ( .A(KEYINPUT96), .ZN(n573) );
  XNOR2_X1 U681 ( .A(n573), .B(G472), .ZN(n574) );
  XNOR2_X1 U682 ( .A(n575), .B(KEYINPUT28), .ZN(n576) );
  INV_X1 U683 ( .A(KEYINPUT42), .ZN(n577) );
  NOR2_X1 U684 ( .A1(n709), .A2(n579), .ZN(n580) );
  INV_X1 U685 ( .A(n724), .ZN(n581) );
  INV_X1 U686 ( .A(KEYINPUT99), .ZN(n583) );
  XNOR2_X1 U687 ( .A(n596), .B(n583), .ZN(n593) );
  INV_X1 U688 ( .A(n595), .ZN(n592) );
  XOR2_X1 U689 ( .A(KEYINPUT108), .B(KEYINPUT40), .Z(n584) );
  XNOR2_X1 U690 ( .A(n585), .B(n354), .ZN(n601) );
  INV_X1 U691 ( .A(KEYINPUT6), .ZN(n587) );
  INV_X1 U692 ( .A(n633), .ZN(n710) );
  NAND2_X1 U693 ( .A1(n598), .A2(n724), .ZN(n590) );
  NOR2_X1 U694 ( .A1(n699), .A2(n702), .ZN(n728) );
  NAND2_X1 U695 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U696 ( .A(n597), .B(KEYINPUT105), .ZN(n637) );
  AND2_X1 U697 ( .A1(n360), .A2(n637), .ZN(n599) );
  AND2_X1 U698 ( .A1(n599), .A2(n350), .ZN(n695) );
  NAND2_X1 U699 ( .A1(n601), .A2(n600), .ZN(n603) );
  INV_X1 U700 ( .A(KEYINPUT48), .ZN(n602) );
  XNOR2_X1 U701 ( .A(n603), .B(n602), .ZN(n609) );
  XNOR2_X1 U702 ( .A(KEYINPUT107), .B(n604), .ZN(n605) );
  NAND2_X1 U703 ( .A1(n605), .A2(n710), .ZN(n606) );
  XNOR2_X1 U704 ( .A(n606), .B(KEYINPUT43), .ZN(n608) );
  NAND2_X1 U705 ( .A1(n608), .A2(n607), .ZN(n708) );
  NAND2_X1 U706 ( .A1(n609), .A2(n708), .ZN(n611) );
  INV_X1 U707 ( .A(KEYINPUT82), .ZN(n610) );
  INV_X1 U708 ( .A(KEYINPUT103), .ZN(n621) );
  NOR2_X1 U709 ( .A1(G898), .A2(n612), .ZN(n613) );
  NOR2_X1 U710 ( .A1(n727), .A2(n617), .ZN(n618) );
  AND2_X1 U711 ( .A1(n624), .A2(n643), .ZN(n622) );
  XOR2_X1 U712 ( .A(KEYINPUT102), .B(n624), .Z(n713) );
  INV_X1 U713 ( .A(n631), .ZN(n642) );
  INV_X1 U714 ( .A(n709), .ZN(n632) );
  NAND2_X1 U715 ( .A1(n633), .A2(n632), .ZN(n644) );
  NOR2_X1 U716 ( .A1(n644), .A2(n639), .ZN(n635) );
  XNOR2_X1 U717 ( .A(KEYINPUT104), .B(KEYINPUT33), .ZN(n634) );
  XNOR2_X1 U718 ( .A(n635), .B(n634), .ZN(n739) );
  NOR2_X1 U719 ( .A1(n642), .A2(n739), .ZN(n636) );
  INV_X1 U720 ( .A(n643), .ZN(n718) );
  NOR2_X1 U721 ( .A1(n709), .A2(n718), .ZN(n640) );
  NOR2_X1 U722 ( .A1(n642), .A2(n641), .ZN(n687) );
  NAND2_X1 U723 ( .A1(n657), .A2(KEYINPUT2), .ZN(n645) );
  XOR2_X1 U724 ( .A(KEYINPUT78), .B(n645), .Z(n646) );
  INV_X1 U725 ( .A(KEYINPUT65), .ZN(n649) );
  NAND2_X1 U726 ( .A1(n747), .A2(G478), .ZN(n652) );
  XNOR2_X1 U727 ( .A(n652), .B(n651), .ZN(n654) );
  INV_X1 U728 ( .A(G952), .ZN(n653) );
  AND2_X1 U729 ( .A1(n653), .A2(G953), .ZN(n757) );
  XNOR2_X1 U730 ( .A(n656), .B(n655), .ZN(G63) );
  XNOR2_X1 U731 ( .A(n657), .B(G134), .ZN(G36) );
  XOR2_X1 U732 ( .A(n658), .B(G131), .Z(G33) );
  NAND2_X1 U733 ( .A1(n747), .A2(G472), .ZN(n663) );
  XOR2_X1 U734 ( .A(KEYINPUT89), .B(KEYINPUT110), .Z(n659) );
  XNOR2_X1 U735 ( .A(n659), .B(KEYINPUT62), .ZN(n660) );
  XNOR2_X1 U736 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U737 ( .A(KEYINPUT90), .B(KEYINPUT63), .ZN(n665) );
  XOR2_X1 U738 ( .A(n665), .B(KEYINPUT86), .Z(n666) );
  XNOR2_X1 U739 ( .A(n667), .B(n666), .ZN(G57) );
  NAND2_X1 U740 ( .A1(n747), .A2(G475), .ZN(n671) );
  XOR2_X1 U741 ( .A(KEYINPUT66), .B(KEYINPUT59), .Z(n668) );
  XNOR2_X1 U742 ( .A(n671), .B(n670), .ZN(n672) );
  XNOR2_X1 U743 ( .A(n673), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U744 ( .A1(n747), .A2(G210), .ZN(n678) );
  XNOR2_X1 U745 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n675) );
  XNOR2_X1 U746 ( .A(n678), .B(n677), .ZN(n679) );
  XNOR2_X1 U747 ( .A(n680), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U748 ( .A(G101), .B(n681), .ZN(G3) );
  XOR2_X1 U749 ( .A(G104), .B(KEYINPUT111), .Z(n683) );
  NAND2_X1 U750 ( .A1(n687), .A2(n699), .ZN(n682) );
  XNOR2_X1 U751 ( .A(n683), .B(n682), .ZN(G6) );
  XOR2_X1 U752 ( .A(KEYINPUT27), .B(KEYINPUT113), .Z(n685) );
  XNOR2_X1 U753 ( .A(G107), .B(KEYINPUT112), .ZN(n684) );
  XNOR2_X1 U754 ( .A(n685), .B(n684), .ZN(n686) );
  XOR2_X1 U755 ( .A(KEYINPUT26), .B(n686), .Z(n689) );
  NAND2_X1 U756 ( .A1(n687), .A2(n702), .ZN(n688) );
  XNOR2_X1 U757 ( .A(n689), .B(n688), .ZN(G9) );
  XOR2_X1 U758 ( .A(n690), .B(G110), .Z(n691) );
  XNOR2_X1 U759 ( .A(KEYINPUT114), .B(n691), .ZN(G12) );
  INV_X1 U760 ( .A(n702), .ZN(n692) );
  XNOR2_X1 U761 ( .A(G128), .B(KEYINPUT29), .ZN(n693) );
  XNOR2_X1 U762 ( .A(n694), .B(n693), .ZN(G30) );
  XNOR2_X1 U763 ( .A(G143), .B(n695), .ZN(n696) );
  XNOR2_X1 U764 ( .A(n696), .B(KEYINPUT115), .ZN(G45) );
  XOR2_X1 U765 ( .A(G146), .B(n698), .Z(G48) );
  NAND2_X1 U766 ( .A1(n703), .A2(n699), .ZN(n700) );
  XNOR2_X1 U767 ( .A(n700), .B(KEYINPUT116), .ZN(n701) );
  XNOR2_X1 U768 ( .A(G113), .B(n701), .ZN(G15) );
  XOR2_X1 U769 ( .A(G116), .B(KEYINPUT117), .Z(n705) );
  NAND2_X1 U770 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U771 ( .A(n705), .B(n704), .ZN(G18) );
  XNOR2_X1 U772 ( .A(G125), .B(n706), .ZN(n707) );
  XNOR2_X1 U773 ( .A(n707), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U774 ( .A(G140), .B(n708), .ZN(G42) );
  NAND2_X1 U775 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U776 ( .A(KEYINPUT50), .B(n711), .ZN(n717) );
  NOR2_X1 U777 ( .A1(n713), .A2(n712), .ZN(n715) );
  XNOR2_X1 U778 ( .A(KEYINPUT118), .B(KEYINPUT49), .ZN(n714) );
  XNOR2_X1 U779 ( .A(n715), .B(n714), .ZN(n716) );
  NAND2_X1 U780 ( .A1(n717), .A2(n716), .ZN(n719) );
  NOR2_X1 U781 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U782 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U783 ( .A(KEYINPUT51), .B(n722), .Z(n723) );
  NOR2_X1 U784 ( .A1(n356), .A2(n724), .ZN(n726) );
  NOR2_X1 U785 ( .A1(n727), .A2(n726), .ZN(n731) );
  XOR2_X1 U786 ( .A(KEYINPUT119), .B(n729), .Z(n730) );
  NOR2_X1 U787 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U788 ( .A1(n739), .A2(n732), .ZN(n733) );
  NOR2_X1 U789 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U790 ( .A(n735), .B(KEYINPUT52), .ZN(n736) );
  NOR2_X1 U791 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U792 ( .A(n738), .B(KEYINPUT120), .ZN(n740) );
  NOR2_X1 U793 ( .A1(n740), .A2(n352), .ZN(n741) );
  NAND2_X1 U794 ( .A1(n741), .A2(n779), .ZN(n745) );
  XNOR2_X1 U795 ( .A(n742), .B(KEYINPUT79), .ZN(n743) );
  NOR2_X1 U796 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U797 ( .A(n746), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U798 ( .A1(n753), .A2(G469), .ZN(n751) );
  XOR2_X1 U799 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n750) );
  XNOR2_X1 U800 ( .A(n748), .B(KEYINPUT121), .ZN(n749) );
  NOR2_X1 U801 ( .A1(n757), .A2(n752), .ZN(G54) );
  NAND2_X1 U802 ( .A1(n753), .A2(G217), .ZN(n755) );
  XNOR2_X1 U803 ( .A(n755), .B(n754), .ZN(n756) );
  NOR2_X1 U804 ( .A1(n757), .A2(n756), .ZN(G66) );
  NAND2_X1 U805 ( .A1(G953), .A2(G224), .ZN(n758) );
  XNOR2_X1 U806 ( .A(KEYINPUT61), .B(n758), .ZN(n759) );
  NAND2_X1 U807 ( .A1(n759), .A2(G898), .ZN(n760) );
  NAND2_X1 U808 ( .A1(n761), .A2(n760), .ZN(n768) );
  XNOR2_X1 U809 ( .A(G101), .B(n762), .ZN(n764) );
  XNOR2_X1 U810 ( .A(n764), .B(n763), .ZN(n766) );
  NOR2_X1 U811 ( .A1(G898), .A2(n779), .ZN(n765) );
  NOR2_X1 U812 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U813 ( .A(n768), .B(n767), .ZN(n769) );
  XNOR2_X1 U814 ( .A(KEYINPUT124), .B(n769), .ZN(G69) );
  XOR2_X1 U815 ( .A(n772), .B(n771), .Z(n773) );
  XNOR2_X1 U816 ( .A(KEYINPUT125), .B(n773), .ZN(n774) );
  XOR2_X1 U817 ( .A(n770), .B(n774), .Z(n778) );
  XNOR2_X1 U818 ( .A(n778), .B(G227), .ZN(n775) );
  NAND2_X1 U819 ( .A1(n775), .A2(G900), .ZN(n776) );
  NAND2_X1 U820 ( .A1(G953), .A2(n776), .ZN(n777) );
  XNOR2_X1 U821 ( .A(n777), .B(KEYINPUT126), .ZN(n782) );
  NAND2_X1 U822 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U823 ( .A1(n782), .A2(n781), .ZN(G72) );
  XNOR2_X1 U824 ( .A(n345), .B(G122), .ZN(n783) );
  XNOR2_X1 U825 ( .A(n783), .B(KEYINPUT127), .ZN(G24) );
  XOR2_X1 U826 ( .A(n784), .B(G119), .Z(G21) );
  XOR2_X1 U827 ( .A(n785), .B(G137), .Z(G39) );
endmodule

