

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585;

  XOR2_X1 U323 ( .A(n345), .B(n453), .Z(n520) );
  XNOR2_X1 U324 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U325 ( .A(n374), .B(n373), .Z(n291) );
  INV_X1 U326 ( .A(KEYINPUT54), .ZN(n432) );
  XNOR2_X1 U327 ( .A(G169GAT), .B(G36GAT), .ZN(n331) );
  XNOR2_X1 U328 ( .A(n432), .B(KEYINPUT119), .ZN(n433) );
  XNOR2_X1 U329 ( .A(n375), .B(n291), .ZN(n376) );
  XNOR2_X1 U330 ( .A(n377), .B(n376), .ZN(n379) );
  NOR2_X1 U331 ( .A1(n516), .A2(n515), .ZN(n517) );
  XOR2_X1 U332 ( .A(n313), .B(n312), .Z(n532) );
  XOR2_X1 U333 ( .A(KEYINPUT28), .B(n474), .Z(n534) );
  XNOR2_X1 U334 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n458) );
  XNOR2_X1 U335 ( .A(n459), .B(n458), .ZN(G1351GAT) );
  XOR2_X1 U336 ( .A(KEYINPUT0), .B(KEYINPUT82), .Z(n293) );
  XNOR2_X1 U337 ( .A(KEYINPUT81), .B(G127GAT), .ZN(n292) );
  XNOR2_X1 U338 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U339 ( .A(G113GAT), .B(n294), .Z(n330) );
  NAND2_X1 U340 ( .A1(G227GAT), .A2(G233GAT), .ZN(n300) );
  XOR2_X1 U341 ( .A(KEYINPUT85), .B(KEYINPUT20), .Z(n296) );
  XNOR2_X1 U342 ( .A(G99GAT), .B(KEYINPUT84), .ZN(n295) );
  XNOR2_X1 U343 ( .A(n296), .B(n295), .ZN(n298) );
  XOR2_X1 U344 ( .A(G43GAT), .B(G134GAT), .Z(n297) );
  XNOR2_X1 U345 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U346 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U347 ( .A(n330), .B(n301), .ZN(n313) );
  XOR2_X1 U348 ( .A(KEYINPUT18), .B(G190GAT), .Z(n303) );
  XNOR2_X1 U349 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n302) );
  XNOR2_X1 U350 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U351 ( .A(KEYINPUT19), .B(n304), .Z(n341) );
  XOR2_X1 U352 ( .A(KEYINPUT86), .B(KEYINPUT87), .Z(n306) );
  XNOR2_X1 U353 ( .A(G120GAT), .B(G176GAT), .ZN(n305) );
  XNOR2_X1 U354 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U355 ( .A(n341), .B(n307), .ZN(n311) );
  XOR2_X1 U356 ( .A(G71GAT), .B(KEYINPUT83), .Z(n309) );
  XNOR2_X1 U357 ( .A(G169GAT), .B(G15GAT), .ZN(n308) );
  XNOR2_X1 U358 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U359 ( .A(n311), .B(n310), .ZN(n312) );
  INV_X1 U360 ( .A(n532), .ZN(n475) );
  XNOR2_X1 U361 ( .A(G29GAT), .B(G85GAT), .ZN(n314) );
  XOR2_X1 U362 ( .A(G120GAT), .B(G57GAT), .Z(n365) );
  XNOR2_X1 U363 ( .A(n314), .B(n365), .ZN(n318) );
  XOR2_X1 U364 ( .A(KEYINPUT94), .B(G148GAT), .Z(n316) );
  XNOR2_X1 U365 ( .A(G1GAT), .B(G141GAT), .ZN(n315) );
  XNOR2_X1 U366 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U367 ( .A(n318), .B(n317), .Z(n328) );
  XOR2_X1 U368 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n320) );
  XNOR2_X1 U369 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n319) );
  XNOR2_X1 U370 ( .A(n320), .B(n319), .ZN(n326) );
  XOR2_X1 U371 ( .A(G134GAT), .B(KEYINPUT76), .Z(n409) );
  XOR2_X1 U372 ( .A(G155GAT), .B(KEYINPUT2), .Z(n322) );
  XNOR2_X1 U373 ( .A(G162GAT), .B(KEYINPUT3), .ZN(n321) );
  XNOR2_X1 U374 ( .A(n322), .B(n321), .ZN(n442) );
  XOR2_X1 U375 ( .A(n409), .B(n442), .Z(n324) );
  NAND2_X1 U376 ( .A1(G225GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U377 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U378 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U379 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U380 ( .A(n330), .B(n329), .Z(n472) );
  INV_X1 U381 ( .A(n472), .ZN(n518) );
  XNOR2_X1 U382 ( .A(n331), .B(G8GAT), .ZN(n380) );
  XNOR2_X1 U383 ( .A(n380), .B(KEYINPUT97), .ZN(n333) );
  XOR2_X1 U384 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n332) );
  XNOR2_X1 U385 ( .A(n333), .B(n332), .ZN(n337) );
  XOR2_X1 U386 ( .A(KEYINPUT75), .B(G64GAT), .Z(n335) );
  XNOR2_X1 U387 ( .A(G176GAT), .B(G92GAT), .ZN(n334) );
  XNOR2_X1 U388 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U389 ( .A(G204GAT), .B(n336), .ZN(n378) );
  XNOR2_X1 U390 ( .A(n337), .B(n378), .ZN(n339) );
  NAND2_X1 U391 ( .A1(G226GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U392 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U393 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U394 ( .A(KEYINPUT21), .B(G218GAT), .Z(n343) );
  XNOR2_X1 U395 ( .A(KEYINPUT90), .B(G211GAT), .ZN(n342) );
  XNOR2_X1 U396 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U397 ( .A(G197GAT), .B(n344), .Z(n453) );
  XNOR2_X1 U398 ( .A(n520), .B(KEYINPUT118), .ZN(n431) );
  XNOR2_X1 U399 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n430) );
  XOR2_X1 U400 ( .A(G57GAT), .B(G155GAT), .Z(n347) );
  XNOR2_X1 U401 ( .A(G8GAT), .B(G211GAT), .ZN(n346) );
  XNOR2_X1 U402 ( .A(n347), .B(n346), .ZN(n351) );
  XOR2_X1 U403 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n349) );
  XNOR2_X1 U404 ( .A(G64GAT), .B(KEYINPUT78), .ZN(n348) );
  XNOR2_X1 U405 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U406 ( .A(n351), .B(n350), .ZN(n362) );
  XNOR2_X1 U407 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n352) );
  XNOR2_X1 U408 ( .A(n352), .B(KEYINPUT72), .ZN(n364) );
  XOR2_X1 U409 ( .A(n364), .B(G78GAT), .Z(n354) );
  XNOR2_X1 U410 ( .A(G127GAT), .B(G183GAT), .ZN(n353) );
  XNOR2_X1 U411 ( .A(n354), .B(n353), .ZN(n360) );
  XNOR2_X1 U412 ( .A(G15GAT), .B(G1GAT), .ZN(n355) );
  XNOR2_X1 U413 ( .A(n355), .B(KEYINPUT70), .ZN(n383) );
  XOR2_X1 U414 ( .A(KEYINPUT12), .B(n383), .Z(n357) );
  NAND2_X1 U415 ( .A1(G231GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U416 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U417 ( .A(G22GAT), .B(n358), .Z(n359) );
  XNOR2_X1 U418 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U419 ( .A(n362), .B(n361), .Z(n551) );
  INV_X1 U420 ( .A(n551), .ZN(n578) );
  XOR2_X1 U421 ( .A(KEYINPUT46), .B(KEYINPUT111), .Z(n398) );
  INV_X1 U422 ( .A(n365), .ZN(n363) );
  NAND2_X1 U423 ( .A1(n364), .A2(n363), .ZN(n368) );
  INV_X1 U424 ( .A(n364), .ZN(n366) );
  NAND2_X1 U425 ( .A1(n366), .A2(n365), .ZN(n367) );
  NAND2_X1 U426 ( .A1(n368), .A2(n367), .ZN(n370) );
  NAND2_X1 U427 ( .A1(G230GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U428 ( .A(n370), .B(n369), .ZN(n377) );
  XNOR2_X1 U429 ( .A(G106GAT), .B(G78GAT), .ZN(n371) );
  XNOR2_X1 U430 ( .A(n371), .B(G148GAT), .ZN(n447) );
  XNOR2_X1 U431 ( .A(G99GAT), .B(G85GAT), .ZN(n372) );
  XNOR2_X1 U432 ( .A(n372), .B(KEYINPUT74), .ZN(n408) );
  XNOR2_X1 U433 ( .A(n447), .B(n408), .ZN(n375) );
  XOR2_X1 U434 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n374) );
  XNOR2_X1 U435 ( .A(KEYINPUT73), .B(KEYINPUT32), .ZN(n373) );
  XOR2_X1 U436 ( .A(n379), .B(n378), .Z(n575) );
  XNOR2_X1 U437 ( .A(n575), .B(KEYINPUT41), .ZN(n501) );
  INV_X1 U438 ( .A(n501), .ZN(n396) );
  XOR2_X1 U439 ( .A(n380), .B(G197GAT), .Z(n382) );
  XOR2_X1 U440 ( .A(G141GAT), .B(G22GAT), .Z(n443) );
  XNOR2_X1 U441 ( .A(G113GAT), .B(n443), .ZN(n381) );
  XNOR2_X1 U442 ( .A(n382), .B(n381), .ZN(n387) );
  XOR2_X1 U443 ( .A(n383), .B(KEYINPUT68), .Z(n385) );
  NAND2_X1 U444 ( .A1(G229GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U445 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U446 ( .A(n387), .B(n386), .Z(n395) );
  XOR2_X1 U447 ( .A(KEYINPUT7), .B(G50GAT), .Z(n389) );
  XNOR2_X1 U448 ( .A(G43GAT), .B(G29GAT), .ZN(n388) );
  XNOR2_X1 U449 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U450 ( .A(KEYINPUT8), .B(n390), .Z(n413) );
  XOR2_X1 U451 ( .A(KEYINPUT69), .B(KEYINPUT30), .Z(n392) );
  XNOR2_X1 U452 ( .A(KEYINPUT29), .B(KEYINPUT67), .ZN(n391) );
  XNOR2_X1 U453 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U454 ( .A(n413), .B(n393), .ZN(n394) );
  XOR2_X1 U455 ( .A(n395), .B(n394), .Z(n546) );
  INV_X1 U456 ( .A(n546), .ZN(n572) );
  NAND2_X1 U457 ( .A1(n396), .A2(n572), .ZN(n397) );
  XOR2_X1 U458 ( .A(n398), .B(n397), .Z(n399) );
  NOR2_X1 U459 ( .A1(n578), .A2(n399), .ZN(n418) );
  XOR2_X1 U460 ( .A(KEYINPUT11), .B(G106GAT), .Z(n401) );
  XNOR2_X1 U461 ( .A(G36GAT), .B(G190GAT), .ZN(n400) );
  XNOR2_X1 U462 ( .A(n401), .B(n400), .ZN(n417) );
  XOR2_X1 U463 ( .A(G92GAT), .B(KEYINPUT77), .Z(n403) );
  XNOR2_X1 U464 ( .A(G218GAT), .B(G162GAT), .ZN(n402) );
  XNOR2_X1 U465 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U466 ( .A(KEYINPUT65), .B(KEYINPUT9), .Z(n405) );
  XNOR2_X1 U467 ( .A(KEYINPUT10), .B(KEYINPUT66), .ZN(n404) );
  XNOR2_X1 U468 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U469 ( .A(n407), .B(n406), .Z(n415) );
  XNOR2_X1 U470 ( .A(n409), .B(n408), .ZN(n411) );
  AND2_X1 U471 ( .A1(G232GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U472 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U473 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U474 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U475 ( .A(n417), .B(n416), .ZN(n541) );
  INV_X1 U476 ( .A(n541), .ZN(n554) );
  NAND2_X1 U477 ( .A1(n418), .A2(n554), .ZN(n420) );
  XOR2_X1 U478 ( .A(KEYINPUT112), .B(KEYINPUT47), .Z(n419) );
  XNOR2_X1 U479 ( .A(n420), .B(n419), .ZN(n428) );
  XOR2_X1 U480 ( .A(KEYINPUT45), .B(KEYINPUT113), .Z(n423) );
  XNOR2_X1 U481 ( .A(KEYINPUT36), .B(KEYINPUT102), .ZN(n421) );
  XOR2_X1 U482 ( .A(n421), .B(n554), .Z(n580) );
  NAND2_X1 U483 ( .A1(n578), .A2(n580), .ZN(n422) );
  XNOR2_X1 U484 ( .A(n423), .B(n422), .ZN(n424) );
  NOR2_X1 U485 ( .A1(n424), .A2(n575), .ZN(n425) );
  XNOR2_X1 U486 ( .A(KEYINPUT114), .B(n425), .ZN(n426) );
  XOR2_X1 U487 ( .A(KEYINPUT71), .B(n546), .Z(n527) );
  NAND2_X1 U488 ( .A1(n426), .A2(n527), .ZN(n427) );
  NAND2_X1 U489 ( .A1(n428), .A2(n427), .ZN(n429) );
  XNOR2_X1 U490 ( .A(n430), .B(n429), .ZN(n529) );
  NAND2_X1 U491 ( .A1(n431), .A2(n529), .ZN(n434) );
  NOR2_X1 U492 ( .A1(n518), .A2(n435), .ZN(n570) );
  XOR2_X1 U493 ( .A(KEYINPUT89), .B(G204GAT), .Z(n437) );
  XNOR2_X1 U494 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n436) );
  XNOR2_X1 U495 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U496 ( .A(KEYINPUT92), .B(KEYINPUT24), .Z(n439) );
  XNOR2_X1 U497 ( .A(G50GAT), .B(KEYINPUT88), .ZN(n438) );
  XNOR2_X1 U498 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U499 ( .A(n441), .B(n440), .ZN(n451) );
  XOR2_X1 U500 ( .A(n443), .B(n442), .Z(n445) );
  NAND2_X1 U501 ( .A1(G228GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U502 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U503 ( .A(n446), .B(KEYINPUT93), .Z(n449) );
  XNOR2_X1 U504 ( .A(n447), .B(KEYINPUT91), .ZN(n448) );
  XNOR2_X1 U505 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U506 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U507 ( .A(n453), .B(n452), .ZN(n474) );
  NAND2_X1 U508 ( .A1(n570), .A2(n474), .ZN(n455) );
  INV_X1 U509 ( .A(KEYINPUT55), .ZN(n454) );
  XNOR2_X1 U510 ( .A(n455), .B(n454), .ZN(n456) );
  NOR2_X1 U511 ( .A1(n475), .A2(n456), .ZN(n457) );
  XNOR2_X1 U512 ( .A(KEYINPUT120), .B(n457), .ZN(n563) );
  NAND2_X1 U513 ( .A1(n563), .A2(n541), .ZN(n459) );
  OR2_X1 U514 ( .A1(n527), .A2(n575), .ZN(n491) );
  NAND2_X1 U515 ( .A1(n578), .A2(n554), .ZN(n462) );
  XNOR2_X1 U516 ( .A(KEYINPUT16), .B(KEYINPUT80), .ZN(n460) );
  XNOR2_X1 U517 ( .A(n460), .B(KEYINPUT79), .ZN(n461) );
  XNOR2_X1 U518 ( .A(n462), .B(n461), .ZN(n479) );
  NAND2_X1 U519 ( .A1(n532), .A2(n520), .ZN(n463) );
  XOR2_X1 U520 ( .A(KEYINPUT99), .B(n463), .Z(n464) );
  NAND2_X1 U521 ( .A1(n474), .A2(n464), .ZN(n465) );
  XOR2_X1 U522 ( .A(KEYINPUT25), .B(n465), .Z(n466) );
  XNOR2_X1 U523 ( .A(n466), .B(KEYINPUT100), .ZN(n470) );
  XNOR2_X1 U524 ( .A(KEYINPUT27), .B(n520), .ZN(n473) );
  NOR2_X1 U525 ( .A1(n532), .A2(n474), .ZN(n468) );
  XNOR2_X1 U526 ( .A(KEYINPUT26), .B(KEYINPUT98), .ZN(n467) );
  XNOR2_X1 U527 ( .A(n468), .B(n467), .ZN(n569) );
  NAND2_X1 U528 ( .A1(n473), .A2(n569), .ZN(n469) );
  NAND2_X1 U529 ( .A1(n470), .A2(n469), .ZN(n471) );
  NAND2_X1 U530 ( .A1(n472), .A2(n471), .ZN(n478) );
  NAND2_X1 U531 ( .A1(n473), .A2(n518), .ZN(n528) );
  NOR2_X1 U532 ( .A1(n528), .A2(n534), .ZN(n476) );
  NAND2_X1 U533 ( .A1(n476), .A2(n475), .ZN(n477) );
  NAND2_X1 U534 ( .A1(n478), .A2(n477), .ZN(n488) );
  NAND2_X1 U535 ( .A1(n479), .A2(n488), .ZN(n502) );
  NOR2_X1 U536 ( .A1(n491), .A2(n502), .ZN(n486) );
  NAND2_X1 U537 ( .A1(n518), .A2(n486), .ZN(n480) );
  XNOR2_X1 U538 ( .A(n480), .B(KEYINPUT34), .ZN(n481) );
  XNOR2_X1 U539 ( .A(G1GAT), .B(n481), .ZN(G1324GAT) );
  NAND2_X1 U540 ( .A1(n520), .A2(n486), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n482), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U542 ( .A(KEYINPUT101), .B(KEYINPUT35), .Z(n484) );
  NAND2_X1 U543 ( .A1(n486), .A2(n532), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n484), .B(n483), .ZN(n485) );
  XOR2_X1 U545 ( .A(G15GAT), .B(n485), .Z(G1326GAT) );
  NAND2_X1 U546 ( .A1(n534), .A2(n486), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n487), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U548 ( .A(G29GAT), .B(KEYINPUT39), .Z(n494) );
  NAND2_X1 U549 ( .A1(n488), .A2(n580), .ZN(n489) );
  NOR2_X1 U550 ( .A1(n489), .A2(n578), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n490), .B(KEYINPUT37), .ZN(n516) );
  NOR2_X1 U552 ( .A1(n491), .A2(n516), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n492), .B(KEYINPUT38), .ZN(n499) );
  NAND2_X1 U554 ( .A1(n499), .A2(n518), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(G1328GAT) );
  XOR2_X1 U556 ( .A(G36GAT), .B(KEYINPUT103), .Z(n496) );
  NAND2_X1 U557 ( .A1(n499), .A2(n520), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(G1329GAT) );
  NAND2_X1 U559 ( .A1(n499), .A2(n532), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n497), .B(KEYINPUT40), .ZN(n498) );
  XNOR2_X1 U561 ( .A(G43GAT), .B(n498), .ZN(G1330GAT) );
  NAND2_X1 U562 ( .A1(n499), .A2(n534), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n500), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U564 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n504) );
  NAND2_X1 U565 ( .A1(n546), .A2(n396), .ZN(n515) );
  NOR2_X1 U566 ( .A1(n515), .A2(n502), .ZN(n512) );
  NAND2_X1 U567 ( .A1(n512), .A2(n518), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n504), .B(n503), .ZN(G1332GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n506) );
  NAND2_X1 U570 ( .A1(n512), .A2(n520), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U572 ( .A(G64GAT), .B(n507), .ZN(G1333GAT) );
  NAND2_X1 U573 ( .A1(n512), .A2(n532), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n508), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U575 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n510) );
  XNOR2_X1 U576 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n509) );
  XNOR2_X1 U577 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U578 ( .A(KEYINPUT106), .B(n511), .Z(n514) );
  NAND2_X1 U579 ( .A1(n512), .A2(n534), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(G1335GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT109), .B(n517), .Z(n523) );
  NAND2_X1 U582 ( .A1(n523), .A2(n518), .ZN(n519) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(n519), .ZN(G1336GAT) );
  NAND2_X1 U584 ( .A1(n520), .A2(n523), .ZN(n521) );
  XNOR2_X1 U585 ( .A(n521), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U586 ( .A1(n523), .A2(n532), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n522), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U588 ( .A1(n523), .A2(n534), .ZN(n525) );
  XOR2_X1 U589 ( .A(KEYINPUT44), .B(KEYINPUT110), .Z(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U591 ( .A(G106GAT), .B(n526), .Z(G1339GAT) );
  INV_X1 U592 ( .A(n527), .ZN(n557) );
  INV_X1 U593 ( .A(n528), .ZN(n530) );
  NAND2_X1 U594 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U595 ( .A(KEYINPUT115), .B(n531), .ZN(n545) );
  NAND2_X1 U596 ( .A1(n532), .A2(n545), .ZN(n533) );
  NOR2_X1 U597 ( .A1(n534), .A2(n533), .ZN(n542) );
  NAND2_X1 U598 ( .A1(n557), .A2(n542), .ZN(n535) );
  XNOR2_X1 U599 ( .A(KEYINPUT116), .B(n535), .ZN(n536) );
  XNOR2_X1 U600 ( .A(G113GAT), .B(n536), .ZN(G1340GAT) );
  XOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT49), .Z(n538) );
  NAND2_X1 U602 ( .A1(n542), .A2(n396), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n538), .B(n537), .ZN(G1341GAT) );
  NAND2_X1 U604 ( .A1(n578), .A2(n542), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n539), .B(KEYINPUT50), .ZN(n540) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n540), .ZN(G1342GAT) );
  XOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT51), .Z(n544) );
  NAND2_X1 U608 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  NAND2_X1 U610 ( .A1(n569), .A2(n545), .ZN(n553) );
  NOR2_X1 U611 ( .A1(n546), .A2(n553), .ZN(n547) );
  XOR2_X1 U612 ( .A(G141GAT), .B(n547), .Z(G1344GAT) );
  NOR2_X1 U613 ( .A1(n501), .A2(n553), .ZN(n549) );
  XNOR2_X1 U614 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(n550), .ZN(G1345GAT) );
  NOR2_X1 U617 ( .A1(n551), .A2(n553), .ZN(n552) );
  XOR2_X1 U618 ( .A(G155GAT), .B(n552), .Z(G1346GAT) );
  NOR2_X1 U619 ( .A1(n554), .A2(n553), .ZN(n556) );
  XNOR2_X1 U620 ( .A(G162GAT), .B(KEYINPUT117), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n556), .B(n555), .ZN(G1347GAT) );
  XOR2_X1 U622 ( .A(G169GAT), .B(KEYINPUT121), .Z(n559) );
  NAND2_X1 U623 ( .A1(n557), .A2(n563), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(G1348GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n561) );
  XNOR2_X1 U626 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U628 ( .A(KEYINPUT122), .B(n562), .Z(n565) );
  NAND2_X1 U629 ( .A1(n563), .A2(n396), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(G1349GAT) );
  NAND2_X1 U631 ( .A1(n563), .A2(n578), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n568) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n574) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U637 ( .A(KEYINPUT124), .B(n571), .Z(n581) );
  NAND2_X1 U638 ( .A1(n581), .A2(n572), .ZN(n573) );
  XOR2_X1 U639 ( .A(n574), .B(n573), .Z(G1352GAT) );
  XOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT61), .Z(n577) );
  NAND2_X1 U641 ( .A1(n581), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NAND2_X1 U643 ( .A1(n581), .A2(n578), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(G211GAT), .ZN(G1354GAT) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n585) );
  XOR2_X1 U646 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n583) );
  NAND2_X1 U647 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(G1355GAT) );
endmodule

