//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0 1 1 0 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 0 1 0 1 1 1 1 0 1 1 1 0 0 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:55 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1208, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  XOR2_X1   g0006(.A(KEYINPUT65), .B(G244), .Z(new_n207));
  AOI22_X1  g0007(.A1(new_n207), .A2(G77), .B1(G116), .B2(G270), .ZN(new_n208));
  INV_X1    g0008(.A(G50), .ZN(new_n209));
  INV_X1    g0009(.A(G226), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  OAI221_X1 g0012(.A(new_n208), .B1(new_n209), .B2(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(KEYINPUT66), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AND2_X1   g0015(.A1(new_n213), .A2(new_n214), .ZN(new_n216));
  AOI211_X1 g0016(.A(new_n215), .B(new_n216), .C1(G87), .C2(G250), .ZN(new_n217));
  INV_X1    g0017(.A(G58), .ZN(new_n218));
  INV_X1    g0018(.A(G232), .ZN(new_n219));
  INV_X1    g0019(.A(G97), .ZN(new_n220));
  INV_X1    g0020(.A(G257), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AND2_X1   g0022(.A1(G107), .A2(G264), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n206), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT1), .Z(new_n225));
  INV_X1    g0025(.A(KEYINPUT64), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n226), .B1(new_n206), .B2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(G13), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n205), .A2(KEYINPUT64), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n230), .B(G250), .C1(G257), .C2(G264), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT0), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n234), .A2(G20), .ZN(new_n235));
  NOR2_X1   g0035(.A1(G58), .A2(G68), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g0037(.A1(new_n237), .A2(G50), .ZN(new_n238));
  OAI211_X1 g0038(.A(new_n225), .B(new_n232), .C1(new_n235), .C2(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n239), .B(KEYINPUT67), .Z(G361));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G264), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n242), .B(G270), .Z(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT2), .B(G226), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n219), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G238), .B(G244), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n243), .B(new_n247), .Z(G358));
  XOR2_X1   g0048(.A(G50), .B(G58), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT68), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G68), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G87), .B(G97), .ZN(new_n253));
  XNOR2_X1  g0053(.A(G107), .B(G116), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n252), .B(new_n255), .ZN(G351));
  OAI21_X1  g0056(.A(G20), .B1(new_n237), .B2(G50), .ZN(new_n257));
  INV_X1    g0057(.A(G150), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n204), .A2(G33), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT8), .B(G58), .ZN(new_n262));
  OAI221_X1 g0062(.A(new_n257), .B1(new_n258), .B2(new_n260), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n233), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n209), .ZN(new_n269));
  AND3_X1   g0069(.A1(new_n267), .A2(new_n233), .A3(new_n264), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT70), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n271), .B1(new_n204), .B2(G1), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n203), .A2(KEYINPUT70), .A3(G20), .ZN(new_n273));
  AND3_X1   g0073(.A1(new_n270), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G50), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n266), .A2(new_n269), .A3(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT3), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G222), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G223), .A2(G1698), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n281), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n233), .B1(G33), .B2(G41), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n285), .B(new_n286), .C1(G77), .C2(new_n281), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n203), .B(G274), .C1(G41), .C2(G45), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT69), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n288), .B(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G41), .ZN(new_n291));
  OAI211_X1 g0091(.A(G1), .B(G13), .C1(new_n278), .C2(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n287), .B(new_n290), .C1(new_n210), .C2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n295), .A2(G179), .ZN(new_n296));
  OR2_X1    g0096(.A1(new_n296), .A2(KEYINPUT71), .ZN(new_n297));
  INV_X1    g0097(.A(G169), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(KEYINPUT71), .ZN(new_n300));
  AND4_X1   g0100(.A1(new_n276), .A2(new_n297), .A3(new_n299), .A4(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n274), .A2(G77), .ZN(new_n302));
  XOR2_X1   g0102(.A(KEYINPUT15), .B(G87), .Z(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n304), .A2(new_n261), .ZN(new_n305));
  INV_X1    g0105(.A(G77), .ZN(new_n306));
  OAI22_X1  g0106(.A1(new_n262), .A2(new_n260), .B1(new_n204), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n265), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n302), .B(new_n308), .C1(G77), .C2(new_n267), .ZN(new_n309));
  NAND2_X1  g0109(.A1(G238), .A2(G1698), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n281), .B(new_n310), .C1(new_n219), .C2(G1698), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n311), .B(new_n286), .C1(G107), .C2(new_n281), .ZN(new_n312));
  INV_X1    g0112(.A(new_n294), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(new_n207), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n312), .A2(new_n290), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G190), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI211_X1 g0117(.A(new_n309), .B(new_n317), .C1(G200), .C2(new_n315), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n295), .A2(new_n316), .ZN(new_n319));
  XNOR2_X1  g0119(.A(new_n319), .B(KEYINPUT74), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT73), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n321), .B1(new_n295), .B2(G200), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT72), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n276), .A2(new_n323), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n266), .A2(new_n275), .A3(KEYINPUT72), .A4(new_n269), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n324), .A2(KEYINPUT9), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(KEYINPUT9), .B1(new_n324), .B2(new_n325), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n320), .B(new_n322), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT10), .ZN(new_n330));
  INV_X1    g0130(.A(new_n328), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n326), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT10), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n332), .A2(new_n333), .A3(new_n320), .A4(new_n322), .ZN(new_n334));
  AOI211_X1 g0134(.A(new_n301), .B(new_n318), .C1(new_n330), .C2(new_n334), .ZN(new_n335));
  XNOR2_X1  g0135(.A(new_n288), .B(KEYINPUT69), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n336), .B1(G238), .B2(new_n313), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT13), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n210), .A2(new_n282), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n281), .B(new_n339), .C1(G232), .C2(new_n282), .ZN(new_n340));
  NAND2_X1  g0140(.A1(G33), .A2(G97), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n286), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n337), .A2(new_n338), .A3(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n290), .B1(new_n212), .B2(new_n294), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n292), .B1(new_n340), .B2(new_n341), .ZN(new_n346));
  OAI21_X1  g0146(.A(KEYINPUT13), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(G190), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT75), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n344), .A2(new_n347), .A3(new_n350), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n337), .A2(new_n343), .A3(KEYINPUT75), .A4(new_n338), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(G200), .A3(new_n352), .ZN(new_n353));
  OAI22_X1  g0153(.A1(new_n260), .A2(new_n209), .B1(new_n204), .B2(G68), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n261), .A2(new_n306), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n265), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  XOR2_X1   g0156(.A(KEYINPUT76), .B(KEYINPUT11), .Z(new_n357));
  XNOR2_X1  g0157(.A(new_n356), .B(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n274), .A2(G68), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n268), .A2(new_n211), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n360), .B(KEYINPUT12), .ZN(new_n361));
  AND3_X1   g0161(.A1(new_n358), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n349), .A2(new_n353), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n351), .A2(G169), .A3(new_n352), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT77), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n366), .A2(KEYINPUT14), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n348), .A2(G179), .B1(new_n366), .B2(KEYINPUT14), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n351), .A2(G169), .A3(new_n367), .A4(new_n352), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n362), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n364), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OR2_X1    g0174(.A1(new_n315), .A2(G179), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n315), .A2(new_n298), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n375), .A2(new_n309), .A3(new_n376), .ZN(new_n377));
  AND2_X1   g0177(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT16), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n279), .A2(new_n204), .A3(new_n280), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT7), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n279), .A2(KEYINPUT7), .A3(new_n204), .A4(new_n280), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n211), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n218), .A2(new_n211), .ZN(new_n385));
  OAI21_X1  g0185(.A(G20), .B1(new_n385), .B2(new_n236), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n259), .A2(G159), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n379), .B1(new_n384), .B2(new_n388), .ZN(new_n389));
  AND2_X1   g0189(.A1(KEYINPUT3), .A2(G33), .ZN(new_n390));
  NOR2_X1   g0190(.A1(KEYINPUT3), .A2(G33), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(KEYINPUT7), .B1(new_n392), .B2(new_n204), .ZN(new_n393));
  INV_X1    g0193(.A(new_n383), .ZN(new_n394));
  OAI21_X1  g0194(.A(G68), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n388), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n395), .A2(KEYINPUT16), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n389), .A2(new_n397), .A3(new_n265), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n262), .A2(new_n268), .ZN(new_n399));
  INV_X1    g0199(.A(new_n262), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n274), .A2(new_n400), .ZN(new_n401));
  AND3_X1   g0201(.A1(new_n398), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n210), .A2(G1698), .ZN(new_n403));
  OAI221_X1 g0203(.A(new_n403), .B1(G223), .B2(G1698), .C1(new_n390), .C2(new_n391), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G87), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n292), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n294), .A2(new_n219), .ZN(new_n407));
  NOR3_X1   g0207(.A1(new_n406), .A2(new_n336), .A3(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(G200), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  XNOR2_X1  g0211(.A(KEYINPUT79), .B(G190), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n408), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n402), .A2(KEYINPUT17), .A3(new_n411), .A4(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n398), .A2(new_n399), .A3(new_n401), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n408), .A2(G169), .ZN(new_n416));
  NOR4_X1   g0216(.A1(new_n406), .A2(new_n336), .A3(new_n407), .A4(G179), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  XOR2_X1   g0219(.A(KEYINPUT78), .B(KEYINPUT18), .Z(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT17), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n398), .A2(new_n413), .A3(new_n399), .A4(new_n401), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n422), .B1(new_n423), .B2(new_n410), .ZN(new_n424));
  NOR2_X1   g0224(.A1(KEYINPUT78), .A2(KEYINPUT18), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n415), .A2(new_n418), .A3(new_n425), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n414), .A2(new_n421), .A3(new_n424), .A4(new_n426), .ZN(new_n427));
  XNOR2_X1  g0227(.A(new_n427), .B(KEYINPUT80), .ZN(new_n428));
  AND3_X1   g0228(.A1(new_n335), .A2(new_n378), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT87), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n212), .A2(new_n282), .ZN(new_n431));
  INV_X1    g0231(.A(G244), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(G1698), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n431), .B(new_n433), .C1(new_n390), .C2(new_n391), .ZN(new_n434));
  AND2_X1   g0234(.A1(G33), .A2(G116), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n286), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT85), .ZN(new_n439));
  INV_X1    g0239(.A(G250), .ZN(new_n440));
  INV_X1    g0240(.A(G45), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n440), .B1(new_n441), .B2(G1), .ZN(new_n442));
  INV_X1    g0242(.A(G274), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n203), .A2(new_n443), .A3(G45), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n292), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n438), .A2(new_n439), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n292), .B1(new_n434), .B2(new_n436), .ZN(new_n447));
  INV_X1    g0247(.A(new_n445), .ZN(new_n448));
  OAI21_X1  g0248(.A(KEYINPUT85), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n446), .A2(new_n449), .A3(G200), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT82), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT81), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n452), .B1(new_n203), .B2(G33), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n452), .A2(new_n203), .A3(G33), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n270), .A2(new_n451), .A3(new_n454), .A4(new_n455), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n455), .A2(new_n267), .A3(new_n233), .A4(new_n264), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT82), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n456), .A2(new_n458), .A3(G87), .ZN(new_n459));
  NOR2_X1   g0259(.A1(G97), .A2(G107), .ZN(new_n460));
  INV_X1    g0260(.A(G87), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n341), .A2(new_n204), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n462), .A2(new_n463), .A3(KEYINPUT19), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n204), .B(G68), .C1(new_n390), .C2(new_n391), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT19), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n466), .B1(new_n341), .B2(G20), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n464), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n468), .A2(new_n265), .B1(new_n268), .B2(new_n304), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n450), .A2(new_n459), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n439), .B1(new_n438), .B2(new_n445), .ZN(new_n471));
  NOR3_X1   g0271(.A1(new_n447), .A2(new_n448), .A3(KEYINPUT85), .ZN(new_n472));
  OAI21_X1  g0272(.A(G190), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(KEYINPUT86), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n446), .A2(new_n449), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT86), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n475), .A2(new_n476), .A3(G190), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n470), .B1(new_n474), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n475), .A2(G169), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n456), .A2(new_n458), .A3(new_n303), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n480), .A2(new_n469), .ZN(new_n481));
  AOI21_X1  g0281(.A(G179), .B1(new_n446), .B2(new_n449), .ZN(new_n482));
  NOR3_X1   g0282(.A1(new_n479), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n430), .B1(new_n478), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n482), .A2(new_n481), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n471), .A2(new_n472), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n298), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n476), .B1(new_n475), .B2(G190), .ZN(new_n489));
  AOI211_X1 g0289(.A(KEYINPUT86), .B(new_n316), .C1(new_n446), .C2(new_n449), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n488), .B(KEYINPUT87), .C1(new_n491), .C2(new_n470), .ZN(new_n492));
  NAND2_X1  g0292(.A1(G264), .A2(G1698), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n281), .B(new_n493), .C1(new_n221), .C2(G1698), .ZN(new_n494));
  XOR2_X1   g0294(.A(KEYINPUT88), .B(G303), .Z(new_n495));
  OAI211_X1 g0295(.A(new_n494), .B(new_n286), .C1(new_n281), .C2(new_n495), .ZN(new_n496));
  XNOR2_X1  g0296(.A(KEYINPUT5), .B(G41), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n441), .A2(G1), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n497), .A2(G274), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n286), .B1(new_n497), .B2(new_n498), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G270), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n496), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(G179), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(G116), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n268), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n270), .A2(G116), .A3(new_n454), .A4(new_n455), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G283), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT83), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT83), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n510), .A2(G33), .A3(G283), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n204), .B1(new_n220), .B2(G33), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n264), .A2(new_n233), .B1(G20), .B2(new_n505), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n515), .A2(KEYINPUT20), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT20), .B1(new_n515), .B2(new_n516), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n506), .B(new_n507), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n504), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n519), .A2(new_n502), .A3(G169), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT21), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n502), .A2(G200), .ZN(new_n524));
  INV_X1    g0324(.A(new_n519), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n496), .A2(new_n412), .A3(new_n501), .A4(new_n499), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n519), .A2(new_n502), .A3(KEYINPUT21), .A4(G169), .ZN(new_n528));
  AND4_X1   g0328(.A1(new_n520), .A2(new_n523), .A3(new_n527), .A4(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n484), .A2(new_n492), .A3(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT84), .ZN(new_n531));
  OAI211_X1 g0331(.A(G244), .B(new_n282), .C1(new_n390), .C2(new_n391), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT4), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n281), .A2(KEYINPUT4), .A3(G244), .A4(new_n282), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n281), .A2(G250), .A3(G1698), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n512), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n286), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n500), .A2(G257), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n539), .A2(G190), .A3(new_n499), .A4(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n267), .A2(G97), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(G107), .B1(new_n393), .B2(new_n394), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n260), .A2(new_n306), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT6), .ZN(new_n547));
  AND2_X1   g0347(.A1(G97), .A2(G107), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n547), .B1(new_n548), .B2(new_n460), .ZN(new_n549));
  INV_X1    g0349(.A(G107), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n550), .A2(KEYINPUT6), .A3(G97), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n204), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n544), .A2(new_n546), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n265), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n456), .A2(new_n458), .A3(G97), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n541), .A2(new_n543), .A3(new_n555), .A4(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n534), .A2(new_n535), .A3(new_n512), .A4(new_n537), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n558), .A2(new_n286), .B1(G257), .B2(new_n500), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n409), .B1(new_n559), .B2(new_n499), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n531), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n550), .B1(new_n382), .B2(new_n383), .ZN(new_n562));
  NOR3_X1   g0362(.A1(new_n562), .A2(new_n545), .A3(new_n552), .ZN(new_n563));
  INV_X1    g0363(.A(new_n265), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n543), .B(new_n556), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n539), .A2(new_n499), .A3(new_n540), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(G200), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n566), .A2(KEYINPUT84), .A3(new_n568), .A4(new_n541), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n561), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n567), .A2(new_n298), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n559), .A2(new_n503), .A3(new_n499), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n571), .A2(new_n565), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(KEYINPUT90), .B1(new_n204), .B2(G107), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT23), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n576), .A2(new_n577), .B1(new_n204), .B2(new_n435), .ZN(new_n578));
  OAI211_X1 g0378(.A(KEYINPUT90), .B(KEYINPUT23), .C1(new_n204), .C2(G107), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n204), .B(G87), .C1(new_n390), .C2(new_n391), .ZN(new_n580));
  XNOR2_X1  g0380(.A(KEYINPUT89), .B(KEYINPUT22), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n578), .B(new_n579), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT89), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT22), .ZN(new_n584));
  AND3_X1   g0384(.A1(new_n580), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(KEYINPUT24), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  OR2_X1    g0386(.A1(new_n580), .A2(new_n581), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n576), .A2(new_n577), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n435), .A2(new_n204), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n588), .A2(new_n579), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT24), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n580), .A2(new_n583), .A3(new_n584), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n587), .A2(new_n590), .A3(new_n591), .A4(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n586), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n265), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n456), .A2(new_n458), .A3(G107), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n267), .A2(G107), .ZN(new_n597));
  XNOR2_X1  g0397(.A(new_n597), .B(KEYINPUT25), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n595), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n499), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n221), .A2(G1698), .ZN(new_n601));
  OAI221_X1 g0401(.A(new_n601), .B1(G250), .B2(G1698), .C1(new_n390), .C2(new_n391), .ZN(new_n602));
  NAND2_X1  g0402(.A1(G33), .A2(G294), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n600), .B1(new_n604), .B2(new_n286), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n500), .A2(G264), .ZN(new_n606));
  AOI21_X1  g0406(.A(G169), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n606), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n607), .B1(new_n609), .B2(new_n503), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n599), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n596), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n612), .B1(new_n594), .B2(new_n265), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n608), .A2(G200), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n605), .A2(G190), .A3(new_n606), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n613), .A2(new_n598), .A3(new_n614), .A4(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n530), .A2(new_n575), .A3(new_n617), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n429), .A2(new_n618), .ZN(G372));
  NAND2_X1  g0419(.A1(new_n459), .A2(new_n469), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n438), .A2(new_n445), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n620), .B1(G200), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n622), .B1(new_n489), .B2(new_n490), .ZN(new_n623));
  AOI21_X1  g0423(.A(G169), .B1(new_n438), .B2(new_n445), .ZN(new_n624));
  OR3_X1    g0424(.A1(new_n482), .A2(new_n481), .A3(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT26), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n573), .A2(new_n623), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n625), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n484), .A2(new_n492), .A3(new_n573), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n628), .B1(new_n629), .B2(KEYINPUT26), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT91), .ZN(new_n631));
  NOR3_X1   g0431(.A1(new_n482), .A2(new_n481), .A3(new_n624), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n474), .A2(new_n477), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n632), .B1(new_n633), .B2(new_n622), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n599), .A2(new_n610), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n523), .A2(new_n520), .A3(new_n528), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n634), .B(new_n616), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n631), .B1(new_n637), .B2(new_n575), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n573), .B1(new_n561), .B2(new_n569), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n616), .A2(new_n623), .A3(new_n625), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n611), .A2(new_n520), .A3(new_n528), .A4(new_n523), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n639), .A2(new_n640), .A3(new_n641), .A4(KEYINPUT91), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n630), .A2(new_n638), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n429), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n414), .A2(new_n424), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n372), .A2(new_n373), .ZN(new_n646));
  INV_X1    g0446(.A(new_n377), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n363), .B(new_n645), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  XNOR2_X1  g0448(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n415), .A2(new_n418), .A3(KEYINPUT92), .ZN(new_n651));
  AOI21_X1  g0451(.A(KEYINPUT92), .B1(new_n415), .B2(new_n418), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT92), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n419), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n415), .A2(new_n418), .A3(KEYINPUT92), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(new_n656), .A3(new_n649), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n648), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n330), .A2(new_n334), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n301), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n644), .A2(new_n661), .ZN(G369));
  NOR2_X1   g0462(.A1(new_n228), .A2(G20), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  OR3_X1    g0464(.A1(new_n664), .A2(KEYINPUT27), .A3(G1), .ZN(new_n665));
  OAI21_X1  g0465(.A(KEYINPUT27), .B1(new_n664), .B2(G1), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(G213), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(G343), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n519), .A2(new_n669), .ZN(new_n670));
  MUX2_X1   g0470(.A(new_n636), .B(new_n529), .S(new_n670), .Z(new_n671));
  OR2_X1    g0471(.A1(new_n671), .A2(KEYINPUT94), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(KEYINPUT94), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(G330), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n616), .ZN(new_n677));
  INV_X1    g0477(.A(new_n669), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n678), .B1(new_n613), .B2(new_n598), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n611), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n635), .A2(new_n678), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n676), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n636), .A2(new_n678), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n617), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n684), .A2(new_n681), .A3(new_n686), .ZN(G399));
  INV_X1    g0487(.A(new_n230), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(G41), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n462), .A2(G116), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT95), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n689), .A2(new_n691), .A3(new_n203), .ZN(new_n692));
  INV_X1    g0492(.A(new_n238), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n692), .B1(new_n693), .B2(new_n689), .ZN(new_n694));
  XOR2_X1   g0494(.A(new_n694), .B(KEYINPUT96), .Z(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT28), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n484), .A2(new_n492), .A3(new_n626), .A4(new_n573), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n573), .A2(new_n623), .A3(new_n625), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n632), .B1(new_n699), .B2(KEYINPUT26), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n697), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n701), .A2(KEYINPUT29), .A3(new_n678), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n643), .A2(new_n678), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n702), .B1(new_n703), .B2(KEYINPUT29), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n504), .A2(new_n609), .A3(new_n559), .A4(new_n475), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT30), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n609), .A2(G179), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n708), .A2(new_n567), .A3(new_n621), .A4(new_n502), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n486), .A2(new_n608), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n710), .A2(KEYINPUT30), .A3(new_n559), .A4(new_n504), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n707), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n669), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  AOI22_X1  g0514(.A1(new_n618), .A2(new_n678), .B1(KEYINPUT31), .B2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT31), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n675), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n704), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n696), .B1(new_n720), .B2(G1), .ZN(G364));
  AOI21_X1  g0521(.A(new_n203), .B1(new_n663), .B2(G45), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n689), .A2(new_n723), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n204), .A2(new_n503), .A3(new_n409), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n412), .ZN(new_n726));
  INV_X1    g0526(.A(G326), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n204), .A2(G190), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT99), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n730), .A2(G179), .A3(G200), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n412), .A2(G20), .A3(G179), .A4(new_n409), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  AOI22_X1  g0533(.A1(new_n731), .A2(G329), .B1(G322), .B2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(G294), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n316), .A2(G179), .A3(G200), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(new_n204), .ZN(new_n737));
  INV_X1    g0537(.A(G311), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n729), .A2(G179), .A3(new_n409), .ZN(new_n739));
  OAI221_X1 g0539(.A(new_n734), .B1(new_n735), .B2(new_n737), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n409), .A2(G179), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n730), .A2(new_n742), .ZN(new_n743));
  AOI211_X1 g0543(.A(new_n728), .B(new_n740), .C1(G283), .C2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n725), .A2(new_n316), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(G317), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(KEYINPUT33), .ZN(new_n748));
  OR2_X1    g0548(.A1(new_n747), .A2(KEYINPUT33), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n746), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n742), .A2(new_n204), .A3(new_n316), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G303), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n744), .A2(new_n392), .A3(new_n750), .A4(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n737), .A2(new_n220), .ZN(new_n754));
  INV_X1    g0554(.A(new_n751), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n461), .ZN(new_n756));
  INV_X1    g0556(.A(new_n726), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n756), .B1(G50), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n731), .A2(G159), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n758), .B1(KEYINPUT32), .B2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n739), .ZN(new_n761));
  AOI211_X1 g0561(.A(new_n754), .B(new_n760), .C1(G77), .C2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n733), .A2(G58), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n759), .A2(KEYINPUT32), .ZN(new_n764));
  INV_X1    g0564(.A(new_n743), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n550), .ZN(new_n766));
  AOI211_X1 g0566(.A(new_n392), .B(new_n766), .C1(G68), .C2(new_n746), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n762), .A2(new_n763), .A3(new_n764), .A4(new_n767), .ZN(new_n768));
  AND2_X1   g0568(.A1(new_n753), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n298), .A2(KEYINPUT98), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n204), .B1(KEYINPUT98), .B2(new_n298), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n233), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n724), .B1(new_n769), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G13), .A2(G33), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(G20), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n773), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n688), .A2(new_n392), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G355), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n230), .A2(new_n392), .ZN(new_n782));
  XOR2_X1   g0582(.A(new_n782), .B(KEYINPUT97), .Z(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(G45), .B2(new_n238), .ZN(new_n784));
  AND2_X1   g0584(.A1(new_n252), .A2(G45), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n781), .B1(G116), .B2(new_n230), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n775), .B1(new_n779), .B2(new_n786), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n787), .B(KEYINPUT100), .Z(new_n788));
  INV_X1    g0588(.A(new_n778), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n671), .A2(new_n789), .ZN(new_n790));
  AND2_X1   g0590(.A1(new_n672), .A2(new_n673), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(G330), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n676), .A2(new_n724), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n788), .A2(new_n790), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(G396));
  AND2_X1   g0596(.A1(new_n309), .A2(new_n669), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n377), .B1(new_n318), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n647), .A2(new_n678), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n703), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n643), .A2(new_n678), .A3(new_n801), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  OR3_X1    g0604(.A1(new_n802), .A2(new_n719), .A3(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n724), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n719), .B1(new_n802), .B2(new_n804), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n731), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n392), .B1(new_n809), .B2(new_n738), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n765), .A2(new_n461), .ZN(new_n811));
  INV_X1    g0611(.A(G303), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n755), .A2(new_n550), .B1(new_n726), .B2(new_n812), .ZN(new_n813));
  OR4_X1    g0613(.A1(new_n754), .A2(new_n810), .A3(new_n811), .A4(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(G294), .B2(new_n733), .ZN(new_n815));
  INV_X1    g0615(.A(G283), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n815), .B1(new_n505), .B2(new_n739), .C1(new_n816), .C2(new_n745), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n733), .A2(G143), .B1(G159), .B2(new_n761), .ZN(new_n818));
  INV_X1    g0618(.A(G137), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n818), .B1(new_n819), .B2(new_n726), .C1(new_n258), .C2(new_n745), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT101), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT34), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n281), .B1(new_n218), .B2(new_n737), .C1(new_n755), .C2(new_n209), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n765), .A2(new_n211), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n823), .B(new_n824), .C1(G132), .C2(new_n731), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n817), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n806), .B1(new_n827), .B2(new_n773), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n773), .A2(new_n776), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n828), .B1(G77), .B2(new_n830), .C1(new_n777), .C2(new_n801), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n808), .A2(KEYINPUT102), .A3(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(KEYINPUT102), .B1(new_n808), .B2(new_n831), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(G384));
  NAND2_X1  g0636(.A1(new_n549), .A2(new_n551), .ZN(new_n837));
  OAI211_X1 g0637(.A(G20), .B(new_n234), .C1(new_n837), .C2(KEYINPUT35), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n505), .B(new_n838), .C1(KEYINPUT35), .C2(new_n837), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n839), .B(KEYINPUT36), .Z(new_n840));
  OAI21_X1  g0640(.A(G77), .B1(new_n218), .B2(new_n211), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n238), .A2(new_n841), .B1(G50), .B2(new_n211), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n842), .A2(G1), .A3(new_n228), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT103), .Z(new_n845));
  INV_X1    g0645(.A(KEYINPUT39), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n416), .A2(new_n417), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n402), .A2(new_n847), .B1(new_n423), .B2(new_n410), .ZN(new_n848));
  INV_X1    g0648(.A(new_n667), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n415), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(KEYINPUT37), .B1(new_n848), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT104), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT37), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n415), .A2(KEYINPUT104), .A3(new_n849), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n852), .B1(new_n848), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n427), .A2(new_n851), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n858), .A2(KEYINPUT38), .A3(new_n859), .ZN(new_n860));
  NOR3_X1   g0660(.A1(new_n651), .A2(new_n652), .A3(new_n650), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n649), .B1(new_n655), .B2(new_n656), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n645), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n854), .A2(new_n856), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n402), .A2(new_n411), .A3(new_n413), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n655), .A2(new_n865), .A3(new_n656), .ZN(new_n866));
  OAI21_X1  g0666(.A(KEYINPUT37), .B1(new_n866), .B2(new_n864), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n415), .A2(KEYINPUT104), .A3(new_n849), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT104), .B1(new_n415), .B2(new_n849), .ZN(new_n869));
  NOR3_X1   g0669(.A1(new_n868), .A2(new_n869), .A3(KEYINPUT37), .ZN(new_n870));
  INV_X1    g0670(.A(new_n848), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n863), .A2(new_n864), .B1(new_n867), .B2(new_n872), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n846), .B(new_n860), .C1(new_n873), .C2(KEYINPUT38), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n858), .A2(KEYINPUT38), .A3(new_n859), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT38), .B1(new_n858), .B2(new_n859), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT39), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n874), .A2(KEYINPUT105), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n646), .A2(new_n678), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT38), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n868), .A2(new_n869), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n882), .A2(new_n865), .A3(new_n655), .A4(new_n656), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n883), .A2(KEYINPUT37), .B1(new_n871), .B2(new_n870), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n882), .B1(new_n658), .B2(new_n645), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n881), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT105), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n886), .A2(new_n887), .A3(new_n846), .A4(new_n860), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n878), .A2(new_n880), .A3(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n658), .A2(new_n849), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n373), .A2(new_n669), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n374), .A2(new_n891), .B1(new_n646), .B2(new_n669), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n892), .B1(new_n803), .B2(new_n799), .ZN(new_n893));
  OR2_X1    g0693(.A1(new_n875), .A2(new_n876), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n890), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n889), .A2(new_n895), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n429), .B(new_n702), .C1(new_n703), .C2(KEYINPUT29), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n661), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n896), .B(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n886), .A2(new_n860), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n374), .A2(new_n891), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n646), .A2(new_n669), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n800), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n575), .A2(new_n617), .ZN(new_n904));
  INV_X1    g0704(.A(new_n530), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n904), .A2(new_n905), .A3(new_n678), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT106), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n713), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n712), .A2(KEYINPUT106), .A3(new_n669), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n908), .A2(new_n716), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n714), .A2(KEYINPUT31), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n906), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n900), .A2(KEYINPUT40), .A3(new_n903), .A4(new_n912), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n912), .B(new_n903), .C1(new_n875), .C2(new_n876), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT40), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n913), .A2(new_n916), .A3(new_n912), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n913), .A2(new_n916), .A3(G330), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n675), .B1(new_n715), .B2(new_n910), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n429), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n917), .A2(new_n429), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n899), .B(new_n921), .Z(new_n922));
  NOR2_X1   g0722(.A1(new_n663), .A2(new_n203), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n845), .B1(new_n922), .B2(new_n923), .ZN(G367));
  NAND2_X1  g0724(.A1(new_n620), .A2(new_n669), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n634), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n625), .B2(new_n925), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(KEYINPUT43), .ZN(new_n928));
  INV_X1    g0728(.A(new_n685), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n904), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT42), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n639), .B1(new_n566), .B2(new_n678), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n932), .A2(new_n611), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n669), .B1(new_n933), .B2(new_n574), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n928), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n927), .A2(KEYINPUT43), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n935), .B(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n573), .A2(new_n669), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n932), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n684), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n937), .B(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n689), .B(KEYINPUT41), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n686), .B1(new_n683), .B2(new_n929), .C1(new_n674), .C2(new_n675), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n686), .B1(new_n683), .B2(new_n929), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n676), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n947), .A2(new_n719), .A3(new_n704), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT107), .Z(new_n949));
  NAND2_X1  g0749(.A1(new_n686), .A2(new_n681), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n939), .A2(new_n950), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n951), .B(KEYINPUT44), .Z(new_n952));
  NOR2_X1   g0752(.A1(new_n939), .A2(new_n950), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT45), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n952), .B(new_n954), .C1(KEYINPUT108), .C2(new_n684), .ZN(new_n955));
  AND3_X1   g0755(.A1(new_n955), .A2(KEYINPUT108), .A3(new_n684), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n955), .B1(KEYINPUT108), .B2(new_n684), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(KEYINPUT109), .B1(new_n949), .B2(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n948), .B(KEYINPUT107), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT109), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n960), .B(new_n961), .C1(new_n956), .C2(new_n957), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n943), .B1(new_n963), .B2(new_n720), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n941), .B1(new_n964), .B2(new_n723), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n731), .A2(G317), .B1(new_n495), .B2(new_n733), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n966), .B(new_n392), .C1(new_n738), .C2(new_n726), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT46), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n755), .B2(new_n505), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n751), .A2(KEYINPUT46), .A3(G116), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n969), .B(new_n970), .C1(new_n735), .C2(new_n745), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT110), .ZN(new_n972));
  INV_X1    g0772(.A(new_n737), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n967), .B(new_n972), .C1(G107), .C2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n743), .A2(G97), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n974), .B(new_n975), .C1(new_n816), .C2(new_n739), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT111), .Z(new_n977));
  NOR2_X1   g0777(.A1(new_n732), .A2(new_n258), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n765), .A2(new_n306), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n757), .A2(G143), .B1(new_n751), .B2(G58), .ZN(new_n980));
  INV_X1    g0780(.A(G159), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n980), .B1(new_n981), .B2(new_n745), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n979), .B(new_n982), .C1(G50), .C2(new_n761), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n973), .A2(G68), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n731), .A2(G137), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n983), .A2(new_n281), .A3(new_n984), .A4(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n977), .B1(new_n978), .B2(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT47), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n773), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n927), .A2(new_n789), .ZN(new_n990));
  INV_X1    g0790(.A(new_n783), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n779), .B1(new_n230), .B2(new_n304), .C1(new_n991), .C2(new_n243), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n989), .A2(new_n724), .A3(new_n990), .A4(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT112), .Z(new_n994));
  NAND2_X1  g0794(.A1(new_n965), .A2(new_n994), .ZN(G387));
  OAI211_X1 g0795(.A(new_n949), .B(new_n689), .C1(new_n720), .C2(new_n947), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n947), .A2(new_n723), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n683), .A2(new_n789), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n392), .B1(new_n809), .B2(new_n727), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n757), .A2(G322), .B1(new_n746), .B2(G311), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT114), .Z(new_n1001));
  AOI22_X1  g0801(.A1(new_n733), .A2(G317), .B1(new_n495), .B2(new_n761), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT48), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1004), .B1(new_n816), .B2(new_n737), .C1(new_n735), .C2(new_n755), .ZN(new_n1005));
  XOR2_X1   g0805(.A(KEYINPUT115), .B(KEYINPUT49), .Z(new_n1006));
  XNOR2_X1  g0806(.A(new_n1005), .B(new_n1006), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n999), .B(new_n1007), .C1(G116), .C2(new_n743), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n809), .A2(new_n258), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n975), .B1(new_n211), .B2(new_n739), .C1(new_n262), .C2(new_n745), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1009), .B(new_n1010), .C1(G50), .C2(new_n733), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(new_n306), .B2(new_n755), .C1(new_n981), .C2(new_n726), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n304), .A2(new_n737), .ZN(new_n1013));
  NOR3_X1   g0813(.A1(new_n1012), .A2(new_n392), .A3(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n773), .B1(new_n1008), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n247), .A2(G45), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n783), .A2(new_n1016), .B1(new_n691), .B2(new_n780), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n400), .A2(new_n209), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT50), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n211), .A2(new_n306), .ZN(new_n1020));
  NOR4_X1   g0820(.A1(new_n1019), .A2(G45), .A3(new_n691), .A4(new_n1020), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n1017), .A2(new_n1021), .B1(G107), .B2(new_n230), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n806), .B1(new_n1022), .B2(new_n779), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1023), .B(KEYINPUT113), .Z(new_n1024));
  NAND2_X1  g0824(.A1(new_n1015), .A2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT116), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n996), .B(new_n997), .C1(new_n998), .C2(new_n1026), .ZN(G393));
  NAND2_X1  g0827(.A1(new_n949), .A2(new_n958), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n963), .A2(new_n689), .A3(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n958), .A2(new_n722), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n783), .A2(new_n255), .B1(G97), .B2(new_n688), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n779), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n939), .A2(new_n778), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n737), .A2(new_n306), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n1034), .B(new_n811), .C1(G143), .C2(new_n731), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n732), .A2(new_n981), .B1(new_n726), .B2(new_n258), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT51), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n761), .A2(new_n400), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n755), .A2(new_n211), .B1(new_n209), .B2(new_n745), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1039), .A2(new_n392), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1035), .A2(new_n1037), .A3(new_n1038), .A4(new_n1040), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n281), .B(new_n766), .C1(G322), .C2(new_n731), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n732), .A2(new_n738), .B1(new_n726), .B2(new_n747), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT52), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n746), .A2(new_n495), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n751), .A2(G283), .B1(new_n761), .B2(G294), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1042), .A2(new_n1044), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n737), .A2(new_n505), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1041), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n806), .B1(new_n1049), .B2(new_n773), .ZN(new_n1050));
  AND2_X1   g0850(.A1(new_n1033), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1030), .B1(new_n1032), .B2(new_n1051), .ZN(new_n1052));
  AND2_X1   g0852(.A1(new_n1029), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(G390));
  NAND2_X1  g0854(.A1(new_n878), .A2(new_n888), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n880), .B2(new_n893), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT117), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n863), .A2(new_n864), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n867), .A2(new_n872), .ZN(new_n1059));
  AOI21_X1  g0859(.A(KEYINPUT38), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n879), .B1(new_n1060), .B2(new_n875), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n701), .A2(new_n678), .A3(new_n798), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n892), .B1(new_n1062), .B2(new_n799), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1057), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n880), .B1(new_n886), .B2(new_n860), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1062), .A2(new_n799), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n892), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1065), .A2(new_n1068), .A3(KEYINPUT117), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1064), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n718), .A2(new_n801), .A3(new_n1067), .ZN(new_n1071));
  AND3_X1   g0871(.A1(new_n1056), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  AND3_X1   g0872(.A1(new_n912), .A2(new_n903), .A3(G330), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n1056), .B2(new_n1070), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n897), .A2(new_n661), .A3(new_n920), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n803), .A2(new_n799), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1067), .B1(new_n718), .B2(new_n801), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1077), .B1(new_n1078), .B2(new_n1073), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n912), .A2(G330), .A3(new_n801), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n892), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1071), .A2(new_n799), .A3(new_n1062), .A4(new_n1081), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n1079), .A2(new_n1082), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n1072), .A2(new_n1075), .B1(new_n1076), .B2(new_n1083), .ZN(new_n1084));
  NOR3_X1   g0884(.A1(new_n1061), .A2(new_n1057), .A3(new_n1063), .ZN(new_n1085));
  AOI21_X1  g0885(.A(KEYINPUT117), .B1(new_n1065), .B2(new_n1068), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1077), .A2(new_n1067), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n879), .A2(new_n1088), .B1(new_n878), .B2(new_n888), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1073), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1056), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1076), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1084), .A2(new_n689), .A3(new_n1093), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1072), .A2(new_n1075), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1055), .A2(new_n776), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n824), .B1(G294), .B2(new_n731), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT118), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n757), .A2(G283), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1034), .B1(new_n733), .B2(G116), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n220), .B2(new_n739), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n756), .B(new_n1101), .C1(G107), .C2(new_n746), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1098), .A2(new_n392), .A3(new_n1099), .A4(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n743), .A2(G50), .B1(G137), .B2(new_n746), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n731), .A2(G125), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1104), .B(new_n1105), .C1(new_n981), .C2(new_n737), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(G128), .B2(new_n757), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n733), .A2(G132), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n751), .A2(G150), .ZN(new_n1109));
  XOR2_X1   g0909(.A(new_n1109), .B(KEYINPUT53), .Z(new_n1110));
  XOR2_X1   g0910(.A(KEYINPUT54), .B(G143), .Z(new_n1111));
  AOI21_X1  g0911(.A(new_n392), .B1(new_n761), .B2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1107), .A2(new_n1108), .A3(new_n1110), .A4(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n774), .B1(new_n1103), .B2(new_n1113), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n806), .B(new_n1114), .C1(new_n262), .C2(new_n829), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1095), .A2(new_n723), .B1(new_n1096), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1094), .A2(new_n1116), .ZN(G378));
  INV_X1    g0917(.A(new_n301), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n660), .A2(new_n1118), .ZN(new_n1119));
  XOR2_X1   g0919(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n324), .A2(new_n325), .A3(new_n849), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1124));
  OR3_X1    g0924(.A1(new_n1122), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1123), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n776), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n724), .B1(G50), .B2(new_n830), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n757), .A2(G116), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n281), .A2(G41), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n761), .A2(new_n303), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1130), .A2(new_n984), .A3(new_n1131), .A4(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n765), .A2(new_n218), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n1133), .B(new_n1134), .C1(G283), .C2(new_n731), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n746), .A2(G97), .B1(new_n751), .B2(G77), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1135), .B(new_n1136), .C1(new_n550), .C2(new_n732), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1137), .B(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n209), .B1(new_n390), .B2(G41), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n757), .A2(G125), .B1(new_n751), .B2(new_n1111), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n733), .A2(G128), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n746), .A2(G132), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n973), .A2(G150), .B1(new_n761), .B2(G137), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .A4(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n291), .B1(new_n1145), .B2(KEYINPUT59), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(KEYINPUT120), .B(G124), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1146), .B1(new_n731), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1145), .A2(KEYINPUT59), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n743), .A2(G159), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1148), .A2(new_n278), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1139), .A2(new_n1140), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1129), .B1(new_n1152), .B2(new_n773), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1128), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n918), .A2(new_n889), .A3(new_n895), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n918), .B1(new_n889), .B2(new_n895), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1127), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n896), .A2(G330), .A3(new_n916), .A4(new_n913), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1127), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1159), .A2(new_n1160), .A3(new_n1155), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1158), .A2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1154), .B1(new_n1162), .B2(new_n722), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1076), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1093), .A2(new_n1165), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1166), .A2(KEYINPUT57), .A3(new_n1161), .A4(new_n1158), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(new_n689), .ZN(new_n1168));
  AND2_X1   g0968(.A1(new_n1158), .A2(new_n1161), .ZN(new_n1169));
  AOI21_X1  g0969(.A(KEYINPUT57), .B1(new_n1169), .B2(new_n1166), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1164), .B1(new_n1168), .B2(new_n1170), .ZN(G375));
  OAI21_X1  g0971(.A(new_n724), .B1(G68), .B2(new_n830), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT121), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1067), .A2(new_n777), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n746), .A2(new_n1111), .B1(G150), .B2(new_n761), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1175), .B1(new_n819), .B2(new_n732), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(G128), .B2(new_n731), .ZN(new_n1177));
  OAI21_X1  g0977(.A(KEYINPUT122), .B1(new_n1134), .B2(new_n392), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n973), .A2(G50), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n757), .A2(G132), .B1(new_n751), .B2(G159), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  NOR3_X1   g0981(.A1(new_n1134), .A2(KEYINPUT122), .A3(new_n392), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n979), .A2(new_n1013), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n751), .A2(G97), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n281), .B1(new_n733), .B2(G283), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n726), .A2(new_n735), .B1(new_n745), .B2(new_n505), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(new_n731), .B2(G303), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .A4(new_n1187), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n739), .A2(new_n550), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n1181), .A2(new_n1182), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1173), .B(new_n1174), .C1(new_n773), .C2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1083), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1191), .B1(new_n1192), .B2(new_n723), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1079), .A2(new_n1076), .A3(new_n1082), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n942), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1193), .B1(new_n1195), .B2(new_n1092), .ZN(G381));
  NAND3_X1  g0996(.A1(new_n965), .A2(new_n1053), .A3(new_n994), .ZN(new_n1197));
  OR2_X1    g0997(.A1(G384), .A2(G381), .ZN(new_n1198));
  NOR4_X1   g0998(.A1(new_n1197), .A2(G396), .A3(G393), .A4(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT57), .ZN(new_n1200));
  AND2_X1   g1000(.A1(new_n1093), .A2(new_n1165), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1200), .B1(new_n1201), .B2(new_n1162), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1202), .A2(new_n689), .A3(new_n1167), .ZN(new_n1203));
  INV_X1    g1003(.A(G378), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1203), .A2(new_n1204), .A3(new_n1164), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1199), .A2(new_n1206), .ZN(G407));
  OAI21_X1  g1007(.A(new_n1206), .B1(new_n1199), .B2(new_n668), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(G213), .ZN(G409));
  XNOR2_X1  g1009(.A(G393), .B(new_n795), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n965), .A2(new_n1053), .A3(new_n994), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1053), .B1(new_n965), .B2(new_n994), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1210), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(G387), .A2(G390), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1210), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1214), .A2(new_n1197), .A3(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1213), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT123), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1204), .B1(new_n1203), .B2(new_n1164), .ZN(new_n1219));
  NOR3_X1   g1019(.A1(new_n1201), .A2(new_n1162), .A3(new_n943), .ZN(new_n1220));
  NOR3_X1   g1020(.A1(new_n1220), .A2(G378), .A3(new_n1163), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1218), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(G375), .A2(G378), .ZN(new_n1223));
  OR3_X1    g1023(.A1(new_n1220), .A2(G378), .A3(new_n1163), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1223), .A2(KEYINPUT123), .A3(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n668), .A2(G213), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT60), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1194), .B1(new_n1092), .B2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1083), .A2(KEYINPUT60), .A3(new_n1076), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1228), .A2(new_n1229), .A3(new_n689), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT124), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n1193), .ZN(new_n1232));
  OR2_X1    g1032(.A1(new_n835), .A2(KEYINPUT125), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n835), .A2(KEYINPUT125), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1232), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1231), .A2(KEYINPUT125), .A3(new_n835), .A4(new_n1193), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1222), .A2(new_n1225), .A3(new_n1226), .A4(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT127), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT62), .ZN(new_n1240));
  AND3_X1   g1040(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1239), .B1(new_n1238), .B2(new_n1240), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1237), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1223), .A2(new_n1226), .A3(new_n1224), .ZN(new_n1244));
  NOR3_X1   g1044(.A1(new_n1243), .A2(new_n1240), .A3(new_n1244), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(new_n1241), .A2(new_n1242), .A3(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n668), .A2(G213), .A3(G2897), .ZN(new_n1247));
  XOR2_X1   g1047(.A(new_n1237), .B(new_n1247), .Z(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1244), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1217), .B1(new_n1246), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT63), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(new_n1243), .A2(new_n1253), .A3(new_n1244), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1217), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT61), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1222), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1253), .B1(new_n1248), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1238), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1255), .B(new_n1256), .C1(new_n1258), .C2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1252), .A2(new_n1260), .ZN(G405));
  NAND2_X1  g1061(.A1(new_n1217), .A2(new_n1243), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1213), .A2(new_n1216), .A3(new_n1237), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1206), .A2(new_n1219), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1264), .B(new_n1266), .ZN(G402));
endmodule


