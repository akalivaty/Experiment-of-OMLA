//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 1 1 1 1 1 0 1 1 0 1 0 1 0 1 1 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n529, new_n530, new_n531, new_n532, new_n533, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n544, new_n545,
    new_n546, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n605, new_n607, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1140, new_n1141;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT65), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  XNOR2_X1  g029(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT69), .Z(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n461), .B1(G2106), .B2(new_n452), .ZN(G319));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  INV_X1    g041(.A(G113), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  OAI22_X1  g043(.A1(new_n465), .A2(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT70), .A2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g048(.A1(KEYINPUT70), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(G2105), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G137), .ZN(new_n476));
  INV_X1    g051(.A(G2105), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n477), .A2(G101), .A3(G2104), .ZN(new_n478));
  AND3_X1   g053(.A1(new_n470), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT71), .ZN(G160));
  NAND2_X1  g055(.A1(new_n475), .A2(G136), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n477), .B1(new_n473), .B2(new_n474), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n477), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n481), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  NOR2_X1   g062(.A1(new_n477), .A2(G114), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT72), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT72), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n491), .A2(new_n493), .A3(new_n494), .A4(G2104), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  OAI211_X1 g071(.A(G138), .B(new_n477), .C1(new_n463), .C2(new_n464), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n474), .ZN(new_n500));
  AOI21_X1  g075(.A(KEYINPUT3), .B1(KEYINPUT70), .B2(G2104), .ZN(new_n501));
  OAI211_X1 g076(.A(G126), .B(G2105), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  AND2_X1   g077(.A1(KEYINPUT4), .A2(G138), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n477), .B(new_n503), .C1(new_n500), .C2(new_n501), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n496), .A2(new_n499), .A3(new_n502), .A4(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  XNOR2_X1  g081(.A(KEYINPUT6), .B(G651), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT5), .B(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G88), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n507), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G50), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n509), .A2(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n513), .A2(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  NAND3_X1  g093(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT73), .ZN(new_n520));
  INV_X1    g095(.A(new_n509), .ZN(new_n521));
  INV_X1    g096(.A(new_n511), .ZN(new_n522));
  AOI22_X1  g097(.A1(G89), .A2(new_n521), .B1(new_n522), .B2(G51), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT74), .ZN(new_n526));
  XOR2_X1   g101(.A(new_n526), .B(KEYINPUT7), .Z(new_n527));
  NOR2_X1   g102(.A1(new_n524), .A2(new_n527), .ZN(G168));
  INV_X1    g103(.A(G90), .ZN(new_n529));
  INV_X1    g104(.A(G52), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n509), .A2(new_n529), .B1(new_n511), .B2(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n515), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n531), .A2(new_n533), .ZN(G301));
  INV_X1    g109(.A(G301), .ZN(G171));
  XOR2_X1   g110(.A(KEYINPUT75), .B(G81), .Z(new_n536));
  INV_X1    g111(.A(G43), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n509), .A2(new_n536), .B1(new_n511), .B2(new_n537), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n515), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  NAND4_X1  g117(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g118(.A(KEYINPUT76), .B(KEYINPUT8), .Z(new_n544));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n544), .B(new_n545), .ZN(new_n546));
  NAND4_X1  g121(.A1(G319), .A2(G483), .A3(G661), .A4(new_n546), .ZN(G188));
  INV_X1    g122(.A(G65), .ZN(new_n548));
  XOR2_X1   g123(.A(KEYINPUT5), .B(G543), .Z(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(KEYINPUT79), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT79), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n508), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n548), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT80), .ZN(new_n554));
  AND2_X1   g129(.A1(G78), .A2(G543), .ZN(new_n555));
  OR3_X1    g130(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n554), .B1(new_n553), .B2(new_n555), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n556), .A2(G651), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n507), .A2(G53), .A3(G543), .ZN(new_n559));
  OAI21_X1  g134(.A(KEYINPUT9), .B1(new_n559), .B2(KEYINPUT77), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(KEYINPUT77), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n559), .A2(KEYINPUT77), .A3(KEYINPUT9), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n509), .A2(KEYINPUT78), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT78), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n508), .A2(new_n507), .A3(new_n565), .ZN(new_n566));
  AND2_X1   g141(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n562), .A2(new_n563), .B1(new_n567), .B2(G91), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n558), .A2(new_n568), .ZN(G299));
  INV_X1    g144(.A(G168), .ZN(G286));
  NAND2_X1  g145(.A1(new_n567), .A2(G87), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n508), .A2(G74), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n522), .A2(G49), .B1(new_n572), .B2(G651), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n573), .ZN(G288));
  AOI22_X1  g149(.A1(new_n508), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n575), .A2(new_n515), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT81), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n576), .A2(new_n577), .B1(G48), .B2(new_n522), .ZN(new_n578));
  OAI21_X1  g153(.A(KEYINPUT81), .B1(new_n575), .B2(new_n515), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n564), .A2(G86), .A3(new_n566), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G305));
  INV_X1    g156(.A(G85), .ZN(new_n582));
  INV_X1    g157(.A(G47), .ZN(new_n583));
  OAI22_X1  g158(.A1(new_n509), .A2(new_n582), .B1(new_n511), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n515), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n567), .A2(G92), .ZN(new_n590));
  XOR2_X1   g165(.A(new_n590), .B(KEYINPUT10), .Z(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  AND2_X1   g167(.A1(new_n550), .A2(new_n552), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n595), .A2(G651), .B1(G54), .B2(new_n522), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n589), .B1(new_n598), .B2(G868), .ZN(G284));
  OAI21_X1  g174(.A(new_n589), .B1(new_n598), .B2(G868), .ZN(G321));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(G299), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(new_n601), .B2(G168), .ZN(G297));
  OAI21_X1  g178(.A(new_n602), .B1(new_n601), .B2(G168), .ZN(G280));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n598), .B1(new_n605), .B2(G860), .ZN(G148));
  OAI21_X1  g181(.A(KEYINPUT82), .B1(new_n541), .B2(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n598), .A2(new_n605), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  MUX2_X1   g184(.A(KEYINPUT82), .B(new_n607), .S(new_n609), .Z(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g186(.A1(new_n482), .A2(G123), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT83), .Z(new_n613));
  NAND2_X1  g188(.A1(new_n475), .A2(G135), .ZN(new_n614));
  OAI21_X1  g189(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n615), .A2(KEYINPUT84), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(KEYINPUT84), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G111), .B2(new_n477), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n613), .B(new_n614), .C1(new_n616), .C2(new_n618), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(G2096), .Z(new_n620));
  NAND3_X1  g195(.A1(new_n477), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT12), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT13), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2100), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n620), .A2(new_n624), .ZN(G156));
  XNOR2_X1  g200(.A(G2427), .B(G2438), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2430), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT15), .B(G2435), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n629), .A2(KEYINPUT14), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G1341), .B(G1348), .Z(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n631), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT86), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2443), .B(G2446), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT87), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n637), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n635), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(G14), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n635), .A2(new_n640), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n642), .A2(new_n643), .ZN(G401));
  XOR2_X1   g219(.A(G2072), .B(G2078), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT17), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2067), .B(G2678), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(new_n648), .B2(new_n645), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n649), .B1(KEYINPUT88), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n652), .B1(KEYINPUT88), .B2(new_n651), .ZN(new_n653));
  INV_X1    g228(.A(new_n645), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n654), .A2(new_n650), .A3(new_n647), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT18), .Z(new_n656));
  NAND3_X1  g231(.A1(new_n646), .A2(new_n650), .A3(new_n648), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n653), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2096), .B(G2100), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(G227));
  XOR2_X1   g236(.A(G1971), .B(G1976), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT19), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1956), .B(G2474), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1961), .B(G1966), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AND2_X1   g241(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  NOR3_X1   g242(.A1(new_n663), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n663), .A2(new_n666), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT20), .Z(new_n670));
  AOI211_X1 g245(.A(new_n668), .B(new_n670), .C1(new_n663), .C2(new_n667), .ZN(new_n671));
  XOR2_X1   g246(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1991), .B(G1996), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1981), .B(G1986), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(G229));
  INV_X1    g252(.A(G288), .ZN(new_n678));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(new_n679), .B2(G23), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT33), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT90), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n679), .A2(G22), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(G166), .B2(new_n679), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G1971), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n686), .A2(G1971), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n684), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  MUX2_X1   g264(.A(G6), .B(G305), .S(G16), .Z(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT32), .B(G1981), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n681), .A2(new_n683), .ZN(new_n693));
  NOR3_X1   g268(.A1(new_n689), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT34), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g271(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n697));
  INV_X1    g272(.A(G107), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n697), .B1(new_n698), .B2(G2105), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n475), .A2(G131), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT89), .ZN(new_n701));
  AOI211_X1 g276(.A(new_n699), .B(new_n701), .C1(G119), .C2(new_n482), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G29), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G25), .B2(G29), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT35), .B(G1991), .Z(new_n705));
  AND2_X1   g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n704), .A2(new_n705), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n679), .A2(G24), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(new_n587), .B2(new_n679), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G1986), .ZN(new_n710));
  NOR3_X1   g285(.A1(new_n706), .A2(new_n707), .A3(new_n710), .ZN(new_n711));
  AND3_X1   g286(.A1(new_n696), .A2(KEYINPUT91), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(KEYINPUT91), .B1(new_n696), .B2(new_n711), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n694), .A2(new_n695), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT92), .B(KEYINPUT36), .Z(new_n716));
  OR3_X1    g291(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT36), .ZN(new_n718));
  OAI211_X1 g293(.A(KEYINPUT92), .B(new_n718), .C1(new_n714), .C2(new_n715), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n598), .A2(G16), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G4), .B2(G16), .ZN(new_n721));
  INV_X1    g296(.A(G1348), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT94), .B(KEYINPUT25), .Z(new_n724));
  NAND3_X1  g299(.A1(new_n477), .A2(G103), .A3(G2104), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G127), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n465), .A2(new_n727), .ZN(new_n728));
  AND2_X1   g303(.A1(G115), .A2(G2104), .ZN(new_n729));
  OAI21_X1  g304(.A(G2105), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n475), .A2(G139), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n726), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT95), .Z(new_n733));
  MUX2_X1   g308(.A(G33), .B(new_n733), .S(G29), .Z(new_n734));
  AOI21_X1  g309(.A(new_n723), .B1(G2072), .B2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(G29), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G32), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n482), .A2(G129), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT98), .ZN(new_n739));
  AND3_X1   g314(.A1(new_n477), .A2(G105), .A3(G2104), .ZN(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT26), .ZN(new_n742));
  AOI211_X1 g317(.A(new_n740), .B(new_n742), .C1(G141), .C2(new_n475), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n737), .B1(new_n744), .B2(new_n736), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT27), .B(G1996), .Z(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n736), .A2(G26), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT28), .Z(new_n749));
  OR2_X1    g324(.A1(G104), .A2(G2105), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n750), .B(G2104), .C1(G116), .C2(new_n477), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT93), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n475), .A2(G140), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n482), .A2(G128), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n749), .B1(new_n755), .B2(G29), .ZN(new_n756));
  INV_X1    g331(.A(G2067), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n747), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(G168), .A2(new_n679), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n679), .B2(G21), .ZN(new_n761));
  INV_X1    g336(.A(G1966), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(G2078), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n505), .A2(G29), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n736), .A2(G27), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n763), .B1(new_n764), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n764), .B2(new_n767), .ZN(new_n769));
  NOR2_X1   g344(.A1(G171), .A2(new_n679), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G5), .B2(new_n679), .ZN(new_n771));
  INV_X1    g346(.A(G1961), .ZN(new_n772));
  NOR2_X1   g347(.A1(G16), .A2(G19), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n541), .B2(G16), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n771), .A2(new_n772), .B1(G1341), .B2(new_n774), .ZN(new_n775));
  OAI221_X1 g350(.A(new_n775), .B1(new_n736), .B2(new_n619), .C1(G1341), .C2(new_n774), .ZN(new_n776));
  INV_X1    g351(.A(G28), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n777), .A2(KEYINPUT30), .ZN(new_n778));
  AOI21_X1  g353(.A(G29), .B1(new_n777), .B2(KEYINPUT30), .ZN(new_n779));
  OR2_X1    g354(.A1(KEYINPUT31), .A2(G11), .ZN(new_n780));
  NAND2_X1  g355(.A1(KEYINPUT31), .A2(G11), .ZN(new_n781));
  AOI22_X1  g356(.A1(new_n778), .A2(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI221_X1 g357(.A(new_n782), .B1(new_n771), .B2(new_n772), .C1(new_n761), .C2(new_n762), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n776), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n735), .A2(new_n759), .A3(new_n769), .A4(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(G34), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n786), .A2(KEYINPUT24), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n786), .A2(KEYINPUT24), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n736), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G160), .B2(new_n736), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT96), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(G2084), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT97), .Z(new_n793));
  INV_X1    g368(.A(G2090), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n736), .A2(G35), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT99), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n486), .B2(G29), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT100), .B(KEYINPUT29), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n797), .B(new_n798), .Z(new_n799));
  AOI22_X1  g374(.A1(new_n721), .A2(new_n722), .B1(new_n794), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n679), .A2(G20), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT23), .Z(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G299), .B2(G16), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G1956), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n791), .A2(G2084), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n734), .A2(G2072), .ZN(new_n806));
  INV_X1    g381(.A(new_n799), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n806), .B1(G2090), .B2(new_n807), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n800), .A2(new_n804), .A3(new_n805), .A4(new_n808), .ZN(new_n809));
  NOR3_X1   g384(.A1(new_n785), .A2(new_n793), .A3(new_n809), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n717), .A2(new_n719), .A3(new_n810), .ZN(G150));
  INV_X1    g386(.A(G150), .ZN(G311));
  INV_X1    g387(.A(G93), .ZN(new_n813));
  INV_X1    g388(.A(G55), .ZN(new_n814));
  OAI22_X1  g389(.A1(new_n509), .A2(new_n813), .B1(new_n511), .B2(new_n814), .ZN(new_n815));
  AOI22_X1  g390(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n816), .A2(new_n515), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(G860), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT37), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n598), .A2(G559), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT38), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n541), .B(new_n818), .Z(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n823), .B(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT39), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(new_n819), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n826), .A2(new_n827), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n821), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT101), .ZN(G145));
  XNOR2_X1  g407(.A(new_n733), .B(new_n744), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n702), .B(new_n622), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n489), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n494), .B1(new_n836), .B2(new_n493), .ZN(new_n837));
  NOR3_X1   g412(.A1(new_n488), .A2(new_n489), .A3(KEYINPUT72), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n502), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(KEYINPUT102), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n475), .A2(new_n503), .B1(new_n497), .B2(new_n498), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT102), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n496), .A2(new_n842), .A3(new_n502), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n840), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n755), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n475), .A2(G142), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT103), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n482), .A2(G130), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n477), .A2(G118), .ZN(new_n849));
  OAI21_X1  g424(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n847), .B(new_n848), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n845), .B(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n835), .B(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(G160), .B(new_n619), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(G162), .ZN(new_n855));
  AOI21_X1  g430(.A(G37), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n856), .B1(new_n855), .B2(new_n853), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g433(.A(new_n597), .B(G299), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT41), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n608), .B(new_n824), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n862), .B1(new_n861), .B2(new_n859), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n863), .A2(KEYINPUT105), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(KEYINPUT105), .ZN(new_n865));
  XNOR2_X1  g440(.A(G288), .B(G166), .ZN(new_n866));
  XNOR2_X1  g441(.A(G305), .B(new_n587), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT104), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n870), .A2(KEYINPUT42), .ZN(new_n871));
  INV_X1    g446(.A(new_n868), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n872), .A2(KEYINPUT42), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n864), .B1(new_n865), .B2(new_n874), .ZN(new_n875));
  NOR4_X1   g450(.A1(new_n863), .A2(new_n871), .A3(KEYINPUT105), .A4(new_n873), .ZN(new_n876));
  OAI21_X1  g451(.A(G868), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(G868), .B2(new_n818), .ZN(G295));
  OAI21_X1  g453(.A(new_n877), .B1(G868), .B2(new_n818), .ZN(G331));
  XNOR2_X1  g454(.A(new_n825), .B(G171), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(G286), .ZN(new_n881));
  INV_X1    g456(.A(new_n859), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT41), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n859), .B(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n883), .B1(new_n885), .B2(new_n881), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(new_n870), .ZN(new_n887));
  INV_X1    g462(.A(G37), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n883), .B(new_n869), .C1(new_n885), .C2(new_n881), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(KEYINPUT43), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n887), .A2(new_n889), .A3(new_n892), .A4(new_n888), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n891), .A2(KEYINPUT44), .A3(new_n893), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(G397));
  INV_X1    g473(.A(G1384), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT45), .B1(new_n844), .B2(new_n899), .ZN(new_n900));
  XOR2_X1   g475(.A(KEYINPUT106), .B(G40), .Z(new_n901));
  NAND4_X1  g476(.A1(new_n470), .A2(new_n476), .A3(new_n478), .A4(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(KEYINPUT107), .B1(new_n905), .B2(G1996), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT107), .ZN(new_n907));
  INV_X1    g482(.A(G1996), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n904), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(new_n744), .ZN(new_n911));
  OR2_X1    g486(.A1(new_n744), .A2(new_n908), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n755), .B(new_n757), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n911), .B1(new_n905), .B2(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n702), .B(new_n705), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n915), .B1(new_n904), .B2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  XOR2_X1   g493(.A(new_n587), .B(G1986), .Z(new_n919));
  AOI21_X1  g494(.A(new_n918), .B1(new_n904), .B2(new_n919), .ZN(new_n920));
  AOI22_X1  g495(.A1(G126), .A2(new_n482), .B1(new_n490), .B2(new_n495), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n841), .B1(new_n921), .B2(new_n842), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n496), .A2(new_n842), .A3(new_n502), .ZN(new_n923));
  OAI211_X1 g498(.A(KEYINPUT45), .B(new_n899), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n505), .A2(new_n899), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT45), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n902), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(G1971), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n842), .B1(new_n496), .B2(new_n502), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n499), .A2(new_n504), .ZN(new_n932));
  NOR3_X1   g507(.A1(new_n923), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT108), .B1(new_n933), .B2(G1384), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT50), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n844), .A2(new_n936), .A3(new_n899), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n934), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n925), .A2(KEYINPUT50), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(new_n903), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n930), .B1(new_n940), .B2(G2090), .ZN(new_n941));
  NAND2_X1  g516(.A1(G303), .A2(G8), .ZN(new_n942));
  XOR2_X1   g517(.A(new_n942), .B(KEYINPUT55), .Z(new_n943));
  NAND3_X1  g518(.A1(new_n941), .A2(G8), .A3(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n943), .B1(new_n941), .B2(G8), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT63), .ZN(new_n947));
  NOR3_X1   g522(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n678), .A2(G1976), .ZN(new_n949));
  INV_X1    g524(.A(G1976), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT52), .B1(G288), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n934), .A2(new_n903), .A3(new_n937), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n952), .A2(KEYINPUT109), .A3(G8), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT109), .B1(new_n952), .B2(G8), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n949), .B(new_n951), .C1(new_n953), .C2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(KEYINPUT110), .B(G1981), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n578), .A2(new_n579), .A3(new_n580), .A4(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(G86), .ZN(new_n958));
  INV_X1    g533(.A(G48), .ZN(new_n959));
  OAI22_X1  g534(.A1(new_n509), .A2(new_n958), .B1(new_n511), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(G1981), .B1(new_n960), .B2(new_n576), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT111), .B1(new_n957), .B2(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n962), .B(KEYINPUT49), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n963), .B1(new_n953), .B2(new_n954), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n955), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT52), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT109), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n932), .B1(KEYINPUT102), .B2(new_n839), .ZN(new_n968));
  AOI211_X1 g543(.A(KEYINPUT108), .B(G1384), .C1(new_n968), .C2(new_n843), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n936), .B1(new_n844), .B2(new_n899), .ZN(new_n970));
  NOR3_X1   g545(.A1(new_n969), .A2(new_n970), .A3(new_n902), .ZN(new_n971));
  INV_X1    g546(.A(G8), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n967), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n952), .A2(KEYINPUT109), .A3(G8), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n966), .B1(new_n975), .B2(new_n949), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n965), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n902), .A2(G2084), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n938), .A2(new_n939), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT114), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT45), .B1(new_n934), .B2(new_n937), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n903), .B1(new_n926), .B2(new_n925), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n762), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT114), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n938), .A2(new_n984), .A3(new_n939), .A4(new_n978), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n980), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n986), .A2(G8), .A3(G168), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n948), .A2(new_n977), .A3(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT50), .B1(new_n969), .B2(new_n970), .ZN(new_n990));
  INV_X1    g565(.A(new_n925), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n902), .B1(new_n991), .B2(new_n935), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n990), .A2(new_n794), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n972), .B1(new_n993), .B2(new_n930), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n944), .B1(new_n943), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n996), .B1(new_n965), .B2(new_n976), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n949), .B1(new_n953), .B2(new_n954), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT52), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n999), .A2(KEYINPUT113), .A3(new_n955), .A4(new_n964), .ZN(new_n1000));
  AOI211_X1 g575(.A(new_n995), .B(new_n987), .C1(new_n997), .C2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n989), .B1(new_n1001), .B2(KEYINPUT63), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n964), .A2(new_n950), .A3(new_n678), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n957), .ZN(new_n1004));
  XOR2_X1   g579(.A(new_n975), .B(KEYINPUT112), .Z(new_n1005));
  AOI22_X1  g580(.A1(new_n1004), .A2(new_n1005), .B1(new_n977), .B2(new_n945), .ZN(new_n1006));
  AOI21_X1  g581(.A(G1956), .B1(new_n990), .B2(new_n992), .ZN(new_n1007));
  XNOR2_X1  g582(.A(KEYINPUT56), .B(G2072), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n924), .A2(new_n927), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(KEYINPUT115), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT115), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n924), .A2(new_n927), .A3(new_n1011), .A4(new_n1008), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT57), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1014), .B1(new_n558), .B2(new_n568), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n558), .A2(new_n1014), .A3(new_n568), .ZN(new_n1016));
  OAI22_X1  g591(.A1(new_n1007), .A2(new_n1013), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n940), .A2(new_n722), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n971), .A2(new_n757), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT116), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1018), .A2(KEYINPUT116), .A3(new_n1019), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G1956), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n935), .B1(new_n934), .B2(new_n937), .ZN(new_n1026));
  INV_X1    g601(.A(new_n992), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1025), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1016), .A2(new_n1015), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1028), .A2(new_n1029), .A3(new_n1012), .A4(new_n1010), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(new_n598), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1017), .B1(new_n1024), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT118), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1017), .A2(new_n1030), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT61), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1033), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  AOI211_X1 g611(.A(KEYINPUT118), .B(KEYINPUT61), .C1(new_n1017), .C2(new_n1030), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1017), .A2(new_n1030), .A3(KEYINPUT61), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT59), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n1041));
  XOR2_X1   g616(.A(KEYINPUT58), .B(G1341), .Z(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n969), .A2(new_n970), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1043), .B1(new_n1044), .B2(new_n903), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n928), .A2(G1996), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1041), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n952), .A2(new_n1042), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1048), .B(KEYINPUT117), .C1(G1996), .C2(new_n928), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1040), .B1(new_n1050), .B2(new_n541), .ZN(new_n1051));
  INV_X1    g626(.A(new_n541), .ZN(new_n1052));
  AOI211_X1 g627(.A(KEYINPUT59), .B(new_n1052), .C1(new_n1047), .C2(new_n1049), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1039), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1038), .A2(new_n1054), .ZN(new_n1055));
  AOI221_X4 g630(.A(new_n1021), .B1(new_n971), .B2(new_n757), .C1(new_n940), .C2(new_n722), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT116), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1057));
  OR3_X1    g632(.A1(new_n1056), .A2(new_n1057), .A3(KEYINPUT60), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n597), .B1(new_n1024), .B2(KEYINPUT60), .ZN(new_n1059));
  OAI211_X1 g634(.A(KEYINPUT60), .B(new_n597), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1058), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1032), .B1(new_n1055), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT121), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n924), .A2(new_n927), .A3(new_n764), .ZN(new_n1065));
  XOR2_X1   g640(.A(KEYINPUT120), .B(KEYINPUT53), .Z(new_n1066));
  AOI22_X1  g641(.A1(new_n940), .A2(new_n772), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n764), .A2(KEYINPUT53), .ZN(new_n1068));
  OR3_X1    g643(.A1(new_n981), .A2(new_n982), .A3(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1067), .A2(G301), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT54), .ZN(new_n1071));
  INV_X1    g646(.A(G40), .ZN(new_n1072));
  INV_X1    g647(.A(new_n479), .ZN(new_n1073));
  NOR4_X1   g648(.A1(new_n900), .A2(new_n1072), .A3(new_n1073), .A4(new_n1068), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n924), .ZN(new_n1075));
  AOI21_X1  g650(.A(G301), .B1(new_n1067), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1064), .B1(new_n1071), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1076), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1078), .A2(KEYINPUT121), .A3(KEYINPUT54), .A4(new_n1070), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n995), .B1(new_n997), .B2(new_n1000), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1067), .A2(new_n1075), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1083), .A2(G171), .ZN(new_n1084));
  AOI21_X1  g659(.A(G301), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1082), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  AND2_X1   g661(.A1(new_n979), .A2(KEYINPUT114), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n983), .A2(new_n985), .ZN(new_n1088));
  OAI21_X1  g663(.A(G8), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(G168), .A2(new_n972), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT51), .B1(new_n1091), .B2(KEYINPUT119), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1089), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1094));
  OAI211_X1 g669(.A(G8), .B(new_n1092), .C1(new_n986), .C2(G286), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n986), .A2(new_n1090), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1080), .A2(new_n1081), .A3(new_n1086), .A4(new_n1097), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1002), .B(new_n1006), .C1(new_n1063), .C2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1097), .A2(KEYINPUT62), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT62), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1094), .A2(new_n1101), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1100), .A2(new_n1081), .A3(new_n1085), .A4(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT122), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1085), .ZN(new_n1106));
  AOI211_X1 g681(.A(new_n995), .B(new_n1106), .C1(new_n997), .C2(new_n1000), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1107), .A2(KEYINPUT122), .A3(new_n1102), .A4(new_n1100), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n920), .B1(new_n1099), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n702), .A2(new_n705), .ZN(new_n1111));
  XOR2_X1   g686(.A(new_n1111), .B(KEYINPUT123), .Z(new_n1112));
  NOR2_X1   g687(.A1(new_n915), .A2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n755), .A2(G2067), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT124), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT124), .ZN(new_n1116));
  OAI221_X1 g691(.A(new_n1116), .B1(G2067), .B2(new_n755), .C1(new_n915), .C2(new_n1112), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1115), .A2(new_n904), .A3(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n910), .A2(KEYINPUT46), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n913), .A2(new_n744), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1119), .B1(new_n904), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT125), .B1(new_n910), .B2(KEYINPUT46), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n910), .A2(KEYINPUT125), .A3(KEYINPUT46), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1121), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1121), .B(new_n1125), .C1(new_n1122), .C2(new_n1123), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n905), .A2(G1986), .A3(G290), .ZN(new_n1130));
  XOR2_X1   g705(.A(new_n1130), .B(KEYINPUT48), .Z(new_n1131));
  NAND2_X1  g706(.A1(new_n917), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1118), .A2(new_n1129), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT127), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1118), .A2(new_n1129), .A3(KEYINPUT127), .A4(new_n1132), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1110), .A2(new_n1137), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g713(.A1(new_n660), .A2(G319), .ZN(new_n1140));
  NOR3_X1   g714(.A1(G229), .A2(G401), .A3(new_n1140), .ZN(new_n1141));
  NAND3_X1  g715(.A1(new_n894), .A2(new_n857), .A3(new_n1141), .ZN(G225));
  INV_X1    g716(.A(G225), .ZN(G308));
endmodule


