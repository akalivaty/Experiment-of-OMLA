//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 0 0 0 1 1 1 0 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0 0 1 1 0 1 1 0 0 0 0 1 0 0 1 1 1 0 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n818, new_n820, new_n821,
    new_n822, new_n823, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT12), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G229gat), .A2(G233gat), .ZN(new_n208));
  XOR2_X1   g007(.A(G43gat), .B(G50gat), .Z(new_n209));
  INV_X1    g008(.A(KEYINPUT15), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XOR2_X1   g010(.A(new_n211), .B(KEYINPUT88), .Z(new_n212));
  INV_X1    g011(.A(G29gat), .ZN(new_n213));
  INV_X1    g012(.A(G36gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n215), .B(KEYINPUT14), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT89), .B1(new_n213), .B2(new_n214), .ZN(new_n217));
  OR3_X1    g016(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT89), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n209), .A2(new_n210), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n212), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n216), .B1(new_n213), .B2(new_n214), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(new_n220), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G15gat), .B(G22gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT16), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n226), .B1(new_n227), .B2(G1gat), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n228), .B1(G1gat), .B2(new_n226), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(G8gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n225), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT17), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n225), .B(new_n232), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n208), .B(new_n231), .C1(new_n233), .C2(new_n230), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT18), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n225), .B(new_n230), .ZN(new_n236));
  XOR2_X1   g035(.A(new_n208), .B(KEYINPUT13), .Z(new_n237));
  AOI22_X1  g036(.A1(new_n234), .A2(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n231), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n225), .B(KEYINPUT17), .ZN(new_n240));
  INV_X1    g039(.A(new_n230), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n242), .A2(KEYINPUT18), .A3(new_n208), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n207), .B1(new_n238), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n238), .A2(new_n207), .A3(new_n243), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G183gat), .ZN(new_n249));
  INV_X1    g048(.A(G190gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n253));
  OAI22_X1  g052(.A1(new_n249), .A2(new_n250), .B1(new_n253), .B2(KEYINPUT24), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n253), .A2(KEYINPUT24), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n251), .B(new_n252), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT25), .ZN(new_n257));
  INV_X1    g056(.A(G169gat), .ZN(new_n258));
  INV_X1    g057(.A(G176gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT23), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n257), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NOR3_X1   g061(.A1(new_n261), .A2(G169gat), .A3(G176gat), .ZN(new_n263));
  AND2_X1   g062(.A1(G169gat), .A2(G176gat), .ZN(new_n264));
  OAI21_X1  g063(.A(KEYINPUT66), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT66), .ZN(new_n266));
  NAND2_X1  g065(.A1(G169gat), .A2(G176gat), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n266), .B(new_n267), .C1(new_n260), .C2(new_n261), .ZN(new_n268));
  AND4_X1   g067(.A1(new_n256), .A2(new_n262), .A3(new_n265), .A4(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n259), .A2(KEYINPUT23), .ZN(new_n270));
  AND2_X1   g069(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n272));
  NOR3_X1   g071(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NOR2_X1   g072(.A1(G169gat), .A2(G176gat), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n267), .B1(new_n274), .B2(KEYINPUT23), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT65), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n264), .B1(new_n260), .B2(new_n261), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n261), .A2(G176gat), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT64), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(new_n258), .ZN(new_n280));
  NAND2_X1  g079(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n278), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT65), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n277), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n251), .A2(new_n252), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n276), .A2(new_n284), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n269), .B1(new_n289), .B2(new_n257), .ZN(new_n290));
  XNOR2_X1  g089(.A(KEYINPUT27), .B(G183gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n291), .A2(KEYINPUT28), .A3(new_n250), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT68), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(G183gat), .ZN(new_n294));
  AOI21_X1  g093(.A(G190gat), .B1(new_n294), .B2(KEYINPUT27), .ZN(new_n295));
  OR3_X1    g094(.A1(new_n249), .A2(KEYINPUT68), .A3(KEYINPUT27), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n292), .B1(new_n297), .B2(KEYINPUT28), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n264), .B1(new_n260), .B2(KEYINPUT26), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT26), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n274), .A2(new_n300), .ZN(new_n301));
  AOI22_X1  g100(.A1(new_n299), .A2(new_n301), .B1(G183gat), .B2(G190gat), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G226gat), .ZN(new_n304));
  INV_X1    g103(.A(G233gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI22_X1  g105(.A1(new_n290), .A2(new_n303), .B1(KEYINPUT29), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n289), .A2(new_n257), .ZN(new_n308));
  INV_X1    g107(.A(new_n269), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n298), .A2(new_n302), .ZN(new_n311));
  INV_X1    g110(.A(new_n306), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n307), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G211gat), .B(G218gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G211gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT73), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT73), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G211gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT22), .B1(new_n321), .B2(G218gat), .ZN(new_n322));
  XOR2_X1   g121(.A(G197gat), .B(G204gat), .Z(new_n323));
  OAI21_X1  g122(.A(new_n316), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n323), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT73), .B(G211gat), .ZN(new_n326));
  INV_X1    g125(.A(G218gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n315), .B(new_n325), .C1(new_n328), .C2(KEYINPUT22), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n324), .A2(new_n329), .A3(KEYINPUT74), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT74), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n331), .B(new_n316), .C1(new_n322), .C2(new_n323), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT75), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT75), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n330), .A2(new_n335), .A3(new_n332), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n314), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n307), .A2(new_n313), .A3(new_n333), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(KEYINPUT37), .A3(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G8gat), .B(G36gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(G64gat), .B(G92gat), .ZN(new_n341));
  XOR2_X1   g140(.A(new_n340), .B(new_n341), .Z(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n337), .A2(new_n338), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT85), .B(KEYINPUT37), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT86), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT86), .ZN(new_n348));
  AOI211_X1 g147(.A(new_n348), .B(new_n345), .C1(new_n337), .C2(new_n338), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n339), .B(new_n343), .C1(new_n347), .C2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT38), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT37), .ZN(new_n352));
  INV_X1    g151(.A(new_n333), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n352), .B1(new_n314), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n336), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n335), .B1(new_n330), .B2(new_n332), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n307), .B(new_n313), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT38), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n358), .B(new_n343), .C1(new_n347), .C2(new_n349), .ZN(new_n359));
  XNOR2_X1  g158(.A(G1gat), .B(G29gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(KEYINPUT0), .ZN(new_n361));
  XNOR2_X1  g160(.A(G57gat), .B(G85gat), .ZN(new_n362));
  XOR2_X1   g161(.A(new_n361), .B(new_n362), .Z(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(G225gat), .A2(G233gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n365), .B(KEYINPUT79), .ZN(new_n366));
  NAND2_X1  g165(.A1(G155gat), .A2(G162gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT2), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT76), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n367), .A2(KEYINPUT76), .A3(KEYINPUT2), .ZN(new_n371));
  INV_X1    g170(.A(G141gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(G148gat), .ZN(new_n373));
  INV_X1    g172(.A(G148gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(G141gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n370), .A2(new_n371), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(G155gat), .ZN(new_n378));
  INV_X1    g177(.A(G162gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n377), .A2(new_n367), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n367), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT78), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT77), .B1(new_n374), .B2(G141gat), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT77), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n386), .A2(new_n372), .A3(G148gat), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n385), .A2(new_n387), .A3(new_n375), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n380), .A2(KEYINPUT78), .A3(new_n367), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n384), .A2(new_n368), .A3(new_n388), .A4(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n381), .A2(new_n390), .ZN(new_n391));
  XOR2_X1   g190(.A(G127gat), .B(G134gat), .Z(new_n392));
  XNOR2_X1  g191(.A(G113gat), .B(G120gat), .ZN(new_n393));
  OR3_X1    g192(.A1(new_n392), .A2(KEYINPUT1), .A3(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n392), .B1(KEYINPUT1), .B2(new_n393), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n391), .A2(new_n396), .ZN(new_n397));
  AOI22_X1  g196(.A1(new_n381), .A2(new_n390), .B1(new_n394), .B2(new_n395), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n366), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT5), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n391), .A2(KEYINPUT3), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT3), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n381), .A2(new_n402), .A3(new_n390), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n401), .A2(new_n396), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n366), .ZN(new_n405));
  OAI211_X1 g204(.A(KEYINPUT80), .B(KEYINPUT4), .C1(new_n391), .C2(new_n396), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(KEYINPUT4), .B1(new_n391), .B2(new_n396), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n393), .A2(KEYINPUT1), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(new_n392), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT4), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n410), .A2(new_n411), .A3(new_n381), .A4(new_n390), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT80), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n408), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n400), .B1(new_n407), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n410), .B1(new_n391), .B2(KEYINPUT3), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n366), .B1(new_n416), .B2(new_n403), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n408), .A2(new_n412), .A3(KEYINPUT81), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT5), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT81), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n420), .B(KEYINPUT4), .C1(new_n391), .C2(new_n396), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n417), .A2(new_n418), .A3(new_n419), .A4(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n364), .B1(new_n415), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n417), .A2(new_n406), .ZN(new_n425));
  INV_X1    g224(.A(new_n414), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n363), .B(new_n422), .C1(new_n427), .C2(new_n400), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT6), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n424), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  OAI211_X1 g229(.A(KEYINPUT6), .B(new_n364), .C1(new_n415), .C2(new_n423), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n344), .A2(new_n342), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n351), .A2(new_n359), .A3(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT29), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n403), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n436), .B1(new_n355), .B2(new_n356), .ZN(new_n437));
  INV_X1    g236(.A(G228gat), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n438), .A2(new_n305), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n330), .A2(new_n435), .A3(new_n332), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n402), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n391), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n437), .A2(new_n439), .A3(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(G22gat), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n333), .A2(new_n436), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT29), .B1(new_n324), .B2(new_n329), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n391), .B1(new_n446), .B2(KEYINPUT3), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n439), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n443), .A2(new_n444), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n444), .B1(new_n443), .B2(new_n449), .ZN(new_n452));
  OAI21_X1  g251(.A(G78gat), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n443), .A2(new_n449), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(G22gat), .ZN(new_n455));
  INV_X1    g254(.A(G78gat), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n455), .A2(new_n456), .A3(new_n450), .ZN(new_n457));
  XNOR2_X1  g256(.A(KEYINPUT31), .B(G50gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n458), .B(KEYINPUT82), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n459), .B(G106gat), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n453), .A2(new_n457), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n460), .B1(new_n453), .B2(new_n457), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n434), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n418), .A2(new_n421), .ZN(new_n465));
  INV_X1    g264(.A(new_n404), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n366), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OR2_X1    g266(.A1(new_n397), .A2(new_n398), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n467), .B(KEYINPUT39), .C1(new_n366), .C2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT39), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n470), .B(new_n366), .C1(new_n465), .C2(new_n466), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT83), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n471), .A2(new_n472), .A3(new_n363), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n472), .B1(new_n471), .B2(new_n363), .ZN(new_n474));
  OAI211_X1 g273(.A(KEYINPUT40), .B(new_n469), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT30), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n344), .A2(new_n476), .A3(new_n342), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n337), .A2(new_n343), .A3(new_n338), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n432), .A2(KEYINPUT30), .A3(new_n478), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n475), .A2(new_n424), .A3(new_n477), .A4(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT84), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n469), .B1(new_n473), .B2(new_n474), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT40), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n482), .A2(new_n481), .A3(new_n483), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n480), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT87), .B1(new_n464), .B2(new_n487), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n479), .A2(new_n424), .A3(new_n477), .ZN(new_n489));
  INV_X1    g288(.A(new_n486), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n475), .B(new_n489), .C1(new_n490), .C2(new_n484), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT87), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n491), .A2(new_n492), .A3(new_n463), .A4(new_n434), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  XOR2_X1   g293(.A(G15gat), .B(G43gat), .Z(new_n495));
  XNOR2_X1  g294(.A(G71gat), .B(G99gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n495), .B(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n277), .A2(new_n282), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n287), .B1(new_n499), .B2(KEYINPUT65), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT25), .B1(new_n500), .B2(new_n284), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n410), .B(new_n311), .C1(new_n501), .C2(new_n269), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT69), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT69), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n310), .A2(new_n504), .A3(new_n410), .A4(new_n311), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n396), .B1(new_n290), .B2(new_n303), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n503), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(G227gat), .A2(G233gat), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT33), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n498), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT32), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n513), .B1(new_n507), .B2(new_n509), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n503), .A2(new_n505), .A3(new_n508), .A4(new_n506), .ZN(new_n517));
  XOR2_X1   g316(.A(new_n517), .B(KEYINPUT34), .Z(new_n518));
  AOI21_X1  g317(.A(KEYINPUT33), .B1(new_n507), .B2(new_n509), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n514), .B1(new_n519), .B2(new_n498), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n516), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT72), .ZN(new_n522));
  INV_X1    g321(.A(new_n518), .ZN(new_n523));
  NOR3_X1   g322(.A1(new_n514), .A2(new_n519), .A3(new_n498), .ZN(new_n524));
  AOI221_X4 g323(.A(new_n513), .B1(KEYINPUT33), .B2(new_n497), .C1(new_n507), .C2(new_n509), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT72), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n516), .A2(new_n518), .A3(new_n527), .A4(new_n520), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n522), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  OR2_X1    g329(.A1(new_n530), .A2(KEYINPUT36), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT70), .B1(new_n524), .B2(new_n525), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT70), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n516), .A2(new_n533), .A3(new_n520), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(KEYINPUT71), .B1(new_n535), .B2(new_n523), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT71), .ZN(new_n537));
  AOI211_X1 g336(.A(new_n537), .B(new_n518), .C1(new_n532), .C2(new_n534), .ZN(new_n538));
  OAI211_X1 g337(.A(KEYINPUT36), .B(new_n521), .C1(new_n536), .C2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n531), .A2(new_n539), .ZN(new_n540));
  AOI22_X1  g339(.A1(new_n477), .A2(new_n479), .B1(new_n430), .B2(new_n431), .ZN(new_n541));
  OR2_X1    g340(.A1(new_n463), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n494), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n460), .ZN(new_n544));
  NOR3_X1   g343(.A1(new_n451), .A2(new_n452), .A3(G78gat), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n456), .B1(new_n455), .B2(new_n450), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n453), .A2(new_n457), .A3(new_n460), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n547), .A2(new_n521), .A3(new_n548), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n541), .B(new_n549), .C1(new_n536), .C2(new_n538), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT35), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT35), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n541), .A2(new_n547), .A3(new_n552), .A4(new_n548), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n553), .A2(new_n529), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n248), .B1(new_n543), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(G57gat), .ZN(new_n559));
  INV_X1    g358(.A(G64gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G57gat), .A2(G64gat), .ZN(new_n562));
  INV_X1    g361(.A(G71gat), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n563), .A2(new_n456), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n561), .B(new_n562), .C1(new_n564), .C2(KEYINPUT9), .ZN(new_n565));
  NOR2_X1   g364(.A1(G71gat), .A2(G78gat), .ZN(new_n566));
  OR2_X1    g365(.A1(new_n566), .A2(KEYINPUT90), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n564), .A2(new_n566), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n565), .B(new_n567), .C1(new_n564), .C2(new_n566), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n572), .A2(KEYINPUT21), .ZN(new_n573));
  NAND2_X1  g372(.A1(G231gat), .A2(G233gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G127gat), .B(G155gat), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n576), .B(KEYINPUT91), .Z(new_n577));
  XNOR2_X1  g376(.A(new_n575), .B(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(G183gat), .B(G211gat), .Z(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n230), .B1(KEYINPUT21), .B2(new_n572), .ZN(new_n581));
  XNOR2_X1  g380(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n580), .B(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n586));
  INV_X1    g385(.A(new_n225), .ZN(new_n587));
  INV_X1    g386(.A(G85gat), .ZN(new_n588));
  INV_X1    g387(.A(G92gat), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT92), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT7), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n590), .B(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G99gat), .A2(G106gat), .ZN(new_n594));
  AOI22_X1  g393(.A1(KEYINPUT8), .A2(new_n594), .B1(new_n588), .B2(new_n589), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G99gat), .B(G106gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n586), .B1(new_n587), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n600), .B1(new_n240), .B2(new_n599), .ZN(new_n601));
  XOR2_X1   g400(.A(G190gat), .B(G218gat), .Z(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT93), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  OR2_X1    g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n601), .A2(new_n604), .ZN(new_n606));
  XNOR2_X1  g405(.A(G134gat), .B(G162gat), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  AND4_X1   g408(.A1(KEYINPUT94), .A2(new_n605), .A3(new_n606), .A4(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT94), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  AOI22_X1  g411(.A1(new_n612), .A2(new_n609), .B1(new_n605), .B2(new_n606), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G230gat), .A2(G233gat), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n598), .A2(new_n572), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT95), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT10), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n598), .A2(new_n572), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n617), .A2(KEYINPUT95), .A3(KEYINPUT10), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT96), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n616), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n625), .B1(new_n624), .B2(new_n623), .ZN(new_n626));
  XOR2_X1   g425(.A(G120gat), .B(G148gat), .Z(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT97), .ZN(new_n628));
  XOR2_X1   g427(.A(G176gat), .B(G204gat), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n621), .A2(new_n617), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n630), .B1(new_n631), .B2(new_n616), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n616), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n633), .B1(new_n623), .B2(new_n616), .ZN(new_n634));
  AOI22_X1  g433(.A1(new_n626), .A2(new_n632), .B1(new_n634), .B2(new_n630), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n585), .A2(new_n614), .A3(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n558), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n430), .A2(new_n431), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g440(.A1(new_n479), .A2(new_n477), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n558), .A2(new_n642), .A3(new_n636), .ZN(new_n643));
  XOR2_X1   g442(.A(KEYINPUT16), .B(G8gat), .Z(new_n644));
  AND2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(G8gat), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(KEYINPUT42), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n648), .B1(KEYINPUT42), .B2(new_n645), .ZN(G1325gat));
  AOI21_X1  g448(.A(G15gat), .B1(new_n637), .B2(new_n530), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT98), .ZN(new_n651));
  INV_X1    g450(.A(new_n540), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n652), .A2(G15gat), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n651), .B1(new_n637), .B2(new_n653), .ZN(G1326gat));
  INV_X1    g453(.A(new_n463), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n637), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(KEYINPUT43), .B(G22gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(G1327gat));
  AOI21_X1  g457(.A(KEYINPUT102), .B1(new_n551), .B2(new_n555), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT102), .ZN(new_n660));
  AOI211_X1 g459(.A(new_n660), .B(new_n554), .C1(new_n550), .C2(KEYINPUT35), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n543), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT103), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n543), .B(KEYINPUT103), .C1(new_n659), .C2(new_n661), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n614), .A2(KEYINPUT44), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n543), .A2(new_n556), .ZN(new_n668));
  OAI21_X1  g467(.A(KEYINPUT44), .B1(new_n668), .B2(new_n614), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n584), .B(KEYINPUT100), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n635), .B(KEYINPUT101), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n671), .A2(new_n248), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(G29gat), .B1(new_n674), .B2(new_n638), .ZN(new_n675));
  INV_X1    g474(.A(new_n614), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n676), .A2(new_n584), .A3(new_n635), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT99), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n557), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n679), .A2(new_n213), .A3(new_n639), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT45), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n675), .A2(new_n681), .ZN(G1328gat));
  INV_X1    g481(.A(new_n642), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n679), .A2(new_n214), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n684), .B(KEYINPUT46), .Z(new_n685));
  OAI21_X1  g484(.A(G36gat), .B1(new_n674), .B2(new_n642), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(G1329gat));
  INV_X1    g486(.A(G43gat), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n679), .A2(new_n688), .A3(new_n530), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n674), .A2(new_n540), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n689), .B1(new_n690), .B2(new_n688), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT47), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OAI211_X1 g492(.A(KEYINPUT47), .B(new_n689), .C1(new_n690), .C2(new_n688), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(G1330gat));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n696));
  INV_X1    g495(.A(G50gat), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n655), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT104), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n557), .A2(new_n696), .A3(new_n678), .A4(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(KEYINPUT48), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n679), .A2(new_n699), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n701), .B1(new_n702), .B2(KEYINPUT105), .ZN(new_n703));
  INV_X1    g502(.A(new_n673), .ZN(new_n704));
  AOI211_X1 g503(.A(new_n463), .B(new_n704), .C1(new_n667), .C2(new_n669), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n703), .B1(new_n705), .B2(new_n697), .ZN(new_n706));
  INV_X1    g505(.A(new_n702), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n670), .A2(new_n655), .A3(new_n673), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n707), .B1(new_n708), .B2(G50gat), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n706), .B1(new_n709), .B2(KEYINPUT48), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT106), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n706), .B(new_n712), .C1(new_n709), .C2(KEYINPUT48), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(new_n713), .ZN(G1331gat));
  AND2_X1   g513(.A1(new_n664), .A2(new_n665), .ZN(new_n715));
  INV_X1    g514(.A(new_n672), .ZN(new_n716));
  NOR4_X1   g515(.A1(new_n716), .A2(new_n247), .A3(new_n676), .A4(new_n584), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n718), .A2(new_n638), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(new_n559), .ZN(G1332gat));
  INV_X1    g519(.A(new_n718), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n642), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(KEYINPUT107), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT107), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n721), .A2(new_n725), .A3(new_n722), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n724), .A2(new_n728), .A3(new_n726), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(G1333gat));
  OAI21_X1  g531(.A(G71gat), .B1(new_n718), .B2(new_n540), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n530), .A2(new_n563), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n718), .B2(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n735), .B(new_n737), .ZN(G1334gat));
  NOR2_X1   g537(.A1(new_n718), .A2(new_n463), .ZN(new_n739));
  XNOR2_X1  g538(.A(KEYINPUT109), .B(G78gat), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1335gat));
  INV_X1    g540(.A(new_n635), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n248), .A2(new_n584), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT110), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n670), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(G85gat), .B1(new_n745), .B2(new_n638), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n676), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  AND3_X1   g547(.A1(new_n662), .A2(new_n748), .A3(KEYINPUT51), .ZN(new_n749));
  AOI21_X1  g548(.A(KEYINPUT51), .B1(new_n662), .B2(new_n748), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n742), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n639), .A2(new_n588), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n746), .B1(new_n751), .B2(new_n752), .ZN(G1336gat));
  NOR2_X1   g552(.A1(new_n642), .A2(G92gat), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n672), .B(new_n754), .C1(new_n749), .C2(new_n750), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n745), .A2(new_n642), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n755), .B1(new_n756), .B2(new_n589), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT52), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT52), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n759), .B(new_n755), .C1(new_n756), .C2(new_n589), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(G1337gat));
  OAI21_X1  g560(.A(G99gat), .B1(new_n745), .B2(new_n540), .ZN(new_n762));
  OR2_X1    g561(.A1(new_n529), .A2(G99gat), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n762), .B1(new_n751), .B2(new_n763), .ZN(G1338gat));
  OAI21_X1  g563(.A(G106gat), .B1(new_n745), .B2(new_n463), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n463), .A2(G106gat), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n672), .B(new_n766), .C1(new_n749), .C2(new_n750), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT111), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n769), .B1(new_n767), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n765), .B(new_n767), .C1(new_n770), .C2(new_n769), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(G1339gat));
  INV_X1    g573(.A(KEYINPUT113), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n242), .A2(new_n208), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n236), .A2(new_n237), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n205), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n246), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n775), .B1(new_n779), .B2(new_n635), .ZN(new_n780));
  INV_X1    g579(.A(new_n246), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n622), .A2(new_n621), .ZN(new_n782));
  XOR2_X1   g581(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n783));
  NAND4_X1  g582(.A1(new_n782), .A2(new_n615), .A3(new_n620), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n630), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT54), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n786), .B1(new_n623), .B2(new_n616), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n785), .B1(new_n626), .B2(new_n787), .ZN(new_n788));
  OAI22_X1  g587(.A1(new_n781), .A2(new_n244), .B1(new_n788), .B2(KEYINPUT55), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(KEYINPUT55), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n626), .A2(new_n632), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n780), .B1(new_n789), .B2(new_n792), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n779), .A2(new_n775), .A3(new_n635), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n614), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n788), .A2(KEYINPUT55), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n614), .A2(new_n779), .A3(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n792), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n671), .B1(new_n795), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n636), .A2(new_n247), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n802), .A2(new_n463), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n683), .A2(new_n638), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n803), .A2(new_n530), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(G113gat), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n805), .A2(new_n806), .A3(new_n248), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n536), .A2(new_n538), .ZN(new_n808));
  INV_X1    g607(.A(new_n549), .ZN(new_n809));
  INV_X1    g608(.A(new_n804), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n802), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(G113gat), .B1(new_n812), .B2(new_n247), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n807), .A2(new_n813), .ZN(G1340gat));
  OAI21_X1  g613(.A(G120gat), .B1(new_n805), .B2(new_n716), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n635), .A2(G120gat), .ZN(new_n816));
  XOR2_X1   g615(.A(new_n816), .B(KEYINPUT114), .Z(new_n817));
  NAND2_X1  g616(.A1(new_n812), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n815), .A2(new_n818), .ZN(G1341gat));
  INV_X1    g618(.A(new_n671), .ZN(new_n820));
  OAI21_X1  g619(.A(G127gat), .B1(new_n805), .B2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(G127gat), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n812), .A2(new_n822), .A3(new_n585), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(G1342gat));
  INV_X1    g623(.A(G134gat), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n812), .A2(new_n825), .A3(new_n676), .ZN(new_n826));
  OR2_X1    g625(.A1(new_n826), .A2(KEYINPUT56), .ZN(new_n827));
  OAI21_X1  g626(.A(G134gat), .B1(new_n805), .B2(new_n614), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(KEYINPUT56), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(G1343gat));
  NOR2_X1   g629(.A1(new_n652), .A2(new_n810), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n802), .A2(new_n655), .ZN(new_n833));
  XOR2_X1   g632(.A(KEYINPUT115), .B(KEYINPUT57), .Z(new_n834));
  OR2_X1    g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT116), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n742), .A2(new_n836), .A3(new_n246), .A4(new_n778), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT116), .B1(new_n779), .B2(new_n635), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n837), .B(new_n838), .C1(new_n789), .C2(new_n792), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n614), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n585), .B1(new_n840), .B2(new_n799), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n655), .B1(new_n841), .B2(new_n801), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT57), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n832), .B1(new_n835), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n372), .B1(new_n846), .B2(new_n247), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n833), .A2(new_n831), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n247), .A2(new_n372), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(KEYINPUT58), .B1(new_n847), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n833), .A2(new_n834), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n831), .B1(new_n852), .B2(new_n844), .ZN(new_n853));
  OAI21_X1  g652(.A(G141gat), .B1(new_n853), .B2(new_n248), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT58), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n854), .B(new_n855), .C1(new_n848), .C2(new_n849), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n851), .A2(new_n856), .ZN(G1344gat));
  NAND2_X1  g656(.A1(new_n842), .A2(new_n843), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT118), .ZN(new_n859));
  AOI22_X1  g658(.A1(new_n839), .A2(new_n614), .B1(new_n797), .B2(new_n798), .ZN(new_n860));
  OAI22_X1  g659(.A1(new_n860), .A2(new_n585), .B1(new_n247), .B2(new_n636), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT57), .B1(new_n861), .B2(new_n655), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT118), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n655), .B(new_n834), .C1(new_n800), .C2(new_n801), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n859), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n831), .A2(KEYINPUT117), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n831), .A2(KEYINPUT117), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n868), .A2(new_n742), .A3(new_n869), .ZN(new_n870));
  OAI211_X1 g669(.A(KEYINPUT59), .B(G148gat), .C1(new_n867), .C2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(new_n848), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n374), .A3(new_n742), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n374), .B1(new_n846), .B2(new_n742), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n871), .B(new_n873), .C1(new_n874), .C2(KEYINPUT59), .ZN(G1345gat));
  OAI21_X1  g674(.A(G155gat), .B1(new_n853), .B2(new_n820), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n872), .A2(new_n378), .A3(new_n585), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1346gat));
  AOI21_X1  g677(.A(G162gat), .B1(new_n872), .B2(new_n676), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n614), .A2(new_n379), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n879), .B1(new_n846), .B2(new_n880), .ZN(G1347gat));
  NAND2_X1  g680(.A1(new_n683), .A2(new_n638), .ZN(new_n882));
  XOR2_X1   g681(.A(new_n882), .B(KEYINPUT119), .Z(new_n883));
  AND2_X1   g682(.A1(new_n883), .A2(new_n530), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n803), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(G169gat), .B1(new_n885), .B2(new_n248), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n802), .A2(new_n638), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n808), .A2(new_n809), .A3(new_n642), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n247), .A2(new_n280), .A3(new_n281), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n886), .B1(new_n889), .B2(new_n890), .ZN(G1348gat));
  OAI21_X1  g690(.A(new_n259), .B1(new_n889), .B2(new_n635), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT120), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n885), .A2(new_n259), .A3(new_n716), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n893), .A2(new_n894), .ZN(G1349gat));
  NAND4_X1  g694(.A1(new_n802), .A2(new_n463), .A3(new_n671), .A4(new_n884), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n249), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n898), .B1(new_n897), .B2(new_n896), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n887), .A2(new_n291), .A3(new_n585), .A4(new_n888), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT60), .ZN(new_n901));
  AOI22_X1  g700(.A1(new_n899), .A2(new_n900), .B1(KEYINPUT122), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n901), .A2(KEYINPUT122), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n902), .B(new_n903), .ZN(G1350gat));
  OAI21_X1  g703(.A(G190gat), .B1(new_n885), .B2(new_n614), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT61), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n676), .A2(new_n250), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n906), .B1(new_n889), .B2(new_n907), .ZN(G1351gat));
  NOR3_X1   g707(.A1(new_n652), .A2(new_n642), .A3(new_n463), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT123), .ZN(new_n910));
  OR2_X1    g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n910), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n887), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(G197gat), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n913), .A2(new_n914), .A3(new_n247), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n540), .A2(new_n883), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT124), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n865), .B1(new_n862), .B2(new_n863), .ZN(new_n918));
  AOI211_X1 g717(.A(KEYINPUT118), .B(KEYINPUT57), .C1(new_n861), .C2(new_n655), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(KEYINPUT125), .B1(new_n920), .B2(new_n248), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(G197gat), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n920), .A2(KEYINPUT125), .A3(new_n248), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n915), .B1(new_n922), .B2(new_n923), .ZN(G1352gat));
  XNOR2_X1  g723(.A(KEYINPUT126), .B(G204gat), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n913), .A2(new_n742), .A3(new_n925), .ZN(new_n926));
  OR2_X1    g725(.A1(new_n926), .A2(KEYINPUT62), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(KEYINPUT62), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n920), .A2(new_n716), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n927), .B(new_n928), .C1(new_n929), .C2(new_n925), .ZN(G1353gat));
  NAND3_X1  g729(.A1(new_n913), .A2(new_n326), .A3(new_n585), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT127), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n866), .A2(new_n932), .A3(new_n585), .A4(new_n917), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n933), .A2(G211gat), .ZN(new_n934));
  OAI21_X1  g733(.A(KEYINPUT127), .B1(new_n920), .B2(new_n584), .ZN(new_n935));
  AOI21_X1  g734(.A(KEYINPUT63), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AND4_X1   g735(.A1(KEYINPUT63), .A2(new_n935), .A3(G211gat), .A4(new_n933), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n931), .B1(new_n936), .B2(new_n937), .ZN(G1354gat));
  OAI21_X1  g737(.A(G218gat), .B1(new_n920), .B2(new_n614), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n913), .A2(new_n327), .A3(new_n676), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(G1355gat));
endmodule


