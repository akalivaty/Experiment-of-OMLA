//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 0 1 0 1 0 0 1 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972;
  INV_X1    g000(.A(G119), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT23), .B1(new_n187), .B2(G128), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n187), .A2(G128), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  AOI21_X1  g008(.A(KEYINPUT74), .B1(new_n194), .B2(G110), .ZN(new_n195));
  AOI22_X1  g009(.A1(new_n188), .A2(new_n191), .B1(new_n187), .B2(G128), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT74), .ZN(new_n197));
  INV_X1    g011(.A(G110), .ZN(new_n198));
  NOR3_X1   g012(.A1(new_n196), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n195), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n190), .A2(G119), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n193), .A2(new_n201), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT24), .B(G110), .ZN(new_n203));
  OR2_X1    g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  AND2_X1   g018(.A1(G125), .A2(G140), .ZN(new_n205));
  NOR2_X1   g019(.A1(G125), .A2(G140), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT16), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT16), .ZN(new_n208));
  INV_X1    g022(.A(G140), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n209), .A3(G125), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  AOI21_X1  g026(.A(KEYINPUT76), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT76), .ZN(new_n214));
  AOI211_X1 g028(.A(new_n214), .B(G146), .C1(new_n207), .C2(new_n210), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G125), .ZN(new_n217));
  NOR3_X1   g031(.A1(new_n217), .A2(KEYINPUT16), .A3(G140), .ZN(new_n218));
  XNOR2_X1  g032(.A(G125), .B(G140), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n218), .B1(new_n219), .B2(KEYINPUT16), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT75), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n221), .A3(G146), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n207), .A2(G146), .A3(new_n210), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(KEYINPUT75), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n200), .B(new_n204), .C1(new_n216), .C2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT77), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n227), .B1(new_n219), .B2(new_n212), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n227), .B(new_n212), .C1(new_n205), .C2(new_n206), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  OR2_X1    g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n202), .A2(new_n203), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n232), .B1(new_n194), .B2(G110), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n231), .A2(KEYINPUT78), .A3(new_n233), .A4(new_n223), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT78), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n223), .B1(new_n228), .B2(new_n230), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n196), .A2(new_n198), .B1(new_n202), .B2(new_n203), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n226), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT22), .B(G137), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n241), .B(KEYINPUT79), .ZN(new_n242));
  INV_X1    g056(.A(G953), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n243), .A2(G221), .A3(G234), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n242), .B(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n240), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n226), .A2(new_n239), .A3(new_n245), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G902), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(KEYINPUT80), .A3(KEYINPUT25), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT25), .ZN(new_n253));
  AOI21_X1  g067(.A(G902), .B1(new_n247), .B2(new_n248), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT80), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G217), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n257), .B1(G234), .B2(new_n250), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n252), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n258), .A2(G902), .ZN(new_n260));
  XOR2_X1   g074(.A(new_n260), .B(KEYINPUT81), .Z(new_n261));
  NAND2_X1  g075(.A1(new_n249), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT65), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT11), .ZN(new_n265));
  INV_X1    g079(.A(G134), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n265), .B1(new_n266), .B2(G137), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(G137), .ZN(new_n268));
  INV_X1    g082(.A(G137), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(KEYINPUT11), .A3(G134), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n267), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G131), .ZN(new_n272));
  INV_X1    g086(.A(G131), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n267), .A2(new_n270), .A3(new_n273), .A4(new_n268), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT64), .ZN(new_n276));
  XNOR2_X1  g090(.A(G143), .B(G146), .ZN(new_n277));
  XNOR2_X1  g091(.A(KEYINPUT0), .B(G128), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n212), .A2(G143), .ZN(new_n280));
  INV_X1    g094(.A(G143), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G146), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(KEYINPUT0), .A2(G128), .ZN(new_n284));
  OR2_X1    g098(.A1(KEYINPUT0), .A2(G128), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n283), .A2(KEYINPUT64), .A3(new_n284), .A4(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n284), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n277), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n279), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n264), .B1(new_n275), .B2(new_n289), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n266), .A2(G137), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT66), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n273), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n268), .A2(KEYINPUT66), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n293), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT1), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G128), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n297), .A2(new_n281), .A3(G146), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n190), .A2(new_n212), .A3(G143), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n298), .B(new_n299), .C1(new_n283), .C2(new_n297), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n295), .A2(new_n300), .A3(new_n274), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n302));
  AOI22_X1  g116(.A1(new_n302), .A2(new_n276), .B1(new_n277), .B2(new_n287), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n272), .A2(new_n274), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n303), .A2(new_n304), .A3(KEYINPUT65), .A4(new_n286), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n290), .A2(new_n301), .A3(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT30), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT2), .ZN(new_n309));
  INV_X1    g123(.A(G113), .ZN(new_n310));
  OAI21_X1  g124(.A(KEYINPUT67), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT67), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(KEYINPUT2), .A3(G113), .ZN(new_n313));
  AOI22_X1  g127(.A1(new_n311), .A2(new_n313), .B1(new_n309), .B2(new_n310), .ZN(new_n314));
  XNOR2_X1  g128(.A(G116), .B(G119), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n314), .B(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n289), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n304), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(KEYINPUT30), .A3(new_n301), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n308), .A2(new_n316), .A3(new_n319), .ZN(new_n320));
  XOR2_X1   g134(.A(KEYINPUT26), .B(G101), .Z(new_n321));
  NOR2_X1   g135(.A1(G237), .A2(G953), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G210), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n321), .B(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n324), .B(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n311), .A2(new_n313), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n309), .A2(new_n310), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n327), .A2(new_n328), .A3(new_n315), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n315), .B1(new_n327), .B2(new_n328), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n331), .B(new_n301), .C1(new_n275), .C2(new_n289), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT68), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT68), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n318), .A2(new_n334), .A3(new_n331), .A4(new_n301), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n326), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  AND3_X1   g150(.A1(new_n320), .A2(KEYINPUT70), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT70), .B1(new_n320), .B2(new_n336), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT31), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n333), .A2(new_n335), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n306), .A2(new_n316), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT28), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT28), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n332), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n326), .B(KEYINPUT71), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT31), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n320), .A2(new_n350), .A3(new_n336), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n339), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(G472), .A2(G902), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n352), .A2(KEYINPUT32), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(KEYINPUT32), .B1(new_n352), .B2(new_n353), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT29), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n326), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n331), .B1(new_n318), .B2(new_n301), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n359), .B1(new_n333), .B2(new_n335), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n345), .B(new_n358), .C1(new_n360), .C2(new_n344), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n361), .A2(KEYINPUT73), .A3(new_n250), .ZN(new_n362));
  AOI21_X1  g176(.A(KEYINPUT73), .B1(new_n361), .B2(new_n250), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI22_X1  g178(.A1(new_n333), .A2(new_n335), .B1(new_n306), .B2(new_n316), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n347), .B(new_n345), .C1(new_n365), .C2(new_n344), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT72), .ZN(new_n367));
  AOI21_X1  g181(.A(KEYINPUT29), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n343), .A2(KEYINPUT72), .A3(new_n345), .A4(new_n347), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n320), .A2(new_n340), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n326), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n368), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n364), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G472), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n263), .B1(new_n356), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT88), .B1(new_n216), .B2(new_n225), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n214), .B1(new_n220), .B2(G146), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n211), .A2(KEYINPUT76), .A3(new_n212), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT88), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n379), .A2(new_n380), .A3(new_n224), .A4(new_n222), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT17), .ZN(new_n382));
  INV_X1    g196(.A(G237), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(new_n243), .A3(G214), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(KEYINPUT87), .A3(new_n281), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n281), .A2(KEYINPUT87), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(G214), .A3(new_n322), .ZN(new_n387));
  AOI211_X1 g201(.A(new_n382), .B(new_n273), .C1(new_n385), .C2(new_n387), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n385), .A2(new_n273), .A3(new_n387), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n273), .B1(new_n385), .B2(new_n387), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n388), .B1(new_n391), .B2(new_n382), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n376), .A2(new_n381), .A3(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(G113), .B(G122), .ZN(new_n394));
  INV_X1    g208(.A(G104), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n394), .B(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n385), .A2(new_n387), .ZN(new_n397));
  NAND2_X1  g211(.A1(KEYINPUT18), .A2(G131), .ZN(new_n398));
  XOR2_X1   g212(.A(new_n397), .B(new_n398), .Z(new_n399));
  NOR2_X1   g213(.A1(new_n228), .A2(new_n230), .ZN(new_n400));
  INV_X1    g214(.A(new_n219), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n400), .B1(G146), .B2(new_n401), .ZN(new_n402));
  OR2_X1    g216(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  AND3_X1   g217(.A1(new_n393), .A2(new_n396), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n396), .B1(new_n393), .B2(new_n403), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n250), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT90), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI211_X1 g222(.A(KEYINPUT90), .B(new_n250), .C1(new_n404), .C2(new_n405), .ZN(new_n409));
  XNOR2_X1  g223(.A(KEYINPUT89), .B(G475), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n408), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n393), .A2(new_n396), .A3(new_n403), .ZN(new_n413));
  INV_X1    g227(.A(new_n396), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n219), .B(KEYINPUT19), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n223), .B1(new_n416), .B2(G146), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n417), .A2(new_n391), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n399), .A2(new_n402), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n414), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n413), .A2(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(G475), .A2(G902), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(KEYINPUT20), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT20), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n421), .A2(new_n425), .A3(new_n422), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n412), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(G116), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(KEYINPUT14), .A3(G122), .ZN(new_n430));
  INV_X1    g244(.A(G122), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(G116), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n429), .A2(G122), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  OAI211_X1 g248(.A(G107), .B(new_n430), .C1(new_n434), .C2(KEYINPUT14), .ZN(new_n435));
  INV_X1    g249(.A(G107), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n432), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n190), .A2(G143), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n281), .A2(G128), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n266), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n438), .A2(new_n439), .A3(new_n266), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n435), .B(new_n437), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(KEYINPUT9), .B(G234), .ZN(new_n443));
  NOR3_X1   g257(.A1(new_n443), .A2(new_n257), .A3(G953), .ZN(new_n444));
  OR2_X1    g258(.A1(new_n439), .A2(KEYINPUT13), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n438), .A2(new_n439), .A3(KEYINPUT13), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(G134), .A3(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT92), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n441), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n445), .A2(KEYINPUT92), .A3(new_n446), .A4(G134), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n434), .A2(G107), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n437), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT91), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT91), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n453), .A2(new_n437), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n442), .B(new_n444), .C1(new_n452), .C2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n441), .B1(new_n447), .B2(new_n448), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n461), .A2(new_n451), .A3(new_n455), .A4(new_n457), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n444), .B1(new_n462), .B2(new_n442), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n250), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT93), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(G478), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n467), .A2(KEYINPUT15), .ZN(new_n468));
  OAI211_X1 g282(.A(KEYINPUT93), .B(new_n250), .C1(new_n460), .C2(new_n463), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n466), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  OR2_X1    g284(.A1(new_n464), .A2(new_n468), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(G952), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n473), .A2(G953), .ZN(new_n474));
  NAND2_X1  g288(.A1(G234), .A2(G237), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n476), .B(KEYINPUT94), .ZN(new_n477));
  XOR2_X1   g291(.A(KEYINPUT21), .B(G898), .Z(new_n478));
  NAND3_X1  g292(.A1(new_n475), .A2(G902), .A3(G953), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n428), .A2(new_n472), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(G469), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n436), .A2(G104), .ZN(new_n484));
  AND2_X1   g298(.A1(KEYINPUT82), .A2(KEYINPUT3), .ZN(new_n485));
  NOR2_X1   g299(.A1(KEYINPUT82), .A2(KEYINPUT3), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G101), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n395), .A2(G107), .ZN(new_n489));
  NAND2_X1  g303(.A1(KEYINPUT82), .A2(KEYINPUT3), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n490), .A2(G104), .A3(new_n436), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n487), .A2(new_n488), .A3(new_n489), .A4(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n489), .A2(new_n484), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(G101), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(KEYINPUT84), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT84), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n496), .A2(new_n300), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT10), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n497), .B1(new_n492), .B2(new_n494), .ZN(new_n502));
  INV_X1    g316(.A(new_n300), .ZN(new_n503));
  INV_X1    g317(.A(new_n498), .ZN(new_n504));
  NOR3_X1   g318(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT10), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n487), .A2(new_n489), .A3(new_n491), .ZN(new_n507));
  AND2_X1   g321(.A1(KEYINPUT83), .A2(G101), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(KEYINPUT4), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n492), .ZN(new_n510));
  AOI21_X1  g324(.A(KEYINPUT4), .B1(new_n507), .B2(new_n508), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n317), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n501), .A2(new_n506), .A3(new_n275), .A4(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n300), .B1(new_n496), .B2(new_n498), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n304), .B1(new_n514), .B2(new_n505), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT12), .ZN(new_n516));
  XNOR2_X1  g330(.A(G110), .B(G140), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n243), .A2(G227), .ZN(new_n518));
  XOR2_X1   g332(.A(new_n517), .B(new_n518), .Z(new_n519));
  INV_X1    g333(.A(KEYINPUT12), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n520), .B(new_n304), .C1(new_n514), .C2(new_n505), .ZN(new_n521));
  AND4_X1   g335(.A1(new_n513), .A2(new_n516), .A3(new_n519), .A4(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n512), .B1(new_n505), .B2(KEYINPUT10), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n499), .A2(new_n500), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n304), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n519), .B1(new_n525), .B2(new_n513), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n483), .B(new_n250), .C1(new_n522), .C2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(G469), .A2(G902), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n516), .A2(new_n513), .A3(new_n521), .ZN(new_n529));
  INV_X1    g343(.A(new_n519), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n525), .A2(new_n513), .A3(new_n519), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n527), .B(new_n528), .C1(new_n483), .C2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(G221), .B1(new_n443), .B2(G902), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(G214), .B1(G237), .B2(G902), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n316), .B1(new_n510), .B2(new_n511), .ZN(new_n539));
  NOR3_X1   g353(.A1(new_n429), .A2(KEYINPUT5), .A3(G119), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n540), .B1(new_n315), .B2(KEYINPUT5), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n541), .A2(G113), .B1(new_n314), .B2(new_n315), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n496), .A2(new_n498), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  XOR2_X1   g358(.A(G110), .B(G122), .Z(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n545), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n539), .A2(new_n543), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n546), .A2(KEYINPUT6), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n300), .A2(new_n217), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n550), .B1(new_n289), .B2(new_n217), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n243), .A2(G224), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n551), .B(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n547), .B1(new_n539), .B2(new_n543), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT85), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT6), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n555), .B1(new_n554), .B2(new_n556), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n549), .B(new_n553), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n552), .A2(KEYINPUT7), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n551), .B(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n502), .A2(new_n504), .ZN(new_n562));
  XOR2_X1   g376(.A(new_n562), .B(new_n542), .Z(new_n563));
  XNOR2_X1  g377(.A(new_n545), .B(KEYINPUT8), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n548), .B(new_n561), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n559), .A2(new_n250), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(G210), .B1(G237), .B2(G902), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n559), .A2(new_n565), .A3(new_n250), .A4(new_n567), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n538), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OR2_X1    g385(.A1(new_n571), .A2(KEYINPUT86), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(KEYINPUT86), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n536), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n375), .A2(new_n482), .A3(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(G101), .ZN(G3));
  NAND2_X1  g390(.A1(new_n352), .A2(new_n250), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(G472), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(KEYINPUT95), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n352), .A2(new_n353), .ZN(new_n580));
  INV_X1    g394(.A(G472), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n581), .B1(new_n352), .B2(new_n250), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT95), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n580), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NOR4_X1   g398(.A1(new_n579), .A2(new_n584), .A3(new_n263), .A4(new_n536), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n466), .A2(new_n467), .A3(new_n469), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n460), .A2(new_n463), .A3(KEYINPUT33), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT33), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n442), .B1(new_n452), .B2(new_n458), .ZN(new_n589));
  INV_X1    g403(.A(new_n444), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n588), .B1(new_n591), .B2(new_n459), .ZN(new_n592));
  OAI211_X1 g406(.A(G478), .B(new_n250), .C1(new_n587), .C2(new_n592), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n586), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n594), .B1(new_n412), .B2(new_n427), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n571), .A2(new_n480), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n585), .A2(new_n596), .ZN(new_n597));
  XOR2_X1   g411(.A(KEYINPUT34), .B(G104), .Z(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(G6));
  AOI21_X1  g413(.A(new_n410), .B1(new_n406), .B2(new_n407), .ZN(new_n600));
  AOI22_X1  g414(.A1(new_n600), .A2(new_n409), .B1(new_n471), .B2(new_n470), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT96), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n424), .A2(new_n602), .A3(new_n426), .ZN(new_n603));
  OR2_X1    g417(.A1(new_n426), .A2(new_n602), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AND4_X1   g419(.A1(new_n480), .A2(new_n571), .A3(new_n601), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n585), .A2(new_n606), .ZN(new_n607));
  XOR2_X1   g421(.A(KEYINPUT35), .B(G107), .Z(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT97), .B(KEYINPUT98), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G9));
  NOR2_X1   g425(.A1(new_n579), .A2(new_n584), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n245), .A2(KEYINPUT36), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n240), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n261), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n259), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n574), .A2(new_n612), .A3(new_n482), .A4(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(KEYINPUT37), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(new_n198), .ZN(G12));
  INV_X1    g433(.A(KEYINPUT99), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n412), .A2(new_n603), .A3(new_n472), .A4(new_n604), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n477), .B1(G900), .B2(new_n479), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n620), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n569), .A2(new_n570), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n625), .A2(new_n537), .A3(new_n616), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n605), .A2(KEYINPUT99), .A3(new_n601), .A4(new_n622), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n624), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n536), .B1(new_n356), .B2(new_n374), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(G128), .ZN(G30));
  XNOR2_X1  g445(.A(new_n625), .B(KEYINPUT100), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT38), .ZN(new_n633));
  OR2_X1    g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(new_n616), .ZN(new_n637));
  XOR2_X1   g451(.A(new_n622), .B(KEYINPUT39), .Z(new_n638));
  OR2_X1    g452(.A1(new_n536), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(new_n639), .B(KEYINPUT40), .Z(new_n640));
  NAND3_X1  g454(.A1(new_n428), .A2(new_n472), .A3(new_n537), .ZN(new_n641));
  INV_X1    g455(.A(new_n338), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n320), .A2(KEYINPUT70), .A3(new_n336), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n645));
  OR2_X1    g459(.A1(new_n347), .A2(new_n360), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n250), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n645), .B1(new_n644), .B2(new_n646), .ZN(new_n649));
  OAI21_X1  g463(.A(G472), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n641), .B1(new_n356), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n637), .A2(new_n640), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G143), .ZN(G45));
  AOI22_X1  g467(.A1(new_n600), .A2(new_n409), .B1(new_n424), .B2(new_n426), .ZN(new_n654));
  NOR4_X1   g468(.A1(new_n654), .A2(KEYINPUT102), .A3(new_n594), .A4(new_n623), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT102), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n656), .B1(new_n595), .B2(new_n622), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT32), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n580), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n352), .A2(KEYINPUT32), .A3(new_n353), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n660), .A2(new_n374), .A3(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n536), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n658), .A2(new_n662), .A3(new_n663), .A4(new_n626), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G146), .ZN(G48));
  INV_X1    g479(.A(KEYINPUT104), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n250), .B1(new_n522), .B2(new_n526), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(G469), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n668), .A2(new_n535), .A3(new_n527), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT103), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n668), .A2(KEYINPUT103), .A3(new_n535), .A4(new_n527), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n375), .A2(new_n666), .A3(new_n596), .A4(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n263), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n673), .A2(new_n662), .A3(new_n596), .A4(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(KEYINPUT104), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT41), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G113), .ZN(G15));
  NAND4_X1  g494(.A1(new_n606), .A2(new_n673), .A3(new_n675), .A4(new_n662), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G116), .ZN(G18));
  NAND4_X1  g496(.A1(new_n673), .A2(new_n662), .A3(new_n482), .A4(new_n626), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G119), .ZN(G21));
  INV_X1    g498(.A(new_n625), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n641), .A2(new_n685), .A3(new_n481), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n345), .B1(new_n360), .B2(new_n344), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n348), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n339), .A2(new_n351), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n353), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n691), .A2(new_n582), .A3(new_n263), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n686), .A2(new_n692), .A3(new_n673), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G122), .ZN(G24));
  NAND3_X1  g508(.A1(new_n578), .A2(new_n616), .A3(new_n690), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n671), .A2(new_n571), .A3(new_n672), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n658), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G125), .ZN(G27));
  INV_X1    g513(.A(KEYINPUT42), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n529), .A2(new_n701), .A3(new_n530), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n701), .B1(new_n529), .B2(new_n530), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n525), .A2(new_n513), .A3(new_n519), .ZN(new_n705));
  NOR4_X1   g519(.A1(new_n703), .A2(new_n704), .A3(new_n483), .A4(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n527), .A2(new_n528), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n535), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n569), .A2(new_n537), .A3(new_n570), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n662), .A2(new_n710), .A3(new_n675), .ZN(new_n711));
  INV_X1    g525(.A(new_n657), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n595), .A2(new_n656), .A3(new_n622), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n700), .B1(new_n711), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(KEYINPUT106), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT106), .ZN(new_n717));
  OAI211_X1 g531(.A(new_n717), .B(new_n700), .C1(new_n711), .C2(new_n714), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n660), .A2(new_n720), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n374), .B(new_n721), .C1(new_n356), .C2(new_n720), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n722), .A2(new_n675), .ZN(new_n723));
  INV_X1    g537(.A(new_n535), .ZN(new_n724));
  INV_X1    g538(.A(new_n707), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n531), .A2(KEYINPUT105), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n726), .A2(G469), .A3(new_n532), .A4(new_n702), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n724), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n714), .A2(new_n709), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n723), .A2(KEYINPUT42), .A3(new_n728), .A4(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n719), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G131), .ZN(G33));
  NAND2_X1  g546(.A1(new_n624), .A2(new_n627), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n375), .A2(new_n734), .A3(KEYINPUT108), .A4(new_n710), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT108), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n736), .B1(new_n711), .B2(new_n733), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n266), .ZN(G36));
  INV_X1    g553(.A(KEYINPUT45), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n533), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n726), .A2(new_n532), .A3(new_n702), .ZN(new_n742));
  OAI211_X1 g556(.A(G469), .B(new_n741), .C1(new_n742), .C2(new_n740), .ZN(new_n743));
  AOI21_X1  g557(.A(KEYINPUT46), .B1(new_n743), .B2(new_n528), .ZN(new_n744));
  INV_X1    g558(.A(new_n527), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n743), .A2(KEYINPUT46), .A3(new_n528), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n535), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT44), .ZN(new_n750));
  INV_X1    g564(.A(new_n612), .ZN(new_n751));
  INV_X1    g565(.A(new_n594), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n654), .A2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT43), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n751), .A2(new_n755), .A3(new_n616), .ZN(new_n756));
  AOI211_X1 g570(.A(new_n638), .B(new_n749), .C1(new_n750), .C2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n756), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n709), .B1(new_n758), .B2(KEYINPUT44), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(KEYINPUT109), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(new_n269), .ZN(G39));
  INV_X1    g576(.A(KEYINPUT47), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n749), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n748), .A2(KEYINPUT47), .A3(new_n535), .ZN(new_n765));
  AOI211_X1 g579(.A(new_n714), .B(new_n709), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n662), .A2(new_n675), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G140), .ZN(G42));
  NAND2_X1  g583(.A1(new_n675), .A2(new_n537), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n668), .A2(new_n527), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n771), .A2(KEYINPUT49), .ZN(new_n772));
  NOR4_X1   g586(.A1(new_n770), .A2(new_n772), .A3(new_n724), .A4(new_n753), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(KEYINPUT110), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n650), .A2(new_n660), .A3(new_n661), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n771), .A2(KEYINPUT49), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(KEYINPUT111), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n774), .A2(new_n636), .A3(new_n776), .A4(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n634), .A2(new_n635), .A3(new_n538), .ZN(new_n780));
  INV_X1    g594(.A(new_n477), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n755), .A2(new_n781), .A3(new_n673), .A4(new_n692), .ZN(new_n782));
  OR2_X1    g596(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n783));
  OR3_X1    g597(.A1(new_n780), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n709), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n673), .A2(new_n785), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n786), .A2(new_n755), .A3(new_n781), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n696), .ZN(new_n788));
  NAND2_X1  g602(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n783), .B(new_n789), .C1(new_n780), .C2(new_n782), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n263), .A2(new_n477), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n428), .A2(new_n752), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n786), .A2(new_n776), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n784), .A2(new_n788), .A3(new_n790), .A4(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n764), .A2(new_n765), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n668), .A2(new_n724), .A3(new_n527), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n755), .A2(new_n781), .A3(new_n692), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n785), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n795), .A2(new_n802), .A3(KEYINPUT51), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n474), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT51), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n800), .B1(new_n796), .B2(new_n797), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n805), .B1(new_n794), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  OAI211_X1 g623(.A(KEYINPUT117), .B(new_n805), .C1(new_n794), .C2(new_n806), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n804), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n738), .B1(new_n719), .B2(new_n730), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT52), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n630), .A2(new_n664), .A3(new_n698), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n616), .A2(new_n623), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n728), .A2(new_n816), .A3(KEYINPUT113), .ZN(new_n817));
  INV_X1    g631(.A(new_n641), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n775), .A2(new_n817), .A3(new_n625), .A4(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT113), .B1(new_n728), .B2(new_n816), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n814), .B1(new_n815), .B2(new_n821), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n695), .A2(new_n655), .A3(new_n657), .ZN(new_n823));
  AOI22_X1  g637(.A1(new_n697), .A2(new_n823), .B1(new_n628), .B2(new_n629), .ZN(new_n824));
  INV_X1    g638(.A(new_n820), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n651), .A2(new_n825), .A3(new_n625), .A4(new_n817), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n824), .A2(KEYINPUT52), .A3(new_n664), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n822), .A2(new_n827), .ZN(new_n828));
  AND4_X1   g642(.A1(new_n471), .A2(new_n605), .A3(new_n470), .A4(new_n622), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n629), .A2(new_n412), .A3(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n658), .A2(new_n578), .A3(new_n690), .A4(new_n728), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n709), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(new_n616), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n813), .A2(new_n828), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n572), .A2(new_n573), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n654), .A2(new_n472), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n836), .B1(new_n654), .B2(new_n594), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n585), .A2(new_n480), .A3(new_n835), .A4(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n838), .A2(new_n575), .A3(new_n617), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n681), .A2(new_n683), .A3(new_n693), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n678), .A2(new_n841), .A3(KEYINPUT112), .ZN(new_n842));
  AOI21_X1  g656(.A(KEYINPUT112), .B1(new_n678), .B2(new_n841), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n840), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n812), .B1(new_n834), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n678), .A2(new_n841), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT112), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n678), .A2(new_n841), .A3(KEYINPUT112), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n839), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI22_X1  g664(.A1(new_n822), .A2(new_n827), .B1(new_n616), .B2(new_n832), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n850), .A2(KEYINPUT53), .A3(new_n813), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n845), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT54), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n786), .A2(new_n595), .A3(new_n776), .A4(new_n791), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n846), .A2(KEYINPUT114), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT114), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n678), .A2(new_n841), .A3(new_n857), .ZN(new_n858));
  AOI22_X1  g672(.A1(new_n856), .A2(new_n858), .B1(new_n822), .B2(new_n827), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n812), .B1(new_n832), .B2(new_n616), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n859), .A2(new_n813), .A3(new_n840), .A4(new_n860), .ZN(new_n861));
  XNOR2_X1  g675(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n845), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n811), .A2(new_n854), .A3(new_n855), .A4(new_n863), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n799), .A2(new_n697), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n787), .A2(new_n723), .ZN(new_n866));
  XOR2_X1   g680(.A(new_n866), .B(KEYINPUT48), .Z(new_n867));
  NOR3_X1   g681(.A1(new_n864), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(G952), .A2(G953), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n779), .B1(new_n868), .B2(new_n869), .ZN(G75));
  NAND2_X1  g684(.A1(new_n473), .A2(G953), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT119), .Z(new_n872));
  AOI21_X1  g686(.A(new_n250), .B1(new_n845), .B2(new_n861), .ZN(new_n873));
  AOI21_X1  g687(.A(KEYINPUT56), .B1(new_n873), .B2(G210), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n872), .B1(new_n874), .B2(KEYINPUT118), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(KEYINPUT118), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n549), .B1(new_n557), .B2(new_n558), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(new_n553), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT55), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n879), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n874), .A2(KEYINPUT118), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n875), .B1(new_n880), .B2(new_n882), .ZN(G51));
  INV_X1    g697(.A(new_n872), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n522), .A2(new_n526), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n885), .B(KEYINPUT120), .Z(new_n886));
  AND3_X1   g700(.A1(new_n845), .A2(new_n861), .A3(new_n862), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n862), .B1(new_n845), .B2(new_n861), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n528), .B(KEYINPUT57), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n886), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n873), .ZN(new_n892));
  OR2_X1    g706(.A1(new_n892), .A2(new_n743), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n884), .B1(new_n891), .B2(new_n893), .ZN(G54));
  NAND3_X1  g708(.A1(new_n873), .A2(KEYINPUT58), .A3(G475), .ZN(new_n895));
  INV_X1    g709(.A(new_n421), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT121), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n895), .A2(new_n898), .A3(new_n896), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n898), .B1(new_n895), .B2(new_n896), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n872), .B(new_n897), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(G60));
  OR2_X1    g716(.A1(new_n587), .A2(new_n592), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(G478), .A2(G902), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT59), .Z(new_n906));
  NOR2_X1   g720(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n907), .B1(new_n887), .B2(new_n888), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n906), .B1(new_n854), .B2(new_n863), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n872), .B(new_n908), .C1(new_n909), .C2(new_n903), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT54), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n913), .B1(new_n845), .B2(new_n852), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n887), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n904), .B1(new_n915), .B2(new_n906), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n916), .A2(KEYINPUT122), .A3(new_n872), .A4(new_n908), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n912), .A2(new_n917), .ZN(G63));
  NAND2_X1  g732(.A1(new_n845), .A2(new_n861), .ZN(new_n919));
  NAND2_X1  g733(.A1(G217), .A2(G902), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT60), .Z(new_n921));
  NAND3_X1  g735(.A1(new_n919), .A2(new_n614), .A3(new_n921), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n919), .A2(new_n921), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n249), .B(KEYINPUT123), .Z(new_n924));
  OAI211_X1 g738(.A(new_n872), .B(new_n922), .C1(new_n923), .C2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT61), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(G66));
  AOI21_X1  g741(.A(new_n243), .B1(new_n478), .B2(G224), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n928), .B1(new_n844), .B2(new_n243), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n877), .B1(G898), .B2(new_n243), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n929), .B(new_n930), .Z(G69));
  INV_X1    g745(.A(new_n815), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n652), .A2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT62), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n934), .A2(KEYINPUT124), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n652), .A2(new_n932), .A3(new_n935), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI22_X1  g753(.A1(new_n766), .A2(new_n767), .B1(new_n757), .B2(new_n759), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n934), .A2(KEYINPUT124), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n639), .A2(new_n709), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n942), .A2(new_n375), .A3(new_n837), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n939), .A2(new_n940), .A3(new_n941), .A4(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n243), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n308), .A2(new_n319), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(new_n415), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n243), .B1(G227), .B2(G900), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT125), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n947), .ZN(new_n952));
  NAND2_X1  g766(.A1(G900), .A2(G953), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n749), .A2(new_n638), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n954), .A2(new_n625), .A3(new_n818), .A4(new_n723), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n940), .A2(new_n813), .A3(new_n932), .A4(new_n955), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n952), .B(new_n953), .C1(new_n956), .C2(G953), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n948), .A2(new_n951), .A3(new_n957), .ZN(new_n958));
  OR2_X1    g772(.A1(new_n949), .A2(new_n950), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n958), .B(new_n959), .ZN(G72));
  NAND2_X1  g774(.A1(G472), .A2(G902), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT63), .Z(new_n962));
  INV_X1    g776(.A(new_n644), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n371), .B(KEYINPUT127), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n853), .B(new_n962), .C1(new_n963), .C2(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n962), .B1(new_n944), .B2(new_n844), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n370), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n965), .B1(new_n967), .B2(new_n326), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n962), .B1(new_n956), .B2(new_n844), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n969), .A2(new_n340), .A3(new_n326), .A4(new_n320), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n970), .A2(KEYINPUT126), .A3(new_n872), .ZN(new_n971));
  AOI21_X1  g785(.A(KEYINPUT126), .B1(new_n970), .B2(new_n872), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n968), .A2(new_n971), .A3(new_n972), .ZN(G57));
endmodule


