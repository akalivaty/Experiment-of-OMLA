//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 1 0 0 0 1 1 0 0 1 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:10 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998;
  INV_X1    g000(.A(KEYINPUT4), .ZN(new_n187));
  INV_X1    g001(.A(G107), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(KEYINPUT74), .A3(G104), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  NAND4_X1  g005(.A1(new_n188), .A2(KEYINPUT74), .A3(KEYINPUT3), .A4(G104), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT75), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n193), .B1(new_n188), .B2(G104), .ZN(new_n194));
  INV_X1    g008(.A(G104), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(KEYINPUT75), .A3(G107), .ZN(new_n196));
  AOI22_X1  g010(.A1(new_n191), .A2(new_n192), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G101), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n187), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n194), .A2(new_n196), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n195), .A2(G107), .ZN(new_n201));
  AOI21_X1  g015(.A(KEYINPUT3), .B1(new_n201), .B2(KEYINPUT74), .ZN(new_n202));
  INV_X1    g016(.A(new_n192), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n200), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G101), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n199), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT2), .B(G113), .ZN(new_n207));
  XNOR2_X1  g021(.A(G116), .B(G119), .ZN(new_n208));
  XNOR2_X1  g022(.A(new_n207), .B(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n204), .A2(new_n187), .A3(G101), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n206), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n198), .B(new_n200), .C1(new_n202), .C2(new_n203), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT5), .ZN(new_n214));
  INV_X1    g028(.A(G119), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(new_n215), .A3(G116), .ZN(new_n216));
  XOR2_X1   g030(.A(G116), .B(G119), .Z(new_n217));
  OAI211_X1 g031(.A(G113), .B(new_n216), .C1(new_n217), .C2(new_n214), .ZN(new_n218));
  OR2_X1    g032(.A1(new_n217), .A2(new_n207), .ZN(new_n219));
  INV_X1    g033(.A(new_n201), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n195), .A2(G107), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n198), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n213), .A2(new_n218), .A3(new_n219), .A4(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n212), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n213), .A2(new_n223), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n218), .A2(new_n219), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(new_n224), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT8), .ZN(new_n230));
  XOR2_X1   g044(.A(G110), .B(G122), .Z(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n225), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n229), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n231), .B1(new_n234), .B2(KEYINPUT8), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(G143), .B(G146), .ZN(new_n237));
  XNOR2_X1  g051(.A(KEYINPUT0), .B(G128), .ZN(new_n238));
  OAI21_X1  g052(.A(KEYINPUT64), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n237), .A2(KEYINPUT0), .A3(G128), .ZN(new_n240));
  INV_X1    g054(.A(G146), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G143), .ZN(new_n242));
  INV_X1    g056(.A(G143), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G146), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G128), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT0), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT0), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G128), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT64), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n245), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n239), .A2(new_n240), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G125), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n243), .A2(G146), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n241), .A2(G143), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n246), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(KEYINPUT1), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT1), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n242), .A2(new_n244), .A3(new_n259), .A4(G128), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n257), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G125), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n254), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G953), .ZN(new_n265));
  XOR2_X1   g079(.A(KEYINPUT78), .B(G224), .Z(new_n266));
  NAND3_X1  g080(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n265), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n254), .A2(new_n263), .A3(KEYINPUT7), .A4(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT79), .ZN(new_n270));
  AND4_X1   g084(.A1(new_n262), .A2(new_n257), .A3(new_n258), .A4(new_n260), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n271), .B1(G125), .B2(new_n253), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT79), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n272), .A2(new_n273), .A3(KEYINPUT7), .A4(new_n268), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT7), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n264), .A2(new_n275), .ZN(new_n276));
  AND4_X1   g090(.A1(new_n267), .A2(new_n270), .A3(new_n274), .A4(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(G902), .B1(new_n236), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n225), .A2(new_n231), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n212), .A2(new_n224), .A3(new_n232), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n281), .A2(KEYINPUT77), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n279), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n272), .A2(new_n268), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n267), .A2(new_n284), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n225), .B(new_n231), .C1(KEYINPUT77), .C2(new_n281), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n283), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n278), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(G210), .B1(G237), .B2(G902), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT80), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n278), .A2(new_n289), .A3(new_n287), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(G214), .B1(G237), .B2(G902), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n278), .A2(KEYINPUT80), .A3(new_n287), .A4(new_n289), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G140), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n262), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(G125), .A2(G140), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n301), .B(new_n241), .ZN(new_n302));
  INV_X1    g116(.A(G237), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(new_n265), .A3(G214), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n243), .ZN(new_n305));
  NOR2_X1   g119(.A1(G237), .A2(G953), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n306), .A2(G143), .A3(G214), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(KEYINPUT18), .A3(G131), .ZN(new_n309));
  AND2_X1   g123(.A1(KEYINPUT18), .A2(G131), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n302), .B(new_n309), .C1(new_n308), .C2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT19), .ZN(new_n312));
  AND2_X1   g126(.A1(G125), .A2(G140), .ZN(new_n313));
  NOR2_X1   g127(.A1(G125), .A2(G140), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n299), .A2(KEYINPUT19), .A3(new_n300), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(new_n316), .A3(new_n241), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT16), .B1(new_n313), .B2(new_n314), .ZN(new_n318));
  OR3_X1    g132(.A1(new_n262), .A2(KEYINPUT16), .A3(G140), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(new_n319), .A3(G146), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n317), .A2(new_n320), .A3(KEYINPUT82), .ZN(new_n321));
  AND4_X1   g135(.A1(G143), .A2(new_n303), .A3(new_n265), .A4(G214), .ZN(new_n322));
  AOI21_X1  g136(.A(G143), .B1(new_n306), .B2(G214), .ZN(new_n323));
  OAI21_X1  g137(.A(G131), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G131), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n305), .A2(new_n325), .A3(new_n307), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n321), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(KEYINPUT82), .B1(new_n317), .B2(new_n320), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n311), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(G113), .B(G122), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n331), .B(new_n195), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT17), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n324), .A2(new_n335), .A3(new_n326), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n318), .A2(new_n319), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n241), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n308), .A2(KEYINPUT17), .A3(G131), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n336), .A2(new_n338), .A3(new_n320), .A4(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(new_n332), .A3(new_n311), .ZN(new_n341));
  AOI21_X1  g155(.A(KEYINPUT20), .B1(new_n334), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g156(.A1(G475), .A2(G902), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n342), .A2(KEYINPUT84), .A3(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT20), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n317), .A2(new_n320), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT82), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(new_n327), .A3(new_n321), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n332), .B1(new_n349), .B2(new_n311), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n340), .A2(new_n332), .A3(new_n311), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n345), .B(new_n343), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT84), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n343), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT83), .B1(new_n350), .B2(new_n351), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT83), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n334), .A2(new_n357), .A3(new_n341), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n355), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(KEYINPUT81), .B(KEYINPUT20), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n344), .B(new_n354), .C1(new_n359), .C2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n332), .B1(new_n340), .B2(new_n311), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT85), .ZN(new_n364));
  INV_X1    g178(.A(G902), .ZN(new_n365));
  OR2_X1    g179(.A1(new_n351), .A2(KEYINPUT85), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n364), .B(new_n365), .C1(new_n366), .C2(new_n363), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G475), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n362), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT86), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n362), .A2(KEYINPUT86), .A3(new_n368), .ZN(new_n372));
  AND2_X1   g186(.A1(KEYINPUT87), .A2(G122), .ZN(new_n373));
  NOR2_X1   g187(.A1(KEYINPUT87), .A2(G122), .ZN(new_n374));
  OAI21_X1  g188(.A(G116), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G116), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G122), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n375), .A2(new_n188), .A3(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(G128), .B(G143), .ZN(new_n379));
  INV_X1    g193(.A(G134), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n379), .B(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G122), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT14), .B1(new_n382), .B2(G116), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT88), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n377), .A2(KEYINPUT88), .A3(KEYINPUT14), .ZN(new_n386));
  OR3_X1    g200(.A1(new_n382), .A2(KEYINPUT14), .A3(G116), .ZN(new_n387));
  AND4_X1   g201(.A1(new_n375), .A2(new_n385), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n378), .B(new_n381), .C1(new_n388), .C2(new_n188), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n379), .A2(KEYINPUT13), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n243), .A2(G128), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n390), .B(G134), .C1(KEYINPUT13), .C2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n379), .A2(new_n380), .ZN(new_n393));
  INV_X1    g207(.A(new_n378), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n188), .B1(new_n375), .B2(new_n377), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n392), .B(new_n393), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(KEYINPUT9), .B(G234), .ZN(new_n397));
  INV_X1    g211(.A(G217), .ZN(new_n398));
  NOR3_X1   g212(.A1(new_n397), .A2(new_n398), .A3(G953), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n389), .A2(new_n396), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n399), .B1(new_n389), .B2(new_n396), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n365), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G478), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(KEYINPUT15), .ZN(new_n404));
  OR2_X1    g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n402), .A2(new_n404), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G952), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(G953), .ZN(new_n409));
  NAND2_X1  g223(.A1(G234), .A2(G237), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  XOR2_X1   g226(.A(KEYINPUT21), .B(G898), .Z(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n410), .A2(G902), .A3(G953), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n412), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n407), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n371), .A2(new_n372), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(G469), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT76), .ZN(new_n423));
  AOI21_X1  g237(.A(G128), .B1(new_n242), .B2(new_n244), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n244), .A2(new_n259), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n258), .B(KEYINPUT76), .C1(new_n237), .C2(G128), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n260), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n222), .B1(new_n197), .B2(new_n198), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n226), .A2(new_n261), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT11), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n433), .B1(new_n380), .B2(G137), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n380), .A2(G137), .ZN(new_n435));
  INV_X1    g249(.A(G137), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n436), .A2(KEYINPUT11), .A3(G134), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n434), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G131), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n434), .A2(new_n437), .A3(new_n325), .A4(new_n435), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(KEYINPUT12), .B1(new_n432), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT12), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n439), .A2(new_n440), .ZN(new_n444));
  AOI211_X1 g258(.A(new_n443), .B(new_n444), .C1(new_n430), .C2(new_n431), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n253), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n206), .A2(new_n447), .A3(new_n211), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT10), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n430), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n257), .A2(new_n258), .A3(new_n260), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n429), .A2(KEYINPUT10), .A3(new_n451), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n448), .A2(new_n450), .A3(new_n444), .A4(new_n452), .ZN(new_n453));
  XOR2_X1   g267(.A(G110), .B(G140), .Z(new_n454));
  XNOR2_X1  g268(.A(KEYINPUT72), .B(KEYINPUT73), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n454), .B(new_n455), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n265), .A2(G227), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n456), .B(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n446), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n448), .A2(new_n450), .A3(new_n452), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n441), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n458), .B1(new_n462), .B2(new_n453), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n422), .B(new_n365), .C1(new_n460), .C2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n453), .B1(new_n442), .B2(new_n445), .ZN(new_n465));
  INV_X1    g279(.A(new_n458), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n453), .A2(new_n458), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n462), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n467), .A2(new_n469), .A3(G469), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n422), .A2(new_n365), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n464), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(G221), .B1(new_n397), .B2(G902), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n297), .A2(new_n421), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n435), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n380), .A2(G137), .ZN(new_n478));
  OAI21_X1  g292(.A(G131), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n451), .A2(new_n440), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT30), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n480), .B(new_n481), .C1(new_n444), .C2(new_n253), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n441), .A2(new_n240), .A3(new_n252), .A4(new_n239), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n481), .B1(new_n484), .B2(new_n480), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n210), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n480), .B(new_n209), .C1(new_n444), .C2(new_n253), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  XOR2_X1   g302(.A(KEYINPUT26), .B(G101), .Z(new_n489));
  XNOR2_X1  g303(.A(KEYINPUT65), .B(KEYINPUT27), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n489), .B(new_n490), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n306), .A2(G210), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n491), .B(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(KEYINPUT29), .B1(new_n488), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT28), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n480), .B1(new_n444), .B2(new_n253), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n210), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n495), .B1(new_n497), .B2(new_n487), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n487), .A2(new_n495), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(KEYINPUT66), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n487), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n209), .B1(new_n484), .B2(new_n480), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT28), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT66), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n494), .B1(new_n507), .B2(new_n493), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT67), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n497), .A2(new_n509), .A3(new_n487), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n503), .A2(KEYINPUT67), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(KEYINPUT28), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n493), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n512), .A2(KEYINPUT29), .A3(new_n499), .A4(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n508), .A2(new_n365), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(G472), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT32), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n486), .A2(new_n487), .A3(new_n513), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT31), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n496), .A2(KEYINPUT30), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n482), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n502), .B1(new_n522), .B2(new_n210), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n523), .A2(KEYINPUT31), .A3(new_n513), .ZN(new_n524));
  AOI22_X1  g338(.A1(new_n507), .A2(new_n493), .B1(new_n520), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(G472), .A2(G902), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n517), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(KEYINPUT31), .B1(new_n523), .B2(new_n513), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n209), .B1(new_n521), .B2(new_n482), .ZN(new_n530));
  NOR4_X1   g344(.A1(new_n530), .A2(new_n519), .A3(new_n502), .A4(new_n493), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n513), .B1(new_n501), .B2(new_n506), .ZN(new_n533));
  OAI211_X1 g347(.A(KEYINPUT32), .B(new_n526), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n516), .A2(new_n528), .A3(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n265), .A2(G221), .A3(G234), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(G137), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT69), .B(KEYINPUT22), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n537), .B(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n215), .A2(G128), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n540), .B1(KEYINPUT68), .B2(KEYINPUT23), .ZN(new_n541));
  OR2_X1    g355(.A1(new_n540), .A2(KEYINPUT68), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n246), .A2(G119), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT23), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n541), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n540), .A2(new_n543), .ZN(new_n547));
  XOR2_X1   g361(.A(KEYINPUT24), .B(G110), .Z(new_n548));
  OAI22_X1  g362(.A1(new_n546), .A2(G110), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n301), .A2(new_n241), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(new_n320), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n546), .A2(G110), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n338), .A2(new_n320), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n547), .A2(new_n548), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n539), .B1(new_n551), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n551), .A2(new_n555), .A3(new_n539), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n398), .B1(G234), .B2(new_n365), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n560), .A2(G902), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n562), .B(KEYINPUT71), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT25), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT70), .ZN(new_n565));
  INV_X1    g379(.A(new_n558), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n365), .B(new_n565), .C1(new_n566), .C2(new_n556), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n564), .A2(KEYINPUT70), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n568), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n559), .A2(new_n365), .A3(new_n570), .A4(new_n565), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n569), .A2(new_n571), .A3(new_n560), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n563), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n535), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n476), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(G101), .ZN(G3));
  INV_X1    g392(.A(KEYINPUT90), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n291), .A2(new_n579), .A3(new_n295), .ZN(new_n580));
  INV_X1    g394(.A(new_n295), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n581), .A2(KEYINPUT89), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n293), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n289), .B1(new_n278), .B2(new_n287), .ZN(new_n585));
  OAI21_X1  g399(.A(KEYINPUT90), .B1(new_n585), .B2(new_n581), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n580), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n584), .B1(new_n580), .B2(new_n586), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n402), .A2(new_n403), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n400), .A2(new_n401), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n591), .A2(KEYINPUT33), .ZN(new_n592));
  OAI21_X1  g406(.A(KEYINPUT91), .B1(new_n400), .B2(new_n401), .ZN(new_n593));
  OR2_X1    g407(.A1(new_n401), .A2(KEYINPUT91), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(new_n594), .A3(KEYINPUT33), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT92), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n593), .A2(new_n594), .A3(KEYINPUT92), .A4(KEYINPUT33), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n592), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n403), .A2(G902), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n371), .A2(new_n372), .B1(new_n590), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n520), .A2(new_n524), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n505), .B1(new_n504), .B2(new_n499), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n498), .A2(KEYINPUT66), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n493), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(G902), .B1(new_n603), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(G472), .ZN(new_n608));
  OAI22_X1  g422(.A1(new_n607), .A2(new_n608), .B1(new_n525), .B2(new_n527), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n609), .A2(new_n475), .A3(new_n573), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n589), .A2(new_n418), .A3(new_n602), .A4(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT34), .B(G104), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G6));
  AOI21_X1  g427(.A(new_n579), .B1(new_n291), .B2(new_n295), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n585), .A2(KEYINPUT90), .A3(new_n581), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n583), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n580), .A2(new_n584), .A3(new_n586), .ZN(new_n617));
  INV_X1    g431(.A(new_n368), .ZN(new_n618));
  OR2_X1    g432(.A1(new_n359), .A2(new_n361), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n359), .A2(new_n361), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n619), .A2(KEYINPUT93), .A3(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT93), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n359), .A2(new_n361), .ZN(new_n623));
  AOI211_X1 g437(.A(new_n355), .B(new_n360), .C1(new_n356), .C2(new_n358), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  AOI211_X1 g439(.A(new_n618), .B(new_n407), .C1(new_n621), .C2(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n616), .A2(new_n418), .A3(new_n617), .A4(new_n626), .ZN(new_n627));
  AND2_X1   g441(.A1(new_n627), .A2(KEYINPUT94), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n627), .A2(KEYINPUT94), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n610), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT35), .B(G107), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G9));
  NAND2_X1  g446(.A1(new_n551), .A2(new_n555), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n539), .A2(KEYINPUT36), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n561), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n572), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n297), .A2(new_n421), .A3(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n609), .A2(new_n475), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(KEYINPUT37), .B(G110), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT95), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n641), .B(new_n643), .ZN(G12));
  INV_X1    g458(.A(new_n475), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n535), .A2(new_n645), .A3(new_n637), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n589), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n411), .B(KEYINPUT96), .ZN(new_n648));
  INV_X1    g462(.A(G900), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n648), .B1(new_n649), .B2(new_n416), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n626), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT97), .B(G128), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G30));
  XNOR2_X1  g469(.A(new_n650), .B(KEYINPUT39), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n475), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT40), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n637), .A2(new_n581), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n294), .A2(new_n296), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT38), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n294), .A2(KEYINPUT38), .A3(new_n296), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n407), .B1(new_n371), .B2(new_n372), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n510), .A2(new_n493), .A3(new_n511), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n518), .A2(new_n667), .A3(G472), .ZN(new_n668));
  NAND2_X1  g482(.A1(G472), .A2(G902), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n668), .A2(KEYINPUT98), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g484(.A(KEYINPUT98), .B1(new_n668), .B2(new_n669), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n528), .A2(new_n534), .A3(new_n672), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n666), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n659), .A2(new_n660), .A3(new_n665), .A4(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT99), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G143), .ZN(G45));
  NAND2_X1  g491(.A1(new_n371), .A2(new_n372), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n601), .A2(new_n590), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n678), .A2(new_n679), .A3(new_n651), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n647), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(KEYINPUT100), .B(G146), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G48));
  NAND4_X1  g498(.A1(new_n616), .A2(new_n602), .A3(new_n418), .A4(new_n617), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n365), .B1(new_n460), .B2(new_n463), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(G469), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n687), .A2(new_n474), .A3(new_n464), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT101), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n687), .A2(KEYINPUT101), .A3(new_n474), .A4(new_n464), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n692), .A2(new_n535), .A3(new_n574), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n685), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT41), .B(G113), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G15));
  INV_X1    g510(.A(new_n693), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n697), .B1(new_n628), .B2(new_n629), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G116), .ZN(G18));
  NOR3_X1   g513(.A1(new_n587), .A2(new_n588), .A3(new_n688), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT102), .ZN(new_n701));
  INV_X1    g515(.A(new_n372), .ZN(new_n702));
  AOI21_X1  g516(.A(KEYINPUT86), .B1(new_n362), .B2(new_n368), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n702), .A2(new_n703), .A3(new_n419), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n535), .A2(new_n637), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n700), .A2(new_n701), .A3(new_n704), .A4(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n688), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n616), .A2(new_n704), .A3(new_n617), .A4(new_n708), .ZN(new_n709));
  OAI21_X1  g523(.A(KEYINPUT102), .B1(new_n709), .B2(new_n705), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G119), .ZN(G21));
  NAND4_X1  g526(.A1(new_n692), .A2(new_n616), .A3(new_n617), .A4(new_n666), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n607), .A2(new_n608), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n526), .B(KEYINPUT103), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n512), .A2(new_n499), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n493), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n715), .B1(new_n603), .B2(new_n717), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n714), .A2(new_n573), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n418), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n713), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(new_n382), .ZN(G24));
  INV_X1    g536(.A(new_n718), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n723), .B(new_n637), .C1(new_n608), .C2(new_n607), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n589), .A2(new_n681), .A3(new_n708), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G125), .ZN(G27));
  INV_X1    g541(.A(KEYINPUT42), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT104), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n470), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n467), .A2(new_n469), .A3(KEYINPUT104), .A4(G469), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n730), .A2(new_n464), .A3(new_n472), .A4(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n474), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n581), .B1(new_n294), .B2(new_n296), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n734), .A2(new_n735), .A3(new_n602), .A4(new_n651), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n728), .B1(new_n736), .B2(new_n575), .ZN(new_n737));
  INV_X1    g551(.A(new_n528), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT105), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n527), .B1(new_n603), .B2(new_n606), .ZN(new_n740));
  AOI211_X1 g554(.A(new_n739), .B(KEYINPUT106), .C1(new_n740), .C2(KEYINPUT32), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT106), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n742), .B1(new_n534), .B2(KEYINPUT105), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n738), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  AOI211_X1 g558(.A(new_n517), .B(new_n527), .C1(new_n603), .C2(new_n606), .ZN(new_n745));
  OAI21_X1  g559(.A(KEYINPUT106), .B1(new_n745), .B2(new_n739), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n534), .A2(KEYINPUT105), .A3(new_n742), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(new_n528), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n744), .A2(new_n516), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n574), .ZN(new_n750));
  AOI211_X1 g564(.A(new_n581), .B(new_n650), .C1(new_n294), .C2(new_n296), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n751), .A2(KEYINPUT42), .A3(new_n602), .A4(new_n734), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n737), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G131), .ZN(G33));
  NOR2_X1   g568(.A1(new_n575), .A2(new_n733), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n735), .A2(new_n626), .A3(new_n651), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G134), .ZN(G36));
  NAND3_X1  g572(.A1(new_n679), .A2(new_n371), .A3(new_n372), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT43), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT43), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n679), .A2(new_n371), .A3(new_n761), .A4(new_n372), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n609), .A3(new_n637), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(KEYINPUT44), .ZN(new_n765));
  INV_X1    g579(.A(new_n474), .ZN(new_n766));
  INV_X1    g580(.A(new_n464), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT45), .B1(new_n467), .B2(new_n469), .ZN(new_n768));
  OAI21_X1  g582(.A(KEYINPUT107), .B1(new_n768), .B2(new_n422), .ZN(new_n769));
  AOI22_X1  g583(.A1(new_n465), .A2(new_n466), .B1(new_n468), .B2(new_n462), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT45), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT107), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n772), .B(G469), .C1(new_n770), .C2(KEYINPUT45), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n769), .A2(new_n771), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n472), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT46), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n767), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n774), .A2(KEYINPUT46), .A3(new_n472), .ZN(new_n778));
  AOI211_X1 g592(.A(new_n766), .B(new_n656), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n735), .B(KEYINPUT108), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n765), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G137), .ZN(G39));
  AOI21_X1  g597(.A(new_n766), .B1(new_n777), .B2(new_n778), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT109), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(KEYINPUT47), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n785), .A2(KEYINPUT47), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n786), .B1(new_n784), .B2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n751), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n679), .B1(new_n702), .B2(new_n703), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n535), .A2(new_n574), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n787), .A2(new_n789), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G140), .ZN(G42));
  NAND4_X1  g609(.A1(new_n760), .A2(new_n648), .A3(new_n719), .A4(new_n762), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT50), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n295), .B1(KEYINPUT113), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n663), .A2(new_n664), .A3(new_n798), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n796), .A2(new_n799), .A3(new_n688), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n797), .A2(KEYINPUT113), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NOR4_X1   g617(.A1(new_n796), .A2(new_n799), .A3(new_n688), .A4(new_n801), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT51), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n687), .A2(new_n464), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n807), .A2(new_n474), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n808), .B1(new_n787), .B2(new_n789), .ZN(new_n809));
  INV_X1    g623(.A(new_n796), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n781), .A2(new_n810), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n805), .B(new_n806), .C1(new_n809), .C2(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n812), .B1(KEYINPUT115), .B2(new_n806), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n763), .A2(new_n648), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n735), .A2(new_n708), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT114), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n814), .A2(new_n725), .A3(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n673), .A2(new_n573), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n678), .A2(new_n679), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n816), .A2(new_n412), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n813), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n805), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n809), .B(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n811), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n825), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n823), .B1(new_n829), .B2(new_n806), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n576), .A2(new_n476), .B1(new_n639), .B2(new_n640), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n407), .A2(new_n368), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n832), .B1(new_n621), .B2(new_n625), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n535), .A2(new_n645), .A3(new_n637), .A4(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n791), .A2(new_n733), .A3(new_n724), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n751), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n791), .B1(new_n678), .B2(new_n407), .ZN(new_n838));
  INV_X1    g652(.A(new_n297), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n838), .A2(new_n839), .A3(new_n418), .A4(new_n610), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n831), .A2(new_n837), .A3(new_n757), .A4(new_n840), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n589), .B(new_n646), .C1(new_n652), .C2(new_n681), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n673), .A2(new_n638), .A3(new_n651), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n589), .A2(new_n666), .A3(new_n843), .A4(new_n734), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n842), .A2(new_n726), .A3(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n842), .A2(new_n726), .A3(new_n844), .A4(KEYINPUT52), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n841), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n721), .A2(new_n694), .ZN(new_n850));
  AND4_X1   g664(.A1(new_n698), .A2(new_n753), .A3(new_n711), .A4(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT53), .B1(new_n849), .B2(new_n851), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT54), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n847), .A2(new_n848), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n853), .B1(new_n841), .B2(KEYINPUT111), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n831), .A2(new_n840), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n837), .A2(new_n757), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT111), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  AND4_X1   g676(.A1(new_n851), .A2(new_n857), .A3(new_n858), .A4(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n863), .A2(new_n855), .ZN(new_n864));
  XOR2_X1   g678(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n810), .A2(new_n700), .ZN(new_n868));
  AND4_X1   g682(.A1(new_n412), .A2(new_n816), .A3(new_n602), .A4(new_n818), .ZN(new_n869));
  INV_X1    g683(.A(new_n750), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n870), .A2(new_n814), .A3(new_n816), .ZN(new_n871));
  OR2_X1    g685(.A1(new_n871), .A2(KEYINPUT48), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(KEYINPUT48), .ZN(new_n873));
  AOI211_X1 g687(.A(new_n868), .B(new_n869), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n830), .A2(new_n856), .A3(new_n867), .A4(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n409), .B1(new_n875), .B2(KEYINPUT117), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT117), .ZN(new_n877));
  OAI21_X1  g691(.A(G953), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  NOR4_X1   g692(.A1(new_n759), .A2(new_n573), .A3(new_n766), .A4(new_n581), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT110), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n807), .A2(KEYINPUT49), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n665), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n673), .B1(KEYINPUT49), .B2(new_n807), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n880), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n876), .A2(new_n878), .A3(new_n884), .ZN(G75));
  OAI211_X1 g699(.A(G210), .B(G902), .C1(new_n863), .C2(new_n855), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT56), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n283), .A2(new_n286), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(new_n285), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT55), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n891), .B1(KEYINPUT118), .B2(new_n887), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n888), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n408), .A2(G953), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT119), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n886), .B(new_n887), .C1(KEYINPUT118), .C2(new_n891), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n893), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT120), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT120), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n893), .A2(new_n899), .A3(new_n896), .A4(new_n895), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n898), .A2(new_n900), .ZN(G51));
  INV_X1    g715(.A(new_n895), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n852), .A2(new_n853), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n851), .A2(new_n858), .A3(new_n857), .A4(new_n862), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n865), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n867), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n471), .B(KEYINPUT57), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n909), .B1(new_n463), .B2(new_n460), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n365), .B1(new_n903), .B2(new_n904), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n911), .A2(new_n771), .A3(new_n769), .A4(new_n773), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n902), .B1(new_n910), .B2(new_n912), .ZN(G54));
  NAND2_X1  g727(.A1(new_n356), .A2(new_n358), .ZN(new_n914));
  OAI211_X1 g728(.A(KEYINPUT58), .B(G902), .C1(new_n863), .C2(new_n855), .ZN(new_n915));
  INV_X1    g729(.A(G475), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n914), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n911), .A2(KEYINPUT58), .A3(G475), .A4(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n895), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT121), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n920), .A2(KEYINPUT121), .A3(new_n895), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(G60));
  NAND2_X1  g739(.A1(G478), .A2(G902), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT59), .Z(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n907), .A2(new_n599), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n867), .A2(new_n856), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n599), .B1(new_n930), .B2(new_n928), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n929), .A2(new_n931), .A3(new_n902), .ZN(G63));
  NAND2_X1  g746(.A1(G217), .A2(G902), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT60), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n905), .A2(new_n635), .A3(new_n935), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n936), .A2(new_n895), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n559), .B1(new_n905), .B2(new_n935), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT122), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n937), .A2(new_n939), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n940), .A2(new_n941), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n936), .A2(new_n895), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n943), .B(new_n944), .C1(new_n945), .C2(new_n938), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n942), .A2(new_n946), .ZN(G66));
  AOI21_X1  g761(.A(new_n265), .B1(new_n266), .B2(new_n413), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n859), .A2(new_n698), .A3(new_n711), .A4(new_n850), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n948), .B1(new_n949), .B2(new_n265), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n889), .B1(G898), .B2(new_n265), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n950), .B(new_n951), .Z(G69));
  NAND2_X1  g766(.A1(new_n315), .A2(new_n316), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n522), .B(new_n953), .Z(new_n954));
  AOI21_X1  g768(.A(new_n265), .B1(G227), .B2(G900), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT123), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT62), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n842), .A2(new_n726), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n676), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n956), .A2(new_n957), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n782), .A2(new_n794), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n676), .A2(new_n956), .A3(new_n957), .A4(new_n959), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n575), .A2(new_n657), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n965), .A2(new_n735), .A3(new_n838), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n962), .A2(new_n963), .A3(new_n964), .A4(new_n966), .ZN(new_n967));
  AOI211_X1 g781(.A(new_n954), .B(new_n955), .C1(new_n967), .C2(new_n265), .ZN(new_n968));
  OAI21_X1  g782(.A(G953), .B1(new_n649), .B2(G227), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n870), .A2(new_n779), .A3(new_n589), .A4(new_n666), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n959), .A2(new_n753), .A3(new_n757), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n963), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n969), .B(new_n954), .C1(new_n972), .C2(G953), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(KEYINPUT124), .B1(new_n968), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n954), .B1(new_n967), .B2(new_n265), .ZN(new_n976));
  INV_X1    g790(.A(new_n955), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT124), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n978), .A2(new_n979), .A3(new_n973), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n975), .A2(new_n980), .ZN(G72));
  XNOR2_X1  g795(.A(new_n852), .B(new_n853), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n669), .B(KEYINPUT63), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n488), .A2(new_n493), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n518), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n982), .A2(new_n984), .A3(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT127), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n982), .A2(KEYINPUT127), .A3(new_n984), .A4(new_n986), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n984), .B1(new_n967), .B2(new_n949), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n523), .B(KEYINPUT125), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n992), .A2(new_n513), .A3(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n984), .B1(new_n972), .B2(new_n949), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n993), .A2(new_n513), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n996), .B(KEYINPUT126), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n902), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  AND3_X1   g812(.A1(new_n991), .A2(new_n994), .A3(new_n998), .ZN(G57));
endmodule


