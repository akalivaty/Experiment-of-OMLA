

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787;

  BUF_X1 U372 ( .A(G143), .Z(n350) );
  XNOR2_X1 U373 ( .A(n492), .B(n425), .ZN(n771) );
  INV_X1 U374 ( .A(G143), .ZN(n451) );
  AND2_X2 U375 ( .A1(n392), .A2(n445), .ZN(n391) );
  XNOR2_X2 U376 ( .A(n504), .B(n452), .ZN(n534) );
  NOR2_X1 U377 ( .A1(n708), .A2(n711), .ZN(n547) );
  XNOR2_X2 U378 ( .A(KEYINPUT4), .B(KEYINPUT91), .ZN(n428) );
  NOR2_X2 U379 ( .A1(n703), .A2(n649), .ZN(n752) );
  XNOR2_X2 U380 ( .A(n419), .B(n359), .ZN(n588) );
  INV_X2 U381 ( .A(n588), .ZN(n388) );
  XOR2_X2 U382 ( .A(n541), .B(G478), .Z(n568) );
  NAND2_X1 U383 ( .A1(n648), .A2(n647), .ZN(n703) );
  XNOR2_X1 U384 ( .A(n432), .B(n360), .ZN(n621) );
  OR2_X1 U385 ( .A1(n553), .A2(n554), .ZN(n691) );
  AND2_X1 U386 ( .A1(n405), .A2(n404), .ZN(n403) );
  NOR2_X1 U387 ( .A1(G237), .A2(G902), .ZN(n466) );
  INV_X1 U388 ( .A(G134), .ZN(n452) );
  XNOR2_X1 U389 ( .A(n365), .B(G137), .ZN(n491) );
  INV_X1 U390 ( .A(KEYINPUT67), .ZN(n365) );
  XNOR2_X1 U391 ( .A(n534), .B(n453), .ZN(n492) );
  XNOR2_X1 U392 ( .A(G131), .B(KEYINPUT4), .ZN(n453) );
  XNOR2_X1 U393 ( .A(n468), .B(n361), .ZN(n418) );
  OR2_X1 U394 ( .A1(n659), .A2(n401), .ZN(n400) );
  NAND2_X1 U395 ( .A1(n402), .A2(n512), .ZN(n401) );
  NAND2_X1 U396 ( .A1(n517), .A2(n638), .ZN(n404) );
  XNOR2_X1 U397 ( .A(n529), .B(n448), .ZN(n567) );
  XNOR2_X1 U398 ( .A(KEYINPUT3), .B(G119), .ZN(n457) );
  XNOR2_X1 U399 ( .A(G101), .B(KEYINPUT68), .ZN(n455) );
  AND2_X1 U400 ( .A1(n372), .A2(n352), .ZN(n371) );
  NAND2_X1 U401 ( .A1(n556), .A2(KEYINPUT47), .ZN(n372) );
  INV_X1 U402 ( .A(n657), .ZN(n374) );
  XNOR2_X1 U403 ( .A(n376), .B(n375), .ZN(n373) );
  OR2_X1 U404 ( .A1(n514), .A2(n467), .ZN(n705) );
  AND2_X1 U405 ( .A1(n418), .A2(n413), .ZN(n412) );
  NAND2_X1 U406 ( .A1(n385), .A2(n383), .ZN(n382) );
  NAND2_X1 U407 ( .A1(n384), .A2(KEYINPUT19), .ZN(n383) );
  NAND2_X1 U408 ( .A1(n387), .A2(n386), .ZN(n385) );
  INV_X1 U409 ( .A(n705), .ZN(n384) );
  NOR2_X1 U410 ( .A1(n403), .A2(n381), .ZN(n380) );
  INV_X1 U411 ( .A(n386), .ZN(n381) );
  INV_X1 U412 ( .A(KEYINPUT66), .ZN(n406) );
  NOR2_X1 U413 ( .A1(G902), .A2(n745), .ZN(n493) );
  INV_X1 U414 ( .A(G902), .ZN(n462) );
  XNOR2_X1 U415 ( .A(n395), .B(n461), .ZN(n650) );
  NAND2_X1 U416 ( .A1(n397), .A2(n438), .ZN(n395) );
  XNOR2_X1 U417 ( .A(n526), .B(n449), .ZN(n527) );
  XNOR2_X1 U418 ( .A(n424), .B(G140), .ZN(n423) );
  INV_X1 U419 ( .A(KEYINPUT97), .ZN(n424) );
  XNOR2_X1 U420 ( .A(n430), .B(G146), .ZN(n505) );
  INV_X1 U421 ( .A(G125), .ZN(n430) );
  XOR2_X1 U422 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n503) );
  AND2_X1 U423 ( .A1(n373), .A2(n374), .ZN(n773) );
  XNOR2_X1 U424 ( .A(n519), .B(n518), .ZN(n632) );
  XNOR2_X1 U425 ( .A(KEYINPUT71), .B(KEYINPUT39), .ZN(n518) );
  XNOR2_X1 U426 ( .A(n587), .B(n586), .ZN(n594) );
  INV_X1 U427 ( .A(n719), .ZN(n615) );
  INV_X1 U428 ( .A(G107), .ZN(n488) );
  XNOR2_X1 U429 ( .A(KEYINPUT16), .B(G122), .ZN(n508) );
  NAND2_X1 U430 ( .A1(n368), .A2(n716), .ZN(n370) );
  XNOR2_X1 U431 ( .A(n562), .B(n362), .ZN(n368) );
  XNOR2_X1 U432 ( .A(KEYINPUT15), .B(G902), .ZN(n512) );
  NOR2_X1 U433 ( .A1(n566), .A2(n369), .ZN(n572) );
  NAND2_X1 U434 ( .A1(n371), .A2(n370), .ZN(n369) );
  AND2_X1 U435 ( .A1(n705), .A2(n551), .ZN(n386) );
  XNOR2_X1 U436 ( .A(n516), .B(n515), .ZN(n517) );
  NOR2_X1 U437 ( .A1(G953), .A2(G237), .ZN(n459) );
  OR2_X1 U438 ( .A1(n492), .A2(n358), .ZN(n397) );
  NAND2_X1 U439 ( .A1(n492), .A2(n439), .ZN(n438) );
  NAND2_X1 U440 ( .A1(n441), .A2(n440), .ZN(n439) );
  NAND2_X1 U441 ( .A1(n454), .A2(G146), .ZN(n441) );
  NAND2_X1 U442 ( .A1(n442), .A2(n443), .ZN(n440) );
  XNOR2_X1 U443 ( .A(G116), .B(G113), .ZN(n456) );
  XNOR2_X1 U444 ( .A(G113), .B(G131), .ZN(n524) );
  XOR2_X1 U445 ( .A(G104), .B(G122), .Z(n525) );
  INV_X1 U446 ( .A(KEYINPUT89), .ZN(n434) );
  NAND2_X1 U447 ( .A1(G234), .A2(G237), .ZN(n497) );
  XOR2_X1 U448 ( .A(KEYINPUT38), .B(n550), .Z(n706) );
  OR2_X1 U449 ( .A1(n602), .A2(KEYINPUT34), .ZN(n389) );
  XNOR2_X1 U450 ( .A(n364), .B(n356), .ZN(n543) );
  OR2_X1 U451 ( .A1(n755), .A2(G902), .ZN(n364) );
  XOR2_X1 U452 ( .A(KEYINPUT24), .B(G110), .Z(n474) );
  XNOR2_X1 U453 ( .A(G119), .B(G128), .ZN(n473) );
  XNOR2_X1 U454 ( .A(n491), .B(KEYINPUT99), .ZN(n477) );
  XNOR2_X1 U455 ( .A(n505), .B(n444), .ZN(n770) );
  XNOR2_X1 U456 ( .A(G140), .B(KEYINPUT10), .ZN(n444) );
  XNOR2_X1 U457 ( .A(KEYINPUT85), .B(KEYINPUT8), .ZN(n471) );
  XNOR2_X1 U458 ( .A(G116), .B(G122), .ZN(n531) );
  XOR2_X1 U459 ( .A(KEYINPUT106), .B(G107), .Z(n532) );
  INV_X1 U460 ( .A(G953), .ZN(n502) );
  NOR2_X1 U461 ( .A1(n561), .A2(n691), .ZN(n575) );
  AND2_X1 U462 ( .A1(n418), .A2(n415), .ZN(n409) );
  NAND2_X1 U463 ( .A1(n403), .A2(n400), .ZN(n550) );
  NOR2_X1 U464 ( .A1(n382), .A2(n380), .ZN(n379) );
  AND2_X1 U465 ( .A1(n366), .A2(n353), .ZN(n552) );
  XNOR2_X1 U466 ( .A(n367), .B(KEYINPUT28), .ZN(n366) );
  NOR2_X1 U467 ( .A1(n559), .A2(n615), .ZN(n367) );
  INV_X1 U468 ( .A(KEYINPUT105), .ZN(n530) );
  XNOR2_X1 U469 ( .A(n496), .B(n495), .ZN(n601) );
  INV_X1 U470 ( .A(KEYINPUT101), .ZN(n495) );
  XNOR2_X1 U471 ( .A(n594), .B(KEYINPUT96), .ZN(n602) );
  XNOR2_X1 U472 ( .A(n463), .B(KEYINPUT102), .ZN(n464) );
  AND2_X1 U473 ( .A1(n650), .A2(n462), .ZN(n465) );
  NAND2_X1 U474 ( .A1(n621), .A2(n596), .ZN(n617) );
  XNOR2_X1 U475 ( .A(n719), .B(n396), .ZN(n597) );
  INV_X1 U476 ( .A(KEYINPUT6), .ZN(n396) );
  XOR2_X1 U477 ( .A(KEYINPUT62), .B(n650), .Z(n651) );
  XNOR2_X1 U478 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U479 ( .A(n771), .B(n421), .ZN(n745) );
  XNOR2_X1 U480 ( .A(n490), .B(n422), .ZN(n421) );
  XNOR2_X1 U481 ( .A(n487), .B(n423), .ZN(n422) );
  XNOR2_X1 U482 ( .A(n511), .B(n765), .ZN(n659) );
  AND2_X1 U483 ( .A1(n653), .A2(G953), .ZN(n757) );
  NAND2_X1 U484 ( .A1(n643), .A2(n642), .ZN(n648) );
  AND2_X1 U485 ( .A1(n773), .A2(n354), .ZN(n646) );
  BUF_X1 U486 ( .A(n611), .Z(n673) );
  INV_X1 U487 ( .A(n370), .ZN(n697) );
  AND2_X1 U488 ( .A1(n373), .A2(n357), .ZN(n351) );
  OR2_X1 U489 ( .A1(n687), .A2(KEYINPUT84), .ZN(n352) );
  XOR2_X1 U490 ( .A(n558), .B(KEYINPUT110), .Z(n353) );
  BUF_X1 U491 ( .A(n580), .Z(n716) );
  AND2_X1 U492 ( .A1(n645), .A2(KEYINPUT81), .ZN(n354) );
  OR2_X1 U493 ( .A1(n584), .A2(n583), .ZN(n355) );
  XOR2_X1 U494 ( .A(n484), .B(KEYINPUT25), .Z(n356) );
  AND2_X1 U495 ( .A1(n374), .A2(n772), .ZN(n357) );
  AND2_X1 U496 ( .A1(n437), .A2(n436), .ZN(n358) );
  INV_X1 U497 ( .A(G146), .ZN(n443) );
  XOR2_X1 U498 ( .A(n581), .B(KEYINPUT33), .Z(n359) );
  XOR2_X1 U499 ( .A(KEYINPUT64), .B(KEYINPUT22), .Z(n360) );
  XNOR2_X1 U500 ( .A(KEYINPUT109), .B(KEYINPUT30), .ZN(n361) );
  XOR2_X1 U501 ( .A(KEYINPUT90), .B(KEYINPUT36), .Z(n362) );
  INV_X1 U502 ( .A(KEYINPUT76), .ZN(n417) );
  INV_X1 U503 ( .A(KEYINPUT34), .ZN(n589) );
  XNOR2_X1 U504 ( .A(n363), .B(n479), .ZN(n755) );
  XNOR2_X1 U505 ( .A(n478), .B(n480), .ZN(n363) );
  NAND2_X1 U506 ( .A1(n545), .A2(n720), .ZN(n559) );
  INV_X1 U507 ( .A(KEYINPUT48), .ZN(n375) );
  NAND2_X1 U508 ( .A1(n574), .A2(n573), .ZN(n376) );
  NAND2_X1 U509 ( .A1(n379), .A2(n377), .ZN(n585) );
  NAND2_X1 U510 ( .A1(n378), .A2(n403), .ZN(n377) );
  AND2_X1 U511 ( .A1(n400), .A2(KEYINPUT19), .ZN(n378) );
  INV_X1 U512 ( .A(n400), .ZN(n387) );
  NAND2_X1 U513 ( .A1(n585), .A2(n355), .ZN(n587) );
  NAND2_X1 U514 ( .A1(n388), .A2(KEYINPUT34), .ZN(n392) );
  NAND2_X1 U515 ( .A1(n390), .A2(n389), .ZN(n393) );
  NAND2_X1 U516 ( .A1(n394), .A2(n602), .ZN(n390) );
  NAND2_X1 U517 ( .A1(n393), .A2(n391), .ZN(n593) );
  NAND2_X1 U518 ( .A1(n588), .A2(n589), .ZN(n394) );
  INV_X1 U519 ( .A(n729), .ZN(n736) );
  XNOR2_X1 U520 ( .A(n547), .B(n546), .ZN(n729) );
  XNOR2_X2 U521 ( .A(n465), .B(n464), .ZN(n719) );
  NAND2_X1 U522 ( .A1(n408), .A2(n410), .ZN(n570) );
  NAND2_X1 U523 ( .A1(n575), .A2(n550), .ZN(n562) );
  NAND2_X1 U524 ( .A1(n409), .A2(n414), .ZN(n408) );
  NAND2_X2 U525 ( .A1(n758), .A2(n351), .ZN(n701) );
  XNOR2_X1 U526 ( .A(n398), .B(n610), .ZN(n630) );
  NAND2_X1 U527 ( .A1(n399), .A2(n450), .ZN(n398) );
  XNOR2_X1 U528 ( .A(n435), .B(n434), .ZN(n399) );
  NAND2_X1 U529 ( .A1(n752), .A2(G475), .ZN(n669) );
  INV_X1 U530 ( .A(n517), .ZN(n402) );
  NAND2_X1 U531 ( .A1(n659), .A2(n517), .ZN(n405) );
  NAND2_X1 U532 ( .A1(n715), .A2(n494), .ZN(n496) );
  XNOR2_X2 U533 ( .A(n407), .B(n406), .ZN(n715) );
  NAND2_X1 U534 ( .A1(n543), .A2(n720), .ZN(n407) );
  NAND2_X1 U535 ( .A1(n411), .A2(n412), .ZN(n410) );
  NAND2_X1 U536 ( .A1(n414), .A2(n416), .ZN(n411) );
  NAND2_X1 U537 ( .A1(n416), .A2(KEYINPUT76), .ZN(n413) );
  INV_X1 U538 ( .A(n601), .ZN(n414) );
  NOR2_X1 U539 ( .A1(n544), .A2(n417), .ZN(n415) );
  NAND2_X1 U540 ( .A1(n544), .A2(n417), .ZN(n416) );
  NAND2_X1 U541 ( .A1(n570), .A2(n706), .ZN(n519) );
  NAND2_X1 U542 ( .A1(n420), .A2(n597), .ZN(n419) );
  INV_X1 U543 ( .A(n604), .ZN(n420) );
  INV_X1 U544 ( .A(n491), .ZN(n425) );
  XNOR2_X1 U545 ( .A(n426), .B(n503), .ZN(n431) );
  XNOR2_X1 U546 ( .A(n428), .B(n427), .ZN(n426) );
  NAND2_X1 U547 ( .A1(n502), .A2(G224), .ZN(n427) );
  XNOR2_X1 U548 ( .A(n431), .B(n429), .ZN(n507) );
  XNOR2_X1 U549 ( .A(n504), .B(n505), .ZN(n429) );
  NAND2_X1 U550 ( .A1(n594), .A2(n433), .ZN(n432) );
  AND2_X1 U551 ( .A1(n595), .A2(n720), .ZN(n433) );
  XNOR2_X1 U552 ( .A(n593), .B(n446), .ZN(n611) );
  XNOR2_X1 U553 ( .A(n477), .B(n476), .ZN(n478) );
  NAND2_X1 U554 ( .A1(n611), .A2(KEYINPUT44), .ZN(n435) );
  INV_X1 U555 ( .A(n454), .ZN(n442) );
  NAND2_X1 U556 ( .A1(n454), .A2(n443), .ZN(n436) );
  NAND2_X1 U557 ( .A1(n442), .A2(G146), .ZN(n437) );
  XNOR2_X2 U558 ( .A(n631), .B(KEYINPUT45), .ZN(n758) );
  XOR2_X1 U559 ( .A(n591), .B(KEYINPUT78), .Z(n445) );
  XOR2_X1 U560 ( .A(n592), .B(KEYINPUT35), .Z(n446) );
  AND2_X1 U561 ( .A1(n609), .A2(n608), .ZN(n447) );
  XOR2_X1 U562 ( .A(KEYINPUT13), .B(G475), .Z(n448) );
  XOR2_X1 U563 ( .A(n525), .B(n524), .Z(n449) );
  NOR2_X1 U564 ( .A1(n674), .A2(n447), .ZN(n450) );
  XNOR2_X1 U565 ( .A(n510), .B(n460), .ZN(n461) );
  XNOR2_X1 U566 ( .A(n558), .B(n557), .ZN(n580) );
  XNOR2_X1 U567 ( .A(n528), .B(n527), .ZN(n667) );
  XNOR2_X1 U568 ( .A(n567), .B(n530), .ZN(n553) );
  AND2_X1 U569 ( .A1(n600), .A2(n721), .ZN(n674) );
  XNOR2_X2 U570 ( .A(n451), .B(G128), .ZN(n504) );
  XOR2_X1 U571 ( .A(G137), .B(KEYINPUT5), .Z(n454) );
  XNOR2_X1 U572 ( .A(n456), .B(n455), .ZN(n458) );
  XNOR2_X1 U573 ( .A(n458), .B(n457), .ZN(n510) );
  XOR2_X1 U574 ( .A(KEYINPUT75), .B(n459), .Z(n523) );
  NAND2_X1 U575 ( .A1(n523), .A2(G210), .ZN(n460) );
  INV_X1 U576 ( .A(G472), .ZN(n463) );
  XNOR2_X1 U577 ( .A(n466), .B(KEYINPUT74), .ZN(n514) );
  INV_X1 U578 ( .A(G214), .ZN(n467) );
  NAND2_X1 U579 ( .A1(n719), .A2(n705), .ZN(n468) );
  NAND2_X1 U580 ( .A1(n512), .A2(G234), .ZN(n469) );
  XNOR2_X1 U581 ( .A(n469), .B(KEYINPUT20), .ZN(n481) );
  NAND2_X1 U582 ( .A1(G221), .A2(n481), .ZN(n470) );
  XOR2_X1 U583 ( .A(KEYINPUT21), .B(n470), .Z(n720) );
  BUF_X2 U584 ( .A(n502), .Z(n775) );
  NAND2_X1 U585 ( .A1(n775), .A2(G234), .ZN(n472) );
  XNOR2_X1 U586 ( .A(n472), .B(n471), .ZN(n535) );
  NAND2_X1 U587 ( .A1(n535), .A2(G221), .ZN(n480) );
  XNOR2_X1 U588 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U589 ( .A(n770), .B(n475), .ZN(n479) );
  XOR2_X1 U590 ( .A(KEYINPUT23), .B(KEYINPUT98), .Z(n476) );
  XOR2_X1 U591 ( .A(KEYINPUT100), .B(KEYINPUT77), .Z(n483) );
  NAND2_X1 U592 ( .A1(n481), .A2(G217), .ZN(n482) );
  XNOR2_X1 U593 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U594 ( .A(G101), .B(G146), .Z(n486) );
  NAND2_X1 U595 ( .A1(G227), .A2(n775), .ZN(n485) );
  XNOR2_X1 U596 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U597 ( .A(G104), .B(G110), .ZN(n489) );
  XNOR2_X1 U598 ( .A(n489), .B(n488), .ZN(n764) );
  XNOR2_X1 U599 ( .A(n764), .B(KEYINPUT69), .ZN(n506) );
  INV_X1 U600 ( .A(n506), .ZN(n490) );
  XNOR2_X2 U601 ( .A(n493), .B(G469), .ZN(n558) );
  INV_X1 U602 ( .A(n558), .ZN(n494) );
  XOR2_X1 U603 ( .A(KEYINPUT73), .B(KEYINPUT14), .Z(n498) );
  XNOR2_X1 U604 ( .A(n498), .B(n497), .ZN(n499) );
  NAND2_X1 U605 ( .A1(G952), .A2(n499), .ZN(n735) );
  NOR2_X1 U606 ( .A1(n735), .A2(G953), .ZN(n584) );
  NAND2_X1 U607 ( .A1(G902), .A2(n499), .ZN(n582) );
  OR2_X1 U608 ( .A1(n775), .A2(n582), .ZN(n500) );
  NOR2_X1 U609 ( .A1(G900), .A2(n500), .ZN(n501) );
  NOR2_X1 U610 ( .A1(n584), .A2(n501), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n507), .B(n506), .ZN(n511) );
  XNOR2_X1 U612 ( .A(n508), .B(KEYINPUT72), .ZN(n509) );
  XNOR2_X1 U613 ( .A(n510), .B(n509), .ZN(n765) );
  INV_X1 U614 ( .A(n512), .ZN(n638) );
  INV_X1 U615 ( .A(G210), .ZN(n513) );
  OR2_X1 U616 ( .A1(n514), .A2(n513), .ZN(n516) );
  XNOR2_X1 U617 ( .A(KEYINPUT94), .B(KEYINPUT95), .ZN(n515) );
  XOR2_X1 U618 ( .A(KEYINPUT12), .B(KEYINPUT104), .Z(n521) );
  XNOR2_X1 U619 ( .A(n350), .B(KEYINPUT11), .ZN(n520) );
  XNOR2_X1 U620 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U621 ( .A(n770), .B(n522), .Z(n528) );
  NAND2_X1 U622 ( .A1(G214), .A2(n523), .ZN(n526) );
  NOR2_X1 U623 ( .A1(G902), .A2(n667), .ZN(n529) );
  XNOR2_X1 U624 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n539) );
  XNOR2_X1 U625 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U626 ( .A(n534), .B(n533), .Z(n537) );
  NAND2_X1 U627 ( .A1(G217), .A2(n535), .ZN(n536) );
  XNOR2_X1 U628 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U629 ( .A(n539), .B(n538), .ZN(n749) );
  NOR2_X1 U630 ( .A1(G902), .A2(n749), .ZN(n540) );
  XNOR2_X1 U631 ( .A(n540), .B(KEYINPUT107), .ZN(n541) );
  INV_X1 U632 ( .A(n568), .ZN(n554) );
  NOR2_X1 U633 ( .A1(n632), .A2(n691), .ZN(n542) );
  XNOR2_X1 U634 ( .A(n542), .B(KEYINPUT40), .ZN(n786) );
  BUF_X1 U635 ( .A(n543), .Z(n721) );
  NOR2_X1 U636 ( .A1(n544), .A2(n721), .ZN(n545) );
  NAND2_X1 U637 ( .A1(n568), .A2(n567), .ZN(n708) );
  NAND2_X1 U638 ( .A1(n706), .A2(n705), .ZN(n711) );
  XNOR2_X1 U639 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n546) );
  NAND2_X1 U640 ( .A1(n552), .A2(n729), .ZN(n548) );
  XOR2_X1 U641 ( .A(KEYINPUT42), .B(n548), .Z(n784) );
  NOR2_X1 U642 ( .A1(n786), .A2(n784), .ZN(n549) );
  XNOR2_X1 U643 ( .A(n549), .B(KEYINPUT46), .ZN(n574) );
  INV_X1 U644 ( .A(KEYINPUT19), .ZN(n551) );
  NAND2_X1 U645 ( .A1(n552), .A2(n585), .ZN(n687) );
  NAND2_X1 U646 ( .A1(n687), .A2(KEYINPUT84), .ZN(n555) );
  NAND2_X1 U647 ( .A1(n554), .A2(n553), .ZN(n694) );
  NAND2_X1 U648 ( .A1(n691), .A2(n694), .ZN(n608) );
  NAND2_X1 U649 ( .A1(n555), .A2(n608), .ZN(n556) );
  INV_X1 U650 ( .A(KEYINPUT1), .ZN(n557) );
  INV_X1 U651 ( .A(n716), .ZN(n596) );
  INV_X1 U652 ( .A(n597), .ZN(n618) );
  NOR2_X1 U653 ( .A1(n618), .A2(n559), .ZN(n560) );
  NAND2_X1 U654 ( .A1(n560), .A2(n705), .ZN(n561) );
  INV_X1 U655 ( .A(KEYINPUT84), .ZN(n564) );
  INV_X1 U656 ( .A(n608), .ZN(n710) );
  NOR2_X1 U657 ( .A1(n687), .A2(n710), .ZN(n563) );
  NOR2_X1 U658 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U659 ( .A1(KEYINPUT47), .A2(n565), .ZN(n566) );
  NOR2_X1 U660 ( .A1(n568), .A2(n567), .ZN(n590) );
  AND2_X1 U661 ( .A1(n550), .A2(n590), .ZN(n569) );
  AND2_X1 U662 ( .A1(n570), .A2(n569), .ZN(n686) );
  INV_X1 U663 ( .A(n686), .ZN(n571) );
  AND2_X1 U664 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U665 ( .A(n575), .B(KEYINPUT108), .ZN(n576) );
  NAND2_X1 U666 ( .A1(n576), .A2(n596), .ZN(n577) );
  XNOR2_X1 U667 ( .A(KEYINPUT43), .B(n577), .ZN(n579) );
  INV_X1 U668 ( .A(n550), .ZN(n578) );
  AND2_X1 U669 ( .A1(n579), .A2(n578), .ZN(n657) );
  NAND2_X1 U670 ( .A1(n580), .A2(n715), .ZN(n604) );
  INV_X1 U671 ( .A(KEYINPUT70), .ZN(n581) );
  OR2_X1 U672 ( .A1(n775), .A2(G898), .ZN(n766) );
  NOR2_X1 U673 ( .A1(n582), .A2(n766), .ZN(n583) );
  INV_X1 U674 ( .A(KEYINPUT0), .ZN(n586) );
  INV_X1 U675 ( .A(n590), .ZN(n591) );
  INV_X1 U676 ( .A(KEYINPUT86), .ZN(n592) );
  INV_X1 U677 ( .A(n708), .ZN(n595) );
  NOR2_X2 U678 ( .A1(n617), .A2(n597), .ZN(n599) );
  INV_X1 U679 ( .A(KEYINPUT87), .ZN(n598) );
  XNOR2_X1 U680 ( .A(n599), .B(n598), .ZN(n600) );
  NOR2_X1 U681 ( .A1(n601), .A2(n719), .ZN(n603) );
  NAND2_X1 U682 ( .A1(n603), .A2(n602), .ZN(n678) );
  OR2_X1 U683 ( .A1(n604), .A2(n615), .ZN(n726) );
  INV_X1 U684 ( .A(n726), .ZN(n605) );
  NAND2_X1 U685 ( .A1(n594), .A2(n605), .ZN(n607) );
  XNOR2_X1 U686 ( .A(KEYINPUT31), .B(KEYINPUT103), .ZN(n606) );
  XNOR2_X1 U687 ( .A(n607), .B(n606), .ZN(n693) );
  NAND2_X1 U688 ( .A1(n678), .A2(n693), .ZN(n609) );
  INV_X1 U689 ( .A(KEYINPUT88), .ZN(n610) );
  INV_X1 U690 ( .A(n673), .ZN(n613) );
  INV_X1 U691 ( .A(KEYINPUT44), .ZN(n612) );
  NAND2_X1 U692 ( .A1(n613), .A2(n612), .ZN(n625) );
  INV_X1 U693 ( .A(n721), .ZN(n614) );
  NAND2_X1 U694 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U695 ( .A1(n617), .A2(n616), .ZN(n681) );
  XNOR2_X1 U696 ( .A(KEYINPUT32), .B(KEYINPUT79), .ZN(n624) );
  NAND2_X1 U697 ( .A1(n618), .A2(n716), .ZN(n619) );
  NOR2_X1 U698 ( .A1(n721), .A2(n619), .ZN(n620) );
  XNOR2_X1 U699 ( .A(KEYINPUT80), .B(n620), .ZN(n622) );
  NAND2_X1 U700 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U701 ( .A(n624), .B(n623), .ZN(n785) );
  NOR2_X1 U702 ( .A1(n681), .A2(n785), .ZN(n626) );
  NAND2_X1 U703 ( .A1(n625), .A2(n626), .ZN(n628) );
  OR2_X1 U704 ( .A1(n626), .A2(KEYINPUT44), .ZN(n627) );
  NAND2_X1 U705 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U707 ( .A1(n632), .A2(n694), .ZN(n699) );
  INV_X1 U708 ( .A(n699), .ZN(n772) );
  INV_X1 U709 ( .A(KEYINPUT65), .ZN(n633) );
  NAND2_X1 U710 ( .A1(n633), .A2(KEYINPUT2), .ZN(n635) );
  NAND2_X1 U711 ( .A1(n638), .A2(KEYINPUT2), .ZN(n634) );
  NAND2_X1 U712 ( .A1(n634), .A2(KEYINPUT65), .ZN(n637) );
  AND2_X1 U713 ( .A1(n635), .A2(n637), .ZN(n636) );
  NAND2_X1 U714 ( .A1(n701), .A2(n636), .ZN(n641) );
  INV_X1 U715 ( .A(n637), .ZN(n639) );
  OR2_X1 U716 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U717 ( .A1(n641), .A2(n640), .ZN(n649) );
  INV_X1 U718 ( .A(n701), .ZN(n643) );
  INV_X1 U719 ( .A(KEYINPUT2), .ZN(n644) );
  NOR2_X1 U720 ( .A1(n644), .A2(KEYINPUT81), .ZN(n642) );
  OR2_X1 U721 ( .A1(n699), .A2(n644), .ZN(n645) );
  NAND2_X1 U722 ( .A1(n646), .A2(n758), .ZN(n647) );
  NAND2_X1 U723 ( .A1(n752), .A2(G472), .ZN(n652) );
  XNOR2_X1 U724 ( .A(n652), .B(n651), .ZN(n654) );
  INV_X1 U725 ( .A(G952), .ZN(n653) );
  NOR2_X2 U726 ( .A1(n654), .A2(n757), .ZN(n656) );
  XNOR2_X1 U727 ( .A(KEYINPUT63), .B(KEYINPUT93), .ZN(n655) );
  XNOR2_X1 U728 ( .A(n656), .B(n655), .ZN(G57) );
  XOR2_X1 U729 ( .A(n657), .B(G140), .Z(G42) );
  NAND2_X1 U730 ( .A1(n752), .A2(G210), .ZN(n661) );
  XOR2_X1 U731 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n658) );
  XNOR2_X1 U732 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U733 ( .A(n661), .B(n660), .ZN(n662) );
  NOR2_X2 U734 ( .A1(n662), .A2(n757), .ZN(n663) );
  XNOR2_X1 U735 ( .A(n663), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U736 ( .A(KEYINPUT122), .B(KEYINPUT92), .Z(n665) );
  XNOR2_X1 U737 ( .A(KEYINPUT59), .B(KEYINPUT121), .ZN(n664) );
  XOR2_X1 U738 ( .A(n665), .B(n664), .Z(n666) );
  XNOR2_X1 U739 ( .A(n669), .B(n668), .ZN(n670) );
  NOR2_X2 U740 ( .A1(n670), .A2(n757), .ZN(n672) );
  XOR2_X1 U741 ( .A(KEYINPUT123), .B(KEYINPUT60), .Z(n671) );
  XNOR2_X1 U742 ( .A(n672), .B(n671), .ZN(G60) );
  XOR2_X1 U743 ( .A(n673), .B(G122), .Z(G24) );
  XOR2_X1 U744 ( .A(G101), .B(n674), .Z(G3) );
  NOR2_X1 U745 ( .A1(n691), .A2(n678), .ZN(n675) );
  XOR2_X1 U746 ( .A(G104), .B(n675), .Z(G6) );
  XOR2_X1 U747 ( .A(KEYINPUT112), .B(KEYINPUT26), .Z(n677) );
  XNOR2_X1 U748 ( .A(G107), .B(KEYINPUT27), .ZN(n676) );
  XNOR2_X1 U749 ( .A(n677), .B(n676), .ZN(n680) );
  NOR2_X1 U750 ( .A1(n694), .A2(n678), .ZN(n679) );
  XOR2_X1 U751 ( .A(n680), .B(n679), .Z(G9) );
  XOR2_X1 U752 ( .A(G110), .B(n681), .Z(G12) );
  NOR2_X1 U753 ( .A1(n687), .A2(n694), .ZN(n685) );
  XOR2_X1 U754 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n683) );
  XNOR2_X1 U755 ( .A(G128), .B(KEYINPUT29), .ZN(n682) );
  XNOR2_X1 U756 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U757 ( .A(n685), .B(n684), .ZN(G30) );
  XOR2_X1 U758 ( .A(n350), .B(n686), .Z(G45) );
  NOR2_X1 U759 ( .A1(n687), .A2(n691), .ZN(n689) );
  XNOR2_X1 U760 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n688) );
  XNOR2_X1 U761 ( .A(n689), .B(n688), .ZN(n690) );
  XNOR2_X1 U762 ( .A(G146), .B(n690), .ZN(G48) );
  NOR2_X1 U763 ( .A1(n691), .A2(n693), .ZN(n692) );
  XOR2_X1 U764 ( .A(G113), .B(n692), .Z(G15) );
  NOR2_X1 U765 ( .A1(n694), .A2(n693), .ZN(n696) );
  XNOR2_X1 U766 ( .A(G116), .B(KEYINPUT117), .ZN(n695) );
  XNOR2_X1 U767 ( .A(n696), .B(n695), .ZN(G18) );
  XNOR2_X1 U768 ( .A(n697), .B(G125), .ZN(n698) );
  XNOR2_X1 U769 ( .A(n698), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U770 ( .A(G134), .B(n699), .Z(G36) );
  XNOR2_X1 U771 ( .A(KEYINPUT83), .B(KEYINPUT2), .ZN(n700) );
  NAND2_X1 U772 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U773 ( .A(KEYINPUT82), .B(n702), .Z(n704) );
  NOR2_X1 U774 ( .A1(n704), .A2(n703), .ZN(n742) );
  NOR2_X1 U775 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U776 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U777 ( .A(KEYINPUT119), .B(n709), .Z(n713) );
  NOR2_X1 U778 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U779 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U780 ( .A1(n388), .A2(n714), .ZN(n732) );
  NOR2_X1 U781 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U782 ( .A(n717), .B(KEYINPUT50), .ZN(n718) );
  NOR2_X1 U783 ( .A1(n719), .A2(n718), .ZN(n724) );
  NOR2_X1 U784 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U785 ( .A(n722), .B(KEYINPUT49), .ZN(n723) );
  NAND2_X1 U786 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U787 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U788 ( .A(KEYINPUT51), .B(n727), .Z(n728) );
  NAND2_X1 U789 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U790 ( .A(KEYINPUT118), .B(n730), .Z(n731) );
  NOR2_X1 U791 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U792 ( .A(n733), .B(KEYINPUT52), .ZN(n734) );
  NOR2_X1 U793 ( .A1(n735), .A2(n734), .ZN(n738) );
  NOR2_X1 U794 ( .A1(n388), .A2(n736), .ZN(n737) );
  NOR2_X1 U795 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U796 ( .A(n739), .B(KEYINPUT120), .ZN(n740) );
  NAND2_X1 U797 ( .A1(n740), .A2(n775), .ZN(n741) );
  NOR2_X1 U798 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U799 ( .A(n743), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U800 ( .A1(n753), .A2(G469), .ZN(n747) );
  XOR2_X1 U801 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n744) );
  XNOR2_X1 U802 ( .A(n745), .B(n744), .ZN(n746) );
  XNOR2_X1 U803 ( .A(n747), .B(n746), .ZN(n748) );
  NOR2_X1 U804 ( .A1(n748), .A2(n757), .ZN(G54) );
  NAND2_X1 U805 ( .A1(n753), .A2(G478), .ZN(n750) );
  XNOR2_X1 U806 ( .A(n750), .B(n749), .ZN(n751) );
  NOR2_X1 U807 ( .A1(n757), .A2(n751), .ZN(G63) );
  BUF_X1 U808 ( .A(n752), .Z(n753) );
  NAND2_X1 U809 ( .A1(n753), .A2(G217), .ZN(n754) );
  XNOR2_X1 U810 ( .A(n755), .B(n754), .ZN(n756) );
  NOR2_X1 U811 ( .A1(n757), .A2(n756), .ZN(G66) );
  NAND2_X1 U812 ( .A1(n758), .A2(n775), .ZN(n762) );
  NAND2_X1 U813 ( .A1(G953), .A2(G224), .ZN(n759) );
  XNOR2_X1 U814 ( .A(KEYINPUT61), .B(n759), .ZN(n760) );
  NAND2_X1 U815 ( .A1(n760), .A2(G898), .ZN(n761) );
  NAND2_X1 U816 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U817 ( .A(n763), .B(KEYINPUT124), .ZN(n769) );
  XNOR2_X1 U818 ( .A(n765), .B(n764), .ZN(n767) );
  NAND2_X1 U819 ( .A1(n767), .A2(n766), .ZN(n768) );
  XOR2_X1 U820 ( .A(n769), .B(n768), .Z(G69) );
  XNOR2_X1 U821 ( .A(n771), .B(n770), .ZN(n777) );
  AND2_X1 U822 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U823 ( .A(n777), .B(n774), .ZN(n776) );
  NAND2_X1 U824 ( .A1(n776), .A2(n775), .ZN(n782) );
  XNOR2_X1 U825 ( .A(n777), .B(G227), .ZN(n778) );
  XNOR2_X1 U826 ( .A(n778), .B(KEYINPUT125), .ZN(n779) );
  NAND2_X1 U827 ( .A1(n779), .A2(G900), .ZN(n780) );
  NAND2_X1 U828 ( .A1(n780), .A2(G953), .ZN(n781) );
  NAND2_X1 U829 ( .A1(n782), .A2(n781), .ZN(G72) );
  XOR2_X1 U830 ( .A(G137), .B(KEYINPUT126), .Z(n783) );
  XNOR2_X1 U831 ( .A(n784), .B(n783), .ZN(G39) );
  XOR2_X1 U832 ( .A(G119), .B(n785), .Z(G21) );
  XNOR2_X1 U833 ( .A(G131), .B(KEYINPUT127), .ZN(n787) );
  XNOR2_X1 U834 ( .A(n787), .B(n786), .ZN(G33) );
endmodule

