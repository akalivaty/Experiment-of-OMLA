//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 0 1 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 0 1 1 1 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  INV_X1    g0010(.A(G87), .ZN(new_n211));
  INV_X1    g0011(.A(G250), .ZN(new_n212));
  INV_X1    g0012(.A(G116), .ZN(new_n213));
  INV_X1    g0013(.A(G270), .ZN(new_n214));
  OAI22_X1  g0014(.A1(new_n211), .A2(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G77), .A2(G244), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  INV_X1    g0017(.A(G58), .ZN(new_n218));
  INV_X1    g0018(.A(G232), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n216), .B1(new_n202), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI211_X1 g0020(.A(new_n215), .B(new_n220), .C1(G97), .C2(G257), .ZN(new_n221));
  INV_X1    g0021(.A(G107), .ZN(new_n222));
  INV_X1    g0022(.A(G264), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  INV_X1    g0024(.A(KEYINPUT65), .ZN(new_n225));
  INV_X1    g0025(.A(G68), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(KEYINPUT65), .A2(G68), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(new_n207), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n210), .B1(new_n231), .B2(KEYINPUT1), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n231), .A2(KEYINPUT1), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT66), .ZN(new_n234));
  NAND2_X1  g0034(.A1(G1), .A2(G13), .ZN(new_n235));
  INV_X1    g0035(.A(G20), .ZN(new_n236));
  NOR2_X1   g0036(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g0037(.A(new_n201), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n238), .A2(G50), .ZN(new_n239));
  INV_X1    g0039(.A(new_n239), .ZN(new_n240));
  AOI211_X1 g0040(.A(new_n232), .B(new_n234), .C1(new_n237), .C2(new_n240), .ZN(G361));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n219), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT2), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n217), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G250), .B(G257), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G264), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(new_n214), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G358));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(KEYINPUT67), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(new_n211), .ZN(new_n252));
  INV_X1    g0052(.A(G97), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G50), .B(G68), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n255), .B(G58), .ZN(new_n256));
  INV_X1    g0056(.A(G77), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n254), .B(new_n258), .ZN(G351));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n260), .B1(G41), .B2(G45), .ZN(new_n261));
  INV_X1    g0061(.A(G274), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AND2_X1   g0063(.A1(G33), .A2(G41), .ZN(new_n264));
  OR2_X1    g0064(.A1(new_n264), .A2(new_n235), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n265), .A2(new_n261), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n263), .B1(new_n266), .B2(G244), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT70), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n267), .B(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n265), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT3), .B(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G1698), .ZN(new_n272));
  OAI22_X1  g0072(.A1(new_n272), .A2(new_n224), .B1(new_n222), .B2(new_n271), .ZN(new_n273));
  INV_X1    g0073(.A(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT3), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT3), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NOR3_X1   g0078(.A1(new_n278), .A2(new_n219), .A3(G1698), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n270), .B1(new_n273), .B2(new_n279), .ZN(new_n280));
  AND2_X1   g0080(.A1(new_n269), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G179), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G20), .A2(G77), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n236), .A2(G33), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT15), .B(G87), .ZN(new_n286));
  AND2_X1   g0086(.A1(new_n218), .A2(KEYINPUT8), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n218), .A2(KEYINPUT8), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G20), .A2(G33), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  OAI221_X1 g0091(.A(new_n284), .B1(new_n285), .B2(new_n286), .C1(new_n289), .C2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n235), .ZN(new_n294));
  INV_X1    g0094(.A(G13), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n295), .A2(G1), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G20), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  AOI22_X1  g0098(.A1(new_n292), .A2(new_n294), .B1(new_n257), .B2(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n236), .A2(G1), .ZN(new_n300));
  OR2_X1    g0100(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n299), .B1(new_n257), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n269), .A2(new_n280), .ZN(new_n303));
  INV_X1    g0103(.A(G169), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AND3_X1   g0105(.A1(new_n283), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G1698), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n275), .A2(new_n277), .A3(G222), .A4(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n308), .B1(new_n257), .B2(new_n271), .ZN(new_n309));
  AND3_X1   g0109(.A1(new_n271), .A2(G223), .A3(G1698), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n270), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n266), .A2(G226), .ZN(new_n312));
  INV_X1    g0112(.A(new_n263), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n282), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n236), .B(G33), .C1(new_n287), .C2(new_n288), .ZN(new_n317));
  NOR3_X1   g0117(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT69), .B1(new_n318), .B2(new_n236), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n290), .A2(G150), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT69), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n203), .A2(new_n321), .A3(G20), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n317), .A2(new_n319), .A3(new_n320), .A4(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n294), .A2(KEYINPUT68), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT68), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n293), .A2(new_n325), .A3(new_n235), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n298), .A2(new_n202), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n300), .A2(new_n202), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n327), .A2(new_n297), .A3(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n329), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n316), .B(new_n333), .C1(G169), .C2(new_n315), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n306), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n281), .A2(G190), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n302), .B1(new_n303), .B2(G200), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT74), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT14), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n271), .A2(G232), .A3(G1698), .ZN(new_n342));
  NAND2_X1  g0142(.A1(G33), .A2(G97), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n271), .A2(new_n307), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n342), .B(new_n343), .C1(new_n344), .C2(new_n217), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n263), .B1(new_n345), .B2(new_n270), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT13), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n266), .A2(G238), .ZN(new_n348));
  AND3_X1   g0148(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n347), .B1(new_n346), .B2(new_n348), .ZN(new_n350));
  OAI211_X1 g0150(.A(G169), .B(new_n341), .C1(new_n349), .C2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n345), .A2(new_n270), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n352), .A2(new_n313), .A3(new_n348), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(KEYINPUT13), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(G179), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n304), .B1(new_n354), .B2(new_n355), .ZN(new_n357));
  XNOR2_X1  g0157(.A(KEYINPUT74), .B(KEYINPUT14), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n351), .B(new_n356), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT12), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n297), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n226), .B1(new_n301), .B2(KEYINPUT12), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n229), .A2(G20), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NOR3_X1   g0164(.A1(new_n360), .A2(new_n295), .A3(G1), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n362), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  OAI221_X1 g0166(.A(new_n363), .B1(new_n202), .B2(new_n291), .C1(new_n257), .C2(new_n285), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT11), .ZN(new_n368));
  AND3_X1   g0168(.A1(new_n367), .A2(new_n368), .A3(new_n328), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n368), .B1(new_n367), .B2(new_n328), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n361), .B(new_n366), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(KEYINPUT73), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n367), .A2(new_n328), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT11), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n367), .A2(new_n368), .A3(new_n328), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT73), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n376), .A2(new_n377), .A3(new_n361), .A4(new_n366), .ZN(new_n378));
  AND2_X1   g0178(.A1(new_n372), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n359), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n372), .A2(new_n378), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n354), .A2(G190), .A3(new_n355), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT72), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n354), .A2(new_n355), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n383), .B1(new_n384), .B2(G200), .ZN(new_n385));
  INV_X1    g0185(.A(G200), .ZN(new_n386));
  AOI211_X1 g0186(.A(KEYINPUT72), .B(new_n386), .C1(new_n354), .C2(new_n355), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n381), .B(new_n382), .C1(new_n385), .C2(new_n387), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n336), .A2(new_n339), .A3(new_n380), .A4(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT80), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT18), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n328), .A2(new_n298), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n289), .A2(new_n300), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n392), .A2(new_n393), .B1(new_n298), .B2(new_n289), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  AND2_X1   g0195(.A1(new_n293), .A2(new_n235), .ZN(new_n396));
  OAI21_X1  g0196(.A(KEYINPUT7), .B1(new_n271), .B2(G20), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT7), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT75), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT75), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT7), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n278), .A2(new_n402), .A3(new_n236), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n397), .A2(new_n403), .A3(G68), .ZN(new_n404));
  INV_X1    g0204(.A(G159), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n291), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n227), .A2(G58), .A3(new_n228), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n238), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n406), .B1(new_n408), .B2(G20), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n404), .A2(new_n409), .A3(KEYINPUT16), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT76), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT76), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n404), .A2(new_n409), .A3(new_n412), .A4(KEYINPUT16), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n396), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT16), .ZN(new_n415));
  AOI21_X1  g0215(.A(G20), .B1(new_n275), .B2(new_n277), .ZN(new_n416));
  XNOR2_X1  g0216(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT77), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT77), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n402), .B(new_n419), .C1(new_n271), .C2(G20), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT78), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n276), .B2(G33), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n274), .A2(KEYINPUT78), .A3(KEYINPUT3), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n423), .A2(new_n277), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n425), .A2(KEYINPUT7), .A3(new_n236), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n229), .B1(new_n421), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n409), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n415), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n395), .B1(new_n414), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n266), .A2(G232), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n271), .A2(G226), .A3(G1698), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n271), .A2(G223), .A3(new_n307), .ZN(new_n433));
  NAND2_X1  g0233(.A1(G33), .A2(G87), .ZN(new_n434));
  AND3_X1   g0234(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n431), .B(new_n313), .C1(new_n435), .C2(new_n265), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(G169), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n437), .B1(new_n282), .B2(new_n436), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n391), .B1(new_n430), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n411), .A2(new_n413), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n441), .A2(new_n429), .A3(new_n294), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n394), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n443), .A2(KEYINPUT18), .A3(new_n438), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n436), .A2(G200), .ZN(new_n446));
  INV_X1    g0246(.A(G190), .ZN(new_n447));
  OR2_X1    g0247(.A1(new_n436), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n442), .A2(new_n394), .A3(new_n446), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT17), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT17), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n430), .A2(new_n451), .A3(new_n446), .A4(new_n448), .ZN(new_n452));
  AND3_X1   g0252(.A1(new_n450), .A2(KEYINPUT79), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT79), .B1(new_n450), .B2(new_n452), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n445), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n389), .B1(new_n390), .B2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT9), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n333), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT71), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n311), .A2(new_n312), .A3(G190), .A4(new_n313), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n329), .A2(KEYINPUT9), .A3(new_n330), .A4(new_n332), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n458), .A2(new_n459), .A3(new_n460), .A4(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT10), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n314), .A2(G200), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n458), .A2(new_n465), .A3(new_n460), .A4(new_n461), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n466), .A2(new_n462), .A3(new_n463), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n445), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n450), .A2(new_n452), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT79), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n450), .A2(KEYINPUT79), .A3(new_n452), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n471), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n470), .B1(new_n476), .B2(KEYINPUT80), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n456), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G283), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n480), .B(new_n236), .C1(G33), .C2(new_n253), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n396), .B1(KEYINPUT86), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n213), .A2(G20), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n274), .A2(G97), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT86), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n484), .A2(new_n485), .A3(new_n236), .A4(new_n480), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n482), .A2(KEYINPUT20), .A3(new_n483), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n481), .A2(KEYINPUT86), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n488), .A2(new_n294), .A3(new_n483), .A4(new_n486), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT20), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n296), .A2(G20), .A3(new_n213), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n260), .A2(G33), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n396), .A2(new_n297), .A3(G116), .A4(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n492), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n278), .A2(G303), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n497), .B1(new_n272), .B2(new_n223), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n275), .A2(new_n277), .A3(new_n307), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n499), .A2(G257), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n270), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT5), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G41), .ZN(new_n503));
  INV_X1    g0303(.A(G41), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT5), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n503), .A2(new_n505), .A3(new_n260), .A4(G45), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n506), .A2(new_n265), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G270), .ZN(new_n508));
  INV_X1    g0308(.A(new_n505), .ZN(new_n509));
  OR2_X1    g0309(.A1(new_n509), .A2(KEYINPUT83), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n260), .A2(G45), .A3(G274), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n511), .B1(new_n509), .B2(KEYINPUT83), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n510), .A2(new_n503), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n501), .A2(new_n508), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n496), .A2(G169), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(KEYINPUT21), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT21), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n496), .A2(new_n517), .A3(G169), .A4(new_n514), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n492), .A2(new_n493), .A3(new_n495), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(new_n514), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n516), .A2(new_n518), .B1(new_n520), .B2(G179), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n514), .A2(G200), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n522), .B(new_n519), .C1(new_n447), .C2(new_n514), .ZN(new_n523));
  AND2_X1   g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n275), .A2(new_n277), .A3(G244), .A4(new_n307), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT4), .ZN(new_n526));
  AND3_X1   g0326(.A1(new_n525), .A2(KEYINPUT81), .A3(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(KEYINPUT82), .B1(new_n525), .B2(new_n526), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT82), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n499), .A2(new_n529), .A3(KEYINPUT4), .A4(G244), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n527), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT81), .B1(new_n525), .B2(new_n526), .ZN(new_n532));
  NOR3_X1   g0332(.A1(new_n278), .A2(new_n212), .A3(new_n307), .ZN(new_n533));
  INV_X1    g0333(.A(new_n480), .ZN(new_n534));
  NOR3_X1   g0334(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n265), .B1(new_n531), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n507), .A2(G257), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n513), .ZN(new_n538));
  OAI21_X1  g0338(.A(G169), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n530), .A2(new_n528), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n525), .A2(new_n526), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT81), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n534), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n533), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n525), .A2(KEYINPUT81), .A3(new_n526), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n540), .A2(new_n543), .A3(new_n544), .A4(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n270), .ZN(new_n547));
  INV_X1    g0347(.A(new_n538), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n547), .A2(G179), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n539), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n290), .A2(G77), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n222), .A2(KEYINPUT6), .A3(G97), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n253), .A2(new_n222), .ZN(new_n553));
  NOR2_X1   g0353(.A1(G97), .A2(G107), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n552), .B1(new_n555), .B2(KEYINPUT6), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(G20), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n425), .A2(new_n236), .ZN(new_n558));
  AOI22_X1  g0358(.A1(KEYINPUT7), .A2(new_n558), .B1(new_n418), .B2(new_n420), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n551), .B(new_n557), .C1(new_n559), .C2(new_n222), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n294), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n297), .A2(G97), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n327), .A2(new_n297), .A3(new_n494), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G97), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n561), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n550), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n275), .A2(new_n277), .A3(G244), .A4(G1698), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n275), .A2(new_n277), .A3(G238), .A4(new_n307), .ZN(new_n570));
  NAND2_X1  g0370(.A1(G33), .A2(G116), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n270), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT84), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n260), .A2(G45), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n575), .B(G250), .C1(new_n264), .C2(new_n235), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n574), .B1(new_n576), .B2(new_n511), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n576), .A2(new_n574), .A3(new_n511), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n573), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(G200), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n554), .A2(new_n211), .ZN(new_n582));
  NOR2_X1   g0382(.A1(KEYINPUT85), .A2(KEYINPUT19), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n343), .A2(new_n236), .ZN(new_n585));
  NAND2_X1  g0385(.A1(KEYINPUT85), .A2(KEYINPUT19), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n582), .A2(new_n584), .A3(new_n585), .A4(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n586), .ZN(new_n588));
  OAI22_X1  g0388(.A1(new_n588), .A2(new_n583), .B1(new_n285), .B2(new_n253), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n275), .A2(new_n277), .A3(new_n236), .A4(G68), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n587), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n294), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n298), .A2(new_n286), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n327), .A2(G87), .A3(new_n297), .A4(new_n494), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n573), .B(G190), .C1(new_n577), .C2(new_n579), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n581), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n573), .B(new_n282), .C1(new_n577), .C2(new_n579), .ZN(new_n598));
  INV_X1    g0398(.A(new_n286), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n327), .A2(new_n297), .A3(new_n599), .A4(new_n494), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n592), .A2(new_n600), .A3(new_n593), .ZN(new_n601));
  INV_X1    g0401(.A(new_n577), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n602), .A2(new_n578), .B1(new_n572), .B2(new_n270), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n598), .B(new_n601), .C1(new_n603), .C2(G169), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n597), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n562), .B1(new_n560), .B2(new_n294), .ZN(new_n606));
  OAI21_X1  g0406(.A(G200), .B1(new_n536), .B2(new_n538), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n547), .A2(G190), .A3(new_n548), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n606), .A2(new_n607), .A3(new_n608), .A4(new_n566), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n568), .A2(new_n605), .A3(new_n609), .ZN(new_n610));
  AND2_X1   g0410(.A1(KEYINPUT22), .A2(G87), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n275), .A2(new_n277), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n571), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n236), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT24), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n275), .A2(new_n277), .A3(new_n236), .A4(G87), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT22), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT87), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(KEYINPUT23), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT23), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(KEYINPUT87), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n620), .A2(new_n622), .A3(G20), .A4(new_n222), .ZN(new_n623));
  OAI211_X1 g0423(.A(KEYINPUT87), .B(new_n621), .C1(new_n236), .C2(G107), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n614), .A2(new_n615), .A3(new_n618), .A4(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n613), .A2(new_n236), .B1(new_n617), .B2(new_n616), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n615), .B1(new_n628), .B2(new_n625), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n294), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n564), .A2(new_n222), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n298), .A2(new_n222), .ZN(new_n633));
  XNOR2_X1  g0433(.A(new_n633), .B(KEYINPUT25), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n630), .A2(new_n632), .A3(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n271), .A2(G257), .A3(G1698), .ZN(new_n637));
  NAND2_X1  g0437(.A1(G33), .A2(G294), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n275), .A2(new_n277), .A3(G250), .A4(new_n307), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n270), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n507), .A2(G264), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n641), .A2(new_n642), .A3(G179), .A4(new_n513), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n643), .A2(KEYINPUT88), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT88), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n641), .A2(new_n642), .A3(new_n513), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n645), .B1(new_n646), .B2(G169), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n643), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n636), .A2(new_n644), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(KEYINPUT89), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT89), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n636), .A2(new_n648), .A3(new_n651), .A4(new_n644), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n641), .A2(new_n642), .A3(G190), .A4(new_n513), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n630), .A2(new_n653), .A3(new_n632), .A4(new_n635), .ZN(new_n654));
  INV_X1    g0454(.A(new_n646), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n655), .A2(new_n386), .ZN(new_n656));
  OAI21_X1  g0456(.A(KEYINPUT90), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n271), .A2(new_n611), .B1(G33), .B2(G116), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n618), .B(new_n625), .C1(new_n658), .C2(G20), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(KEYINPUT24), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n626), .ZN(new_n661));
  AOI211_X1 g0461(.A(new_n631), .B(new_n634), .C1(new_n661), .C2(new_n294), .ZN(new_n662));
  INV_X1    g0462(.A(new_n656), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT90), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n662), .A2(new_n663), .A3(new_n664), .A4(new_n653), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n650), .A2(new_n652), .B1(new_n657), .B2(new_n665), .ZN(new_n666));
  AND4_X1   g0466(.A1(new_n479), .A2(new_n524), .A3(new_n610), .A4(new_n666), .ZN(G372));
  NAND2_X1  g0467(.A1(new_n657), .A2(new_n665), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n521), .A2(new_n649), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n610), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n567), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n550), .A2(KEYINPUT91), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT91), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n539), .A2(new_n549), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n671), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(KEYINPUT26), .B1(new_n675), .B2(new_n605), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n550), .A2(new_n605), .A3(new_n567), .A4(KEYINPUT26), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT92), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n606), .A2(new_n566), .B1(new_n539), .B2(new_n549), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n680), .A2(KEYINPUT92), .A3(KEYINPUT26), .A4(new_n605), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n670), .B(new_n604), .C1(new_n676), .C2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n479), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n283), .A2(new_n302), .A3(new_n305), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n380), .A2(new_n685), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n388), .B(new_n686), .C1(new_n453), .C2(new_n454), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n445), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT93), .ZN(new_n689));
  AND3_X1   g0489(.A1(new_n466), .A2(new_n462), .A3(new_n463), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n466), .B1(new_n463), .B2(new_n462), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n689), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n468), .A2(KEYINPUT93), .A3(new_n469), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n335), .B1(new_n688), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n684), .A2(new_n695), .ZN(G369));
  INV_X1    g0496(.A(new_n521), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n295), .A2(G20), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n260), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n699), .A2(KEYINPUT27), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(KEYINPUT27), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(G213), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT94), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G343), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(new_n519), .ZN(new_n705));
  MUX2_X1   g0505(.A(new_n524), .B(new_n697), .S(new_n705), .Z(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(G330), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n649), .A2(new_n704), .ZN(new_n708));
  INV_X1    g0508(.A(new_n704), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n636), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n708), .B1(new_n666), .B2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n666), .A2(new_n697), .A3(new_n704), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n631), .B1(new_n661), .B2(new_n294), .ZN(new_n715));
  AOI22_X1  g0515(.A1(new_n715), .A2(new_n635), .B1(new_n643), .B2(new_n647), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n716), .A2(new_n644), .A3(new_n704), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n713), .A2(new_n718), .ZN(G399));
  INV_X1    g0519(.A(new_n208), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(G41), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n582), .A2(G116), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n722), .A2(G1), .A3(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n724), .B1(new_n239), .B2(new_n722), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT28), .ZN(new_n726));
  INV_X1    g0526(.A(G330), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT30), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n547), .A2(G179), .A3(new_n655), .A4(new_n548), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n603), .A2(new_n508), .A3(new_n501), .ZN(new_n730));
  OAI211_X1 g0530(.A(KEYINPUT96), .B(new_n728), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n655), .A2(G179), .A3(new_n603), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n732), .B(new_n514), .C1(new_n536), .C2(new_n538), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n536), .A2(new_n282), .A3(new_n538), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n728), .A2(KEYINPUT96), .ZN(new_n735));
  INV_X1    g0535(.A(new_n730), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n734), .A2(new_n655), .A3(new_n735), .A4(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n731), .A2(new_n733), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(KEYINPUT31), .B1(new_n738), .B2(new_n709), .ZN(new_n739));
  XOR2_X1   g0539(.A(KEYINPUT95), .B(KEYINPUT31), .Z(new_n740));
  AND2_X1   g0540(.A1(new_n738), .A2(new_n709), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n666), .A2(new_n524), .A3(new_n610), .A4(new_n704), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n727), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n683), .A2(new_n704), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT29), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n651), .B1(new_n716), .B2(new_n644), .ZN(new_n748));
  INV_X1    g0548(.A(new_n652), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n521), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n750), .A2(new_n610), .A3(new_n668), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n550), .A2(new_n605), .A3(new_n567), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT26), .ZN(new_n753));
  AOI21_X1  g0553(.A(KEYINPUT97), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n674), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n673), .B1(new_n539), .B2(new_n549), .ZN(new_n756));
  OAI211_X1 g0556(.A(new_n605), .B(new_n567), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n754), .B1(new_n757), .B2(new_n753), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n675), .A2(KEYINPUT97), .A3(KEYINPUT26), .A4(new_n605), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n751), .A2(new_n758), .A3(new_n604), .A4(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n760), .A2(KEYINPUT29), .A3(new_n704), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n744), .B1(new_n747), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n726), .B1(new_n762), .B2(G1), .ZN(G364));
  NOR4_X1   g0563(.A1(new_n236), .A2(new_n282), .A3(new_n447), .A4(new_n386), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(G326), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n236), .A2(G179), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n767), .A2(new_n447), .A3(G200), .ZN(new_n768));
  INV_X1    g0568(.A(G283), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n765), .A2(new_n766), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n236), .A2(new_n282), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n771), .A2(G190), .A3(new_n386), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n271), .B(new_n770), .C1(G322), .C2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G190), .A2(G200), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G311), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n771), .A2(new_n447), .A3(G200), .ZN(new_n778));
  XOR2_X1   g0578(.A(KEYINPUT33), .B(G317), .Z(new_n779));
  NAND3_X1  g0579(.A1(new_n767), .A2(G190), .A3(G200), .ZN(new_n780));
  INV_X1    g0580(.A(G303), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n778), .A2(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n447), .A2(G179), .A3(G200), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n236), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n782), .B1(G294), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n767), .A2(new_n775), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n787), .B(KEYINPUT103), .Z(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G329), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n774), .A2(new_n777), .A3(new_n786), .A4(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n787), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G159), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT32), .ZN(new_n794));
  INV_X1    g0594(.A(new_n778), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n794), .B1(G68), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n271), .B1(new_n772), .B2(new_n218), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(G77), .B2(new_n776), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n780), .A2(new_n211), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n768), .A2(new_n222), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n799), .B(new_n800), .C1(G50), .C2(new_n764), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n796), .A2(new_n798), .A3(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n784), .A2(new_n253), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n791), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n235), .B1(G20), .B2(new_n304), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n260), .B1(new_n698), .B2(G45), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n721), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT98), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n208), .A2(new_n271), .ZN(new_n811));
  INV_X1    g0611(.A(G355), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n811), .A2(new_n812), .B1(G116), .B2(new_n208), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT99), .Z(new_n814));
  NOR2_X1   g0614(.A1(new_n720), .A2(new_n271), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT100), .ZN(new_n816));
  INV_X1    g0616(.A(G45), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n816), .B1(new_n817), .B2(new_n258), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n239), .A2(G45), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n814), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(G13), .A2(G33), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(G20), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n823), .A2(new_n805), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT101), .Z(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT102), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n810), .B1(new_n820), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n823), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n806), .B(new_n827), .C1(new_n706), .C2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n707), .A2(new_n810), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n706), .A2(G330), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(G396));
  NAND4_X1  g0632(.A1(new_n283), .A2(new_n302), .A3(new_n305), .A4(new_n704), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n337), .A2(new_n338), .B1(new_n302), .B2(new_n709), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n833), .B1(new_n306), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n745), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n835), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n683), .A2(new_n704), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(new_n744), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n810), .ZN(new_n841));
  AOI22_X1  g0641(.A1(G137), .A2(new_n764), .B1(new_n776), .B2(G159), .ZN(new_n842));
  INV_X1    g0642(.A(G143), .ZN(new_n843));
  INV_X1    g0643(.A(G150), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n842), .B1(new_n843), .B2(new_n772), .C1(new_n844), .C2(new_n778), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT34), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n271), .B1(new_n768), .B2(new_n226), .C1(new_n784), .C2(new_n218), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(new_n789), .B2(G132), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n846), .B(new_n848), .C1(new_n202), .C2(new_n780), .ZN(new_n849));
  INV_X1    g0649(.A(G294), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n772), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n776), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n278), .B1(new_n852), .B2(new_n213), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n803), .B(new_n853), .C1(G283), .C2(new_n795), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n765), .A2(new_n781), .B1(new_n780), .B2(new_n222), .ZN(new_n855));
  INV_X1    g0655(.A(new_n768), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n855), .B1(G87), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(G311), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n854), .B(new_n857), .C1(new_n858), .C2(new_n788), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n849), .B1(new_n851), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n810), .B1(new_n860), .B2(new_n805), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n805), .A2(new_n821), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n861), .B1(G77), .B2(new_n863), .C1(new_n837), .C2(new_n822), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n841), .A2(new_n864), .ZN(G384));
  NAND2_X1  g0665(.A1(new_n738), .A2(new_n709), .ZN(new_n866));
  INV_X1    g0666(.A(new_n740), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n738), .A2(KEYINPUT31), .A3(new_n709), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n743), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n380), .A2(new_n388), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n381), .A2(new_n704), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n380), .B(new_n388), .C1(new_n381), .C2(new_n704), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n835), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT16), .B1(new_n404), .B2(new_n409), .ZN(new_n877));
  AOI211_X1 g0677(.A(new_n327), .B(new_n877), .C1(new_n411), .C2(new_n413), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n703), .B1(new_n878), .B2(new_n395), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n455), .A2(new_n880), .ZN(new_n881));
  OAI22_X1  g0681(.A1(new_n878), .A2(new_n395), .B1(new_n438), .B2(new_n703), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n449), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(KEYINPUT37), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n443), .A2(new_n438), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n443), .A2(new_n703), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT37), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n885), .A2(new_n886), .A3(new_n887), .A4(new_n449), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT38), .B1(new_n881), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT38), .ZN(new_n892));
  AOI211_X1 g0692(.A(new_n892), .B(new_n889), .C1(new_n455), .C2(new_n880), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n876), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT40), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g0696(.A(KEYINPUT105), .B(KEYINPUT38), .ZN(new_n897));
  INV_X1    g0697(.A(new_n886), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n450), .A2(KEYINPUT106), .A3(new_n452), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n445), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT106), .B1(new_n450), .B2(new_n452), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n885), .A2(new_n886), .A3(new_n449), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(KEYINPUT37), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n888), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n897), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  OAI211_X1 g0706(.A(KEYINPUT40), .B(new_n876), .C1(new_n893), .C2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n896), .A2(new_n907), .ZN(new_n908));
  XOR2_X1   g0708(.A(new_n908), .B(KEYINPUT107), .Z(new_n909));
  NAND2_X1  g0709(.A1(new_n479), .A2(new_n870), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n909), .B(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(G330), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n380), .A2(new_n709), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT39), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n890), .B1(new_n476), .B2(new_n879), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n892), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n881), .A2(KEYINPUT38), .A3(new_n890), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NOR3_X1   g0718(.A1(new_n893), .A2(KEYINPUT39), .A3(new_n906), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n913), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n833), .A2(KEYINPUT104), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n833), .A2(KEYINPUT104), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n838), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n873), .A2(new_n874), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n923), .B(new_n924), .C1(new_n893), .C2(new_n891), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n445), .A2(new_n703), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n920), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n479), .A2(new_n747), .A3(new_n761), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n695), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n928), .B(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n912), .B(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n260), .B2(new_n698), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n213), .B1(new_n556), .B2(KEYINPUT35), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n934), .B(new_n237), .C1(KEYINPUT35), .C2(new_n556), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT36), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n240), .A2(G77), .A3(new_n407), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(G50), .B2(new_n226), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n938), .A2(G1), .A3(new_n295), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n933), .A2(new_n936), .A3(new_n939), .ZN(G367));
  NAND2_X1  g0740(.A1(new_n675), .A2(new_n709), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n568), .B(new_n609), .C1(new_n671), .C2(new_n704), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n650), .A2(new_n652), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n568), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n704), .ZN(new_n947));
  OAI21_X1  g0747(.A(KEYINPUT42), .B1(new_n944), .B2(new_n714), .ZN(new_n948));
  OR3_X1    g0748(.A1(new_n944), .A2(KEYINPUT42), .A3(new_n714), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n712), .A2(new_n943), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n605), .B1(new_n595), .B2(new_n704), .ZN(new_n952));
  OR3_X1    g0752(.A1(new_n704), .A2(new_n604), .A3(new_n595), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n955));
  AND3_X1   g0755(.A1(new_n950), .A2(new_n951), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n951), .B1(new_n950), .B2(new_n955), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  OR3_X1    g0759(.A1(new_n956), .A2(new_n957), .A3(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n959), .B1(new_n956), .B2(new_n957), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n721), .B(KEYINPUT41), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n711), .B1(new_n521), .B2(new_n709), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n714), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(new_n707), .Z(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n762), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n718), .A2(new_n943), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT44), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n718), .A2(new_n943), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT45), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n971), .B(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n712), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n970), .A2(new_n713), .A3(new_n973), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n968), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n963), .B1(new_n977), .B2(new_n762), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n960), .B(new_n961), .C1(new_n978), .C2(new_n808), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n856), .A2(G77), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n405), .B2(new_n778), .ZN(new_n981));
  INV_X1    g0781(.A(G137), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n271), .B1(new_n982), .B2(new_n787), .C1(new_n852), .C2(new_n202), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n981), .B(new_n983), .C1(G143), .C2(new_n764), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n784), .A2(new_n226), .B1(new_n772), .B2(new_n844), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT108), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n984), .B(new_n986), .C1(new_n218), .C2(new_n780), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n852), .A2(new_n769), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n785), .A2(G107), .B1(new_n856), .B2(G97), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n850), .B2(new_n778), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(G311), .B2(new_n764), .ZN(new_n991));
  INV_X1    g0791(.A(new_n780), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n992), .A2(KEYINPUT46), .A3(G116), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n278), .B1(new_n772), .B2(new_n781), .ZN(new_n994));
  AOI21_X1  g0794(.A(KEYINPUT46), .B1(new_n992), .B2(G116), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n994), .B(new_n995), .C1(G317), .C2(new_n792), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n991), .A2(new_n993), .A3(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n987), .B1(new_n988), .B2(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n999));
  XNOR2_X1  g0799(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n810), .B1(new_n1000), .B2(new_n805), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n825), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n816), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1002), .B1(new_n208), .B2(new_n286), .C1(new_n1003), .C2(new_n248), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1001), .B(new_n1004), .C1(new_n828), .C2(new_n954), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n979), .A2(new_n1005), .ZN(G387));
  AOI22_X1  g0806(.A1(G322), .A2(new_n764), .B1(new_n776), .B2(G303), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n773), .A2(G317), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1007), .B(new_n1008), .C1(new_n858), .C2(new_n778), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT48), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1010), .B1(new_n769), .B2(new_n784), .C1(new_n850), .C2(new_n780), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT49), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n271), .B1(new_n856), .B2(G116), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1012), .B(new_n1013), .C1(new_n766), .C2(new_n787), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(KEYINPUT111), .B(G150), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n271), .B1(new_n787), .B2(new_n1015), .C1(new_n852), .C2(new_n226), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n257), .A2(new_n780), .B1(new_n768), .B2(new_n253), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n765), .A2(new_n405), .B1(new_n289), .B2(new_n778), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(new_n599), .B2(new_n785), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1018), .B(new_n1020), .C1(new_n202), .C2(new_n772), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1014), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n810), .B1(new_n1022), .B2(new_n805), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n711), .A2(new_n823), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n245), .A2(new_n817), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n1026), .A2(KEYINPUT110), .ZN(new_n1027));
  OR3_X1    g0827(.A1(new_n289), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1028));
  AOI211_X1 g0828(.A(G116), .B(new_n582), .C1(G68), .C2(G77), .ZN(new_n1029));
  OAI21_X1  g0829(.A(KEYINPUT50), .B1(new_n289), .B2(G50), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .A4(new_n817), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1026), .A2(KEYINPUT110), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1027), .A2(new_n816), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1033), .B1(G107), .B2(new_n208), .C1(new_n723), .C2(new_n811), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1025), .B1(new_n826), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n966), .B2(new_n808), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n721), .B1(new_n966), .B2(new_n762), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1036), .B1(new_n968), .B2(new_n1037), .ZN(G393));
  NAND2_X1  g0838(.A1(new_n975), .A2(new_n976), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n722), .B1(new_n1039), .B2(new_n967), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1040), .A2(new_n977), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1002), .B1(new_n253), .B2(new_n208), .C1(new_n254), .C2(new_n1003), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n852), .A2(new_n850), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n271), .B(new_n1043), .C1(G322), .C2(new_n792), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n795), .A2(G303), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n800), .B1(G116), .B2(new_n785), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n992), .A2(G283), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n773), .A2(G311), .B1(new_n764), .B2(G317), .ZN(new_n1049));
  XOR2_X1   g0849(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n1050));
  XNOR2_X1  g0850(.A(new_n1049), .B(new_n1050), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n765), .A2(new_n844), .B1(new_n405), .B2(new_n772), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT51), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n780), .A2(new_n229), .B1(new_n787), .B2(new_n843), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(KEYINPUT112), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n289), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n278), .B1(new_n1056), .B2(new_n776), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1053), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n784), .A2(new_n257), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(G50), .B2(new_n795), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1060), .B1(KEYINPUT112), .B2(new_n1054), .C1(new_n211), .C2(new_n768), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n1048), .A2(new_n1051), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n810), .B1(new_n1062), .B2(new_n805), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1042), .B(new_n1063), .C1(new_n943), .C2(new_n828), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n1039), .B2(new_n807), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1041), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(G390));
  OR2_X1    g0867(.A1(new_n306), .A2(new_n834), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n760), .A2(new_n704), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n833), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n924), .ZN(new_n1071));
  AND2_X1   g0871(.A1(new_n902), .A2(new_n905), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n917), .B1(new_n1072), .B2(new_n897), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n913), .B(KEYINPUT114), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1071), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(KEYINPUT39), .B1(new_n891), .B2(new_n893), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n917), .B(new_n914), .C1(new_n1072), .C2(new_n897), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n913), .B1(new_n923), .B2(new_n924), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1075), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n835), .A2(new_n727), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n870), .A2(new_n924), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n742), .A2(new_n743), .ZN(new_n1084));
  AND3_X1   g0884(.A1(new_n1084), .A2(new_n924), .A3(new_n1081), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1075), .B(new_n1085), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT116), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n924), .B1(new_n870), .B2(new_n1081), .ZN(new_n1089));
  NOR3_X1   g0889(.A1(new_n1070), .A2(new_n1085), .A3(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1068), .A2(G330), .A3(new_n833), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(new_n742), .B2(new_n743), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1082), .B1(new_n1092), .B2(new_n924), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n923), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(KEYINPUT115), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT115), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1093), .A2(new_n1096), .A3(new_n923), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1090), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n456), .A2(new_n477), .A3(G330), .A4(new_n870), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n747), .A2(new_n761), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n695), .B(new_n1099), .C1(new_n1100), .C2(new_n478), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1088), .B1(new_n1098), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1087), .A2(new_n1102), .ZN(new_n1103));
  OR3_X1    g0903(.A1(new_n1070), .A2(new_n1085), .A3(new_n1089), .ZN(new_n1104));
  AND3_X1   g0904(.A1(new_n1093), .A2(new_n1096), .A3(new_n923), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1096), .B1(new_n1093), .B2(new_n923), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1104), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1101), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1109), .A2(new_n1083), .A3(new_n1088), .A4(new_n1086), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1103), .A2(new_n721), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(G132), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n271), .B1(new_n772), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(new_n789), .B2(G125), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n768), .A2(new_n202), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n784), .A2(new_n405), .B1(new_n778), .B2(new_n982), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n1115), .B(new_n1116), .C1(G128), .C2(new_n764), .ZN(new_n1117));
  XOR2_X1   g0917(.A(KEYINPUT54), .B(G143), .Z(new_n1118));
  NAND2_X1  g0918(.A1(new_n776), .A2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n780), .A2(new_n1015), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT53), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1114), .A2(new_n1117), .A3(new_n1119), .A4(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n278), .B1(new_n852), .B2(new_n253), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n799), .B(new_n1123), .C1(G68), .C2(new_n856), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n778), .A2(new_n222), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n1125), .B(new_n1059), .C1(G283), .C2(new_n764), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1124), .B(new_n1126), .C1(new_n850), .C2(new_n788), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n772), .A2(new_n213), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1122), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n810), .B1(new_n1129), .B2(new_n805), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n1078), .B2(new_n822), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(new_n289), .B2(new_n862), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(new_n1087), .B2(new_n808), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1111), .A2(new_n1133), .ZN(G378));
  NAND2_X1  g0934(.A1(new_n870), .A2(new_n875), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(new_n916), .B2(new_n917), .ZN(new_n1136));
  OAI211_X1 g0936(.A(G330), .B(new_n907), .C1(new_n1136), .C2(KEYINPUT40), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT56), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n692), .A2(new_n334), .A3(new_n693), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n703), .A2(new_n333), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT55), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n692), .A2(new_n693), .A3(new_n334), .A4(new_n1140), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1143), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1138), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(KEYINPUT55), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1149), .A2(KEYINPUT56), .A3(new_n1150), .ZN(new_n1151));
  AND2_X1   g0951(.A1(new_n1147), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1137), .A2(new_n1153), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n896), .A2(G330), .A3(new_n1152), .A4(new_n907), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n928), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n920), .A2(new_n925), .A3(new_n927), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1158), .A2(new_n1155), .A3(new_n1154), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n808), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n504), .B1(new_n780), .B2(new_n257), .C1(new_n222), .C2(new_n772), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n278), .B1(new_n226), .B2(new_n784), .C1(new_n852), .C2(new_n286), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n1162), .B(new_n1163), .C1(G283), .C2(new_n789), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n795), .A2(G97), .B1(new_n764), .B2(G116), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1164), .B(new_n1165), .C1(new_n218), .C2(new_n768), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT58), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n504), .B1(new_n276), .B2(new_n274), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n1166), .A2(new_n1167), .B1(new_n202), .B2(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT117), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G128), .A2(new_n773), .B1(new_n992), .B2(new_n1118), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT119), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n795), .A2(G132), .B1(new_n776), .B2(G137), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT118), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n785), .A2(G150), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n764), .A2(G125), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1172), .A2(new_n1174), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  XOR2_X1   g0977(.A(new_n1177), .B(KEYINPUT59), .Z(new_n1178));
  AOI21_X1  g0978(.A(G41), .B1(new_n856), .B2(G159), .ZN(new_n1179));
  AOI21_X1  g0979(.A(G33), .B1(new_n792), .B2(G124), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1170), .B(new_n1181), .C1(new_n1167), .C2(new_n1166), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n810), .B1(new_n1182), .B2(new_n805), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1183), .B1(G50), .B2(new_n863), .C1(new_n1153), .C2(new_n822), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1161), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1082), .ZN(new_n1187));
  AND2_X1   g0987(.A1(new_n923), .A2(new_n924), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1076), .B(new_n1077), .C1(new_n1188), .C2(new_n913), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1187), .B1(new_n1189), .B2(new_n1075), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1086), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1107), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1192), .A2(new_n1108), .B1(new_n1159), .B2(new_n1157), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n721), .B1(new_n1193), .B2(KEYINPUT57), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1098), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1195));
  OAI21_X1  g0995(.A(KEYINPUT57), .B1(new_n1195), .B2(new_n1101), .ZN(new_n1196));
  AOI21_X1  g0996(.A(KEYINPUT120), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1158), .B1(new_n1155), .B2(new_n1154), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT120), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1196), .B1(new_n1198), .B2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1186), .B1(new_n1194), .B2(new_n1203), .ZN(G375));
  OAI211_X1 g1004(.A(new_n1104), .B(new_n1101), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1109), .A2(new_n962), .A3(new_n1205), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT121), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n784), .A2(new_n202), .B1(new_n768), .B2(new_n218), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n278), .B(new_n1208), .C1(G150), .C2(new_n776), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n765), .A2(new_n1112), .B1(new_n780), .B2(new_n405), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n795), .B2(new_n1118), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n789), .A2(G128), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n773), .A2(G137), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1209), .A2(new_n1211), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n789), .A2(G303), .B1(G97), .B2(new_n992), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1215), .A2(KEYINPUT122), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n980), .B1(new_n286), .B2(new_n784), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n278), .B1(new_n769), .B2(new_n772), .C1(new_n852), .C2(new_n222), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1217), .B(new_n1218), .C1(G116), .C2(new_n795), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1215), .A2(KEYINPUT122), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1216), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n765), .A2(new_n850), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1214), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n810), .B1(new_n1223), .B2(new_n805), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n924), .B2(new_n822), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n226), .B2(new_n862), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n1107), .B2(new_n808), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1207), .A2(new_n1227), .ZN(G381));
  INV_X1    g1028(.A(new_n1159), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n1195), .A2(new_n1101), .B1(new_n1229), .B2(new_n1199), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT57), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n722), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1192), .A2(new_n1108), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1233), .B(KEYINPUT57), .C1(new_n1197), .C2(new_n1201), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1185), .B1(new_n1232), .B2(new_n1234), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1111), .A2(new_n1133), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1066), .A2(new_n1005), .A3(new_n979), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(G393), .A2(G396), .ZN(new_n1239));
  INV_X1    g1039(.A(G384), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1241), .B(KEYINPUT123), .ZN(new_n1242));
  OR4_X1    g1042(.A1(G381), .A2(new_n1237), .A3(new_n1238), .A4(new_n1242), .ZN(G407));
  OAI211_X1 g1043(.A(G407), .B(G213), .C1(G343), .C2(new_n1237), .ZN(G409));
  XOR2_X1   g1044(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1245));
  INV_X1    g1045(.A(G213), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1246), .A2(G343), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n808), .B1(new_n1197), .B2(new_n1201), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1160), .B(new_n962), .C1(new_n1101), .C2(new_n1195), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1236), .A2(new_n1184), .A3(new_n1249), .A4(new_n1250), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1248), .B(new_n1251), .C1(new_n1235), .C2(new_n1236), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT60), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1205), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1255), .A2(KEYINPUT60), .A3(new_n1101), .A4(new_n1104), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1254), .A2(new_n1256), .A3(new_n1109), .A4(new_n721), .ZN(new_n1257));
  AND3_X1   g1057(.A1(new_n1257), .A2(G384), .A3(new_n1227), .ZN(new_n1258));
  AOI21_X1  g1058(.A(G384), .B1(new_n1257), .B2(new_n1227), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1245), .B1(new_n1252), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1247), .A2(G2897), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1263), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1257), .A2(new_n1227), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1240), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1257), .A2(G384), .A3(new_n1227), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1263), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1266), .A2(new_n1267), .A3(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1264), .A2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(KEYINPUT61), .B1(new_n1252), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(G375), .A2(G378), .ZN(new_n1272));
  AND3_X1   g1072(.A1(new_n1249), .A2(new_n1184), .A3(new_n1250), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1247), .B1(new_n1273), .B2(new_n1236), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1272), .A2(new_n1274), .A3(new_n1260), .A4(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1262), .A2(new_n1271), .A3(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1066), .B1(new_n979), .B2(new_n1005), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1239), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(G393), .A2(G396), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT125), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1280), .A2(KEYINPUT125), .A3(new_n1281), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1279), .A2(new_n1286), .A3(new_n1238), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1238), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1285), .B1(new_n1288), .B2(new_n1278), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1277), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1272), .A2(new_n1274), .A3(new_n1260), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT63), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT124), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1264), .A2(new_n1269), .A3(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1294), .B1(new_n1264), .B2(new_n1269), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  AOI22_X1  g1097(.A1(new_n1292), .A2(new_n1293), .B1(new_n1297), .B2(new_n1252), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1229), .A2(new_n1199), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1101), .B1(new_n1087), .B2(new_n1107), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1231), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1234), .A2(new_n721), .A3(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1236), .B1(new_n1302), .B2(new_n1186), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1249), .A2(new_n1184), .A3(new_n1250), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1248), .B1(new_n1304), .B2(G378), .ZN(new_n1305));
  NOR3_X1   g1105(.A1(new_n1303), .A2(new_n1305), .A3(new_n1261), .ZN(new_n1306));
  AOI21_X1  g1106(.A(KEYINPUT61), .B1(new_n1306), .B2(KEYINPUT63), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1298), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1291), .A2(new_n1309), .ZN(G405));
  NAND2_X1  g1110(.A1(new_n1272), .A2(new_n1237), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(new_n1260), .B(KEYINPUT127), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1311), .A2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1312), .A2(new_n1272), .A3(new_n1237), .ZN(new_n1315));
  AND3_X1   g1115(.A1(new_n1314), .A2(new_n1290), .A3(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1290), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1316), .A2(new_n1317), .ZN(G402));
endmodule


