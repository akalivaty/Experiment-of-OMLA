

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580;

  NOR2_X1 U324 ( .A1(n536), .A2(n416), .ZN(n564) );
  XOR2_X1 U325 ( .A(G78GAT), .B(G148GAT), .Z(n292) );
  XNOR2_X1 U326 ( .A(KEYINPUT113), .B(n408), .ZN(n293) );
  XNOR2_X1 U327 ( .A(n409), .B(KEYINPUT46), .ZN(n410) );
  XNOR2_X1 U328 ( .A(n403), .B(n402), .ZN(n404) );
  AND2_X1 U329 ( .A1(n293), .A2(n413), .ZN(n414) );
  XNOR2_X1 U330 ( .A(n405), .B(n404), .ZN(n569) );
  INV_X1 U331 ( .A(G190GAT), .ZN(n451) );
  XOR2_X1 U332 ( .A(n448), .B(n447), .Z(n520) );
  XNOR2_X1 U333 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U334 ( .A(n454), .B(n453), .ZN(G1351GAT) );
  XOR2_X1 U335 ( .A(KEYINPUT70), .B(KEYINPUT8), .Z(n295) );
  XNOR2_X1 U336 ( .A(G50GAT), .B(G43GAT), .ZN(n294) );
  XNOR2_X1 U337 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U338 ( .A(KEYINPUT7), .B(n296), .Z(n363) );
  XOR2_X1 U339 ( .A(G29GAT), .B(G134GAT), .Z(n326) );
  XOR2_X1 U340 ( .A(KEYINPUT79), .B(KEYINPUT78), .Z(n298) );
  XNOR2_X1 U341 ( .A(G218GAT), .B(KEYINPUT80), .ZN(n297) );
  XNOR2_X1 U342 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U343 ( .A(n326), .B(n299), .Z(n301) );
  NAND2_X1 U344 ( .A1(G232GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U345 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U346 ( .A(n363), .B(n302), .ZN(n314) );
  XOR2_X1 U347 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n304) );
  XNOR2_X1 U348 ( .A(G106GAT), .B(G92GAT), .ZN(n303) );
  XNOR2_X1 U349 ( .A(n304), .B(n303), .ZN(n308) );
  XOR2_X1 U350 ( .A(KEYINPUT11), .B(KEYINPUT64), .Z(n306) );
  XNOR2_X1 U351 ( .A(G162GAT), .B(KEYINPUT66), .ZN(n305) );
  XNOR2_X1 U352 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U353 ( .A(n308), .B(n307), .Z(n312) );
  XNOR2_X1 U354 ( .A(G36GAT), .B(G190GAT), .ZN(n309) );
  XNOR2_X1 U355 ( .A(n309), .B(KEYINPUT81), .ZN(n341) );
  XNOR2_X1 U356 ( .A(G99GAT), .B(G85GAT), .ZN(n310) );
  XNOR2_X1 U357 ( .A(n310), .B(KEYINPUT75), .ZN(n390) );
  XNOR2_X1 U358 ( .A(n341), .B(n390), .ZN(n311) );
  XNOR2_X1 U359 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U360 ( .A(n314), .B(n313), .ZN(n450) );
  XOR2_X1 U361 ( .A(KEYINPUT2), .B(KEYINPUT91), .Z(n316) );
  XNOR2_X1 U362 ( .A(G141GAT), .B(G155GAT), .ZN(n315) );
  XNOR2_X1 U363 ( .A(n316), .B(n315), .ZN(n318) );
  XOR2_X1 U364 ( .A(G162GAT), .B(KEYINPUT3), .Z(n317) );
  XOR2_X1 U365 ( .A(n318), .B(n317), .Z(n422) );
  XOR2_X1 U366 ( .A(KEYINPUT4), .B(KEYINPUT1), .Z(n320) );
  XNOR2_X1 U367 ( .A(KEYINPUT95), .B(KEYINPUT6), .ZN(n319) );
  XNOR2_X1 U368 ( .A(n320), .B(n319), .ZN(n333) );
  XOR2_X1 U369 ( .A(KEYINPUT5), .B(KEYINPUT94), .Z(n322) );
  XOR2_X1 U370 ( .A(G120GAT), .B(G57GAT), .Z(n401) );
  XOR2_X1 U371 ( .A(G1GAT), .B(G127GAT), .Z(n384) );
  XNOR2_X1 U372 ( .A(n401), .B(n384), .ZN(n321) );
  XNOR2_X1 U373 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U374 ( .A(n323), .B(G85GAT), .Z(n331) );
  XOR2_X1 U375 ( .A(KEYINPUT88), .B(KEYINPUT0), .Z(n325) );
  XNOR2_X1 U376 ( .A(G113GAT), .B(KEYINPUT87), .ZN(n324) );
  XNOR2_X1 U377 ( .A(n325), .B(n324), .ZN(n432) );
  XOR2_X1 U378 ( .A(n326), .B(n432), .Z(n328) );
  NAND2_X1 U379 ( .A1(G225GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U380 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U381 ( .A(G148GAT), .B(n329), .ZN(n330) );
  XNOR2_X1 U382 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U383 ( .A(n333), .B(n332), .Z(n334) );
  XOR2_X1 U384 ( .A(n422), .B(n334), .Z(n463) );
  XNOR2_X1 U385 ( .A(KEYINPUT96), .B(n463), .ZN(n536) );
  XOR2_X1 U386 ( .A(KEYINPUT21), .B(G218GAT), .Z(n336) );
  XNOR2_X1 U387 ( .A(KEYINPUT90), .B(G211GAT), .ZN(n335) );
  XNOR2_X1 U388 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U389 ( .A(G197GAT), .B(n337), .Z(n418) );
  XOR2_X1 U390 ( .A(G92GAT), .B(G64GAT), .Z(n339) );
  XNOR2_X1 U391 ( .A(G176GAT), .B(KEYINPUT76), .ZN(n338) );
  XNOR2_X1 U392 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U393 ( .A(G204GAT), .B(n340), .Z(n403) );
  XOR2_X1 U394 ( .A(n341), .B(KEYINPUT99), .Z(n343) );
  NAND2_X1 U395 ( .A1(G226GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U396 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U397 ( .A(n403), .B(n344), .ZN(n350) );
  XOR2_X1 U398 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n348) );
  XOR2_X1 U399 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n346) );
  XNOR2_X1 U400 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n345) );
  XNOR2_X1 U401 ( .A(n346), .B(n345), .ZN(n437) );
  XOR2_X1 U402 ( .A(G8GAT), .B(G183GAT), .Z(n377) );
  XNOR2_X1 U403 ( .A(n437), .B(n377), .ZN(n347) );
  XNOR2_X1 U404 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U405 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U406 ( .A(n418), .B(n351), .ZN(n456) );
  XOR2_X1 U407 ( .A(KEYINPUT67), .B(G1GAT), .Z(n353) );
  XNOR2_X1 U408 ( .A(G8GAT), .B(KEYINPUT29), .ZN(n352) );
  XNOR2_X1 U409 ( .A(n353), .B(n352), .ZN(n367) );
  XOR2_X1 U410 ( .A(G197GAT), .B(G141GAT), .Z(n355) );
  XNOR2_X1 U411 ( .A(G29GAT), .B(G36GAT), .ZN(n354) );
  XNOR2_X1 U412 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U413 ( .A(n356), .B(G113GAT), .Z(n358) );
  XOR2_X1 U414 ( .A(G15GAT), .B(G22GAT), .Z(n385) );
  XNOR2_X1 U415 ( .A(G169GAT), .B(n385), .ZN(n357) );
  XNOR2_X1 U416 ( .A(n358), .B(n357), .ZN(n362) );
  XOR2_X1 U417 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n360) );
  NAND2_X1 U418 ( .A1(G229GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U419 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U420 ( .A(n362), .B(n361), .Z(n365) );
  XNOR2_X1 U421 ( .A(n363), .B(KEYINPUT69), .ZN(n364) );
  XNOR2_X1 U422 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U423 ( .A(n367), .B(n366), .ZN(n565) );
  INV_X1 U424 ( .A(n565), .ZN(n540) );
  XOR2_X1 U425 ( .A(G71GAT), .B(KEYINPUT13), .Z(n400) );
  XOR2_X1 U426 ( .A(n400), .B(KEYINPUT12), .Z(n369) );
  NAND2_X1 U427 ( .A1(G231GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U428 ( .A(n369), .B(n368), .ZN(n373) );
  XOR2_X1 U429 ( .A(KEYINPUT14), .B(KEYINPUT82), .Z(n371) );
  XNOR2_X1 U430 ( .A(KEYINPUT86), .B(KEYINPUT15), .ZN(n370) );
  XNOR2_X1 U431 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U432 ( .A(n373), .B(n372), .Z(n379) );
  XOR2_X1 U433 ( .A(KEYINPUT83), .B(KEYINPUT84), .Z(n375) );
  XNOR2_X1 U434 ( .A(G57GAT), .B(KEYINPUT85), .ZN(n374) );
  XNOR2_X1 U435 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U436 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U437 ( .A(n379), .B(n378), .ZN(n383) );
  XOR2_X1 U438 ( .A(G64GAT), .B(G78GAT), .Z(n381) );
  XNOR2_X1 U439 ( .A(G155GAT), .B(G211GAT), .ZN(n380) );
  XNOR2_X1 U440 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U441 ( .A(n383), .B(n382), .Z(n387) );
  XNOR2_X1 U442 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U443 ( .A(n387), .B(n386), .ZN(n573) );
  XNOR2_X1 U444 ( .A(n450), .B(KEYINPUT36), .ZN(n577) );
  NOR2_X1 U445 ( .A1(n573), .A2(n577), .ZN(n388) );
  XNOR2_X1 U446 ( .A(n388), .B(KEYINPUT45), .ZN(n406) );
  XNOR2_X1 U447 ( .A(G106GAT), .B(KEYINPUT74), .ZN(n389) );
  XNOR2_X1 U448 ( .A(n292), .B(n389), .ZN(n417) );
  XNOR2_X1 U449 ( .A(n417), .B(n390), .ZN(n395) );
  XOR2_X1 U450 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n392) );
  NAND2_X1 U451 ( .A1(G230GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U452 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U453 ( .A(n393), .B(KEYINPUT71), .Z(n394) );
  XNOR2_X1 U454 ( .A(n395), .B(n394), .ZN(n399) );
  XOR2_X1 U455 ( .A(KEYINPUT77), .B(KEYINPUT72), .Z(n397) );
  XNOR2_X1 U456 ( .A(KEYINPUT31), .B(KEYINPUT73), .ZN(n396) );
  XNOR2_X1 U457 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U458 ( .A(n399), .B(n398), .Z(n405) );
  XNOR2_X1 U459 ( .A(n401), .B(n400), .ZN(n402) );
  NAND2_X1 U460 ( .A1(n406), .A2(n569), .ZN(n407) );
  NOR2_X1 U461 ( .A1(n540), .A2(n407), .ZN(n408) );
  INV_X1 U462 ( .A(n450), .ZN(n548) );
  XNOR2_X1 U463 ( .A(KEYINPUT41), .B(n569), .ZN(n553) );
  NAND2_X1 U464 ( .A1(n540), .A2(n553), .ZN(n409) );
  NAND2_X1 U465 ( .A1(n410), .A2(n573), .ZN(n411) );
  NOR2_X1 U466 ( .A1(n548), .A2(n411), .ZN(n412) );
  XNOR2_X1 U467 ( .A(n412), .B(KEYINPUT47), .ZN(n413) );
  XNOR2_X1 U468 ( .A(KEYINPUT48), .B(n414), .ZN(n539) );
  NOR2_X1 U469 ( .A1(n456), .A2(n539), .ZN(n415) );
  XOR2_X1 U470 ( .A(KEYINPUT54), .B(n415), .Z(n416) );
  XOR2_X1 U471 ( .A(G204GAT), .B(KEYINPUT93), .Z(n420) );
  XNOR2_X1 U472 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U473 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U474 ( .A(n422), .B(n421), .ZN(n430) );
  NAND2_X1 U475 ( .A1(G228GAT), .A2(G233GAT), .ZN(n428) );
  XOR2_X1 U476 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n424) );
  XNOR2_X1 U477 ( .A(KEYINPUT23), .B(KEYINPUT92), .ZN(n423) );
  XNOR2_X1 U478 ( .A(n424), .B(n423), .ZN(n426) );
  XOR2_X1 U479 ( .A(G50GAT), .B(G22GAT), .Z(n425) );
  XNOR2_X1 U480 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U481 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U482 ( .A(n430), .B(n429), .ZN(n464) );
  NAND2_X1 U483 ( .A1(n564), .A2(n464), .ZN(n431) );
  XNOR2_X1 U484 ( .A(KEYINPUT55), .B(n431), .ZN(n449) );
  XOR2_X1 U485 ( .A(n432), .B(G15GAT), .Z(n434) );
  NAND2_X1 U486 ( .A1(G227GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U487 ( .A(n434), .B(n433), .ZN(n448) );
  XOR2_X1 U488 ( .A(G190GAT), .B(G134GAT), .Z(n436) );
  XNOR2_X1 U489 ( .A(G43GAT), .B(G99GAT), .ZN(n435) );
  XNOR2_X1 U490 ( .A(n436), .B(n435), .ZN(n438) );
  XOR2_X1 U491 ( .A(n438), .B(n437), .Z(n446) );
  XOR2_X1 U492 ( .A(G127GAT), .B(G120GAT), .Z(n440) );
  XNOR2_X1 U493 ( .A(G71GAT), .B(KEYINPUT20), .ZN(n439) );
  XNOR2_X1 U494 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U495 ( .A(G176GAT), .B(G183GAT), .Z(n442) );
  XNOR2_X1 U496 ( .A(KEYINPUT89), .B(KEYINPUT65), .ZN(n441) );
  XNOR2_X1 U497 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U498 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U499 ( .A(n446), .B(n445), .ZN(n447) );
  NAND2_X1 U500 ( .A1(n449), .A2(n520), .ZN(n560) );
  NOR2_X1 U501 ( .A1(n450), .A2(n560), .ZN(n454) );
  XNOR2_X1 U502 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n452) );
  NAND2_X1 U503 ( .A1(n540), .A2(n569), .ZN(n487) );
  XNOR2_X1 U504 ( .A(KEYINPUT27), .B(n456), .ZN(n465) );
  NOR2_X1 U505 ( .A1(n520), .A2(n464), .ZN(n455) );
  XOR2_X1 U506 ( .A(KEYINPUT26), .B(n455), .Z(n562) );
  NOR2_X1 U507 ( .A1(n465), .A2(n562), .ZN(n537) );
  INV_X1 U508 ( .A(n456), .ZN(n511) );
  AND2_X1 U509 ( .A1(n520), .A2(n511), .ZN(n457) );
  XOR2_X1 U510 ( .A(KEYINPUT100), .B(n457), .Z(n458) );
  NAND2_X1 U511 ( .A1(n464), .A2(n458), .ZN(n459) );
  XNOR2_X1 U512 ( .A(n459), .B(KEYINPUT101), .ZN(n460) );
  XOR2_X1 U513 ( .A(KEYINPUT25), .B(n460), .Z(n461) );
  NOR2_X1 U514 ( .A1(n537), .A2(n461), .ZN(n462) );
  NOR2_X1 U515 ( .A1(n463), .A2(n462), .ZN(n468) );
  XOR2_X1 U516 ( .A(KEYINPUT28), .B(n464), .Z(n514) );
  NOR2_X1 U517 ( .A1(n465), .A2(n514), .ZN(n466) );
  NAND2_X1 U518 ( .A1(n466), .A2(n536), .ZN(n519) );
  NOR2_X1 U519 ( .A1(n520), .A2(n519), .ZN(n467) );
  NOR2_X1 U520 ( .A1(n468), .A2(n467), .ZN(n469) );
  XNOR2_X1 U521 ( .A(KEYINPUT102), .B(n469), .ZN(n484) );
  NOR2_X1 U522 ( .A1(n573), .A2(n548), .ZN(n470) );
  XOR2_X1 U523 ( .A(KEYINPUT16), .B(n470), .Z(n471) );
  NOR2_X1 U524 ( .A1(n484), .A2(n471), .ZN(n472) );
  XNOR2_X1 U525 ( .A(KEYINPUT103), .B(n472), .ZN(n497) );
  NOR2_X1 U526 ( .A1(n487), .A2(n497), .ZN(n473) );
  XNOR2_X1 U527 ( .A(n473), .B(KEYINPUT104), .ZN(n482) );
  NAND2_X1 U528 ( .A1(n536), .A2(n482), .ZN(n475) );
  XOR2_X1 U529 ( .A(KEYINPUT34), .B(KEYINPUT105), .Z(n474) );
  XNOR2_X1 U530 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U531 ( .A(G1GAT), .B(n476), .ZN(G1324GAT) );
  NAND2_X1 U532 ( .A1(n511), .A2(n482), .ZN(n477) );
  XNOR2_X1 U533 ( .A(G8GAT), .B(n477), .ZN(G1325GAT) );
  XOR2_X1 U534 ( .A(KEYINPUT35), .B(KEYINPUT107), .Z(n479) );
  NAND2_X1 U535 ( .A1(n520), .A2(n482), .ZN(n478) );
  XNOR2_X1 U536 ( .A(n479), .B(n478), .ZN(n481) );
  XOR2_X1 U537 ( .A(G15GAT), .B(KEYINPUT106), .Z(n480) );
  XNOR2_X1 U538 ( .A(n481), .B(n480), .ZN(G1326GAT) );
  NAND2_X1 U539 ( .A1(n482), .A2(n514), .ZN(n483) );
  XNOR2_X1 U540 ( .A(n483), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U541 ( .A(G29GAT), .B(KEYINPUT39), .Z(n490) );
  NOR2_X1 U542 ( .A1(n577), .A2(n484), .ZN(n485) );
  NAND2_X1 U543 ( .A1(n485), .A2(n573), .ZN(n486) );
  XOR2_X1 U544 ( .A(KEYINPUT37), .B(n486), .Z(n509) );
  NOR2_X1 U545 ( .A1(n509), .A2(n487), .ZN(n488) );
  XNOR2_X1 U546 ( .A(n488), .B(KEYINPUT38), .ZN(n495) );
  NAND2_X1 U547 ( .A1(n495), .A2(n536), .ZN(n489) );
  XNOR2_X1 U548 ( .A(n490), .B(n489), .ZN(G1328GAT) );
  NAND2_X1 U549 ( .A1(n495), .A2(n511), .ZN(n491) );
  XNOR2_X1 U550 ( .A(n491), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U551 ( .A(KEYINPUT40), .B(KEYINPUT108), .Z(n493) );
  NAND2_X1 U552 ( .A1(n520), .A2(n495), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U554 ( .A(G43GAT), .B(n494), .Z(G1330GAT) );
  NAND2_X1 U555 ( .A1(n495), .A2(n514), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n496), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT42), .B(KEYINPUT109), .Z(n499) );
  NAND2_X1 U558 ( .A1(n553), .A2(n565), .ZN(n508) );
  NOR2_X1 U559 ( .A1(n497), .A2(n508), .ZN(n504) );
  NAND2_X1 U560 ( .A1(n504), .A2(n536), .ZN(n498) );
  XNOR2_X1 U561 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U562 ( .A(G57GAT), .B(n500), .ZN(G1332GAT) );
  NAND2_X1 U563 ( .A1(n504), .A2(n511), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n501), .B(KEYINPUT110), .ZN(n502) );
  XNOR2_X1 U565 ( .A(G64GAT), .B(n502), .ZN(G1333GAT) );
  NAND2_X1 U566 ( .A1(n504), .A2(n520), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n503), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT43), .B(KEYINPUT111), .Z(n506) );
  NAND2_X1 U569 ( .A1(n504), .A2(n514), .ZN(n505) );
  XNOR2_X1 U570 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X1 U571 ( .A(G78GAT), .B(n507), .Z(G1335GAT) );
  NOR2_X1 U572 ( .A1(n509), .A2(n508), .ZN(n515) );
  NAND2_X1 U573 ( .A1(n515), .A2(n536), .ZN(n510) );
  XNOR2_X1 U574 ( .A(G85GAT), .B(n510), .ZN(G1336GAT) );
  NAND2_X1 U575 ( .A1(n515), .A2(n511), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n512), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U577 ( .A1(n515), .A2(n520), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n513), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT112), .B(KEYINPUT44), .Z(n517) );
  NAND2_X1 U580 ( .A1(n515), .A2(n514), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n517), .B(n516), .ZN(n518) );
  XOR2_X1 U582 ( .A(G106GAT), .B(n518), .Z(G1339GAT) );
  XOR2_X1 U583 ( .A(G113GAT), .B(KEYINPUT115), .Z(n524) );
  NOR2_X1 U584 ( .A1(n539), .A2(n519), .ZN(n521) );
  NAND2_X1 U585 ( .A1(n521), .A2(n520), .ZN(n522) );
  XOR2_X1 U586 ( .A(KEYINPUT114), .B(n522), .Z(n532) );
  NAND2_X1 U587 ( .A1(n540), .A2(n532), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n524), .B(n523), .ZN(G1340GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n526) );
  NAND2_X1 U590 ( .A1(n553), .A2(n532), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U592 ( .A(G120GAT), .B(n527), .ZN(G1341GAT) );
  INV_X1 U593 ( .A(n573), .ZN(n545) );
  NAND2_X1 U594 ( .A1(n532), .A2(n545), .ZN(n528) );
  XNOR2_X1 U595 ( .A(n528), .B(KEYINPUT50), .ZN(n529) );
  XNOR2_X1 U596 ( .A(G127GAT), .B(n529), .ZN(G1342GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n531) );
  XNOR2_X1 U598 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n530) );
  XNOR2_X1 U599 ( .A(n531), .B(n530), .ZN(n535) );
  NAND2_X1 U600 ( .A1(n532), .A2(n548), .ZN(n533) );
  XNOR2_X1 U601 ( .A(n533), .B(KEYINPUT117), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(G1343GAT) );
  NAND2_X1 U603 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U604 ( .A1(n539), .A2(n538), .ZN(n547) );
  NAND2_X1 U605 ( .A1(n547), .A2(n540), .ZN(n541) );
  XNOR2_X1 U606 ( .A(n541), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n543) );
  NAND2_X1 U608 ( .A1(n547), .A2(n553), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(n544), .ZN(G1345GAT) );
  NAND2_X1 U611 ( .A1(n545), .A2(n547), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n546), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U613 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n549), .B(KEYINPUT120), .ZN(n550) );
  XNOR2_X1 U615 ( .A(G162GAT), .B(n550), .ZN(G1347GAT) );
  NOR2_X1 U616 ( .A1(n565), .A2(n560), .ZN(n552) );
  XNOR2_X1 U617 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(G1348GAT) );
  INV_X1 U619 ( .A(n553), .ZN(n554) );
  NOR2_X1 U620 ( .A1(n554), .A2(n560), .ZN(n559) );
  XOR2_X1 U621 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n556) );
  XNOR2_X1 U622 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U624 ( .A(KEYINPUT56), .B(n557), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(G1349GAT) );
  NOR2_X1 U626 ( .A1(n573), .A2(n560), .ZN(n561) );
  XOR2_X1 U627 ( .A(G183GAT), .B(n561), .Z(G1350GAT) );
  INV_X1 U628 ( .A(n562), .ZN(n563) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n576) );
  NOR2_X1 U630 ( .A1(n565), .A2(n576), .ZN(n567) );
  XNOR2_X1 U631 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(n568), .ZN(G1352GAT) );
  NOR2_X1 U634 ( .A1(n569), .A2(n576), .ZN(n571) );
  XNOR2_X1 U635 ( .A(KEYINPUT61), .B(KEYINPUT125), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XOR2_X1 U637 ( .A(G204GAT), .B(n572), .Z(G1353GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n576), .ZN(n574) );
  XOR2_X1 U639 ( .A(KEYINPUT126), .B(n574), .Z(n575) );
  XNOR2_X1 U640 ( .A(G211GAT), .B(n575), .ZN(G1354GAT) );
  NOR2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n579) );
  XNOR2_X1 U642 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(n580), .ZN(G1355GAT) );
endmodule

