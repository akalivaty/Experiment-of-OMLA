//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 0 1 1 0 0 1 0 1 1 1 1 1 0 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 1 1 1 0 0 1 1 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n445, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n566, new_n567, new_n569, new_n570, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n630,
    new_n631, new_n634, new_n636, new_n637, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n847, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1200;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT64), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n467), .A3(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(KEYINPUT66), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n470), .A2(new_n473), .A3(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G101), .ZN(new_n476));
  NOR3_X1   g051(.A1(new_n476), .A2(new_n464), .A3(G2105), .ZN(new_n477));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n479), .A2(new_n464), .A3(KEYINPUT3), .ZN(new_n480));
  AOI21_X1  g055(.A(KEYINPUT67), .B1(new_n466), .B2(G2104), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n466), .A2(G2104), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n478), .B(new_n480), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n477), .B1(new_n484), .B2(G137), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n475), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G160));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n478), .ZN(new_n489));
  INV_X1    g064(.A(G136), .ZN(new_n490));
  INV_X1    g065(.A(G124), .ZN(new_n491));
  OAI211_X1 g066(.A(G2105), .B(new_n480), .C1(new_n481), .C2(new_n482), .ZN(new_n492));
  OAI221_X1 g067(.A(new_n489), .B1(new_n483), .B2(new_n490), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n494));
  XNOR2_X1  g069(.A(new_n493), .B(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G162));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  OAI21_X1  g072(.A(KEYINPUT4), .B1(new_n483), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n465), .A2(new_n467), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(new_n478), .A3(G138), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G126), .ZN(new_n505));
  NOR2_X1   g080(.A1(G102), .A2(G2105), .ZN(new_n506));
  OAI21_X1  g081(.A(G2104), .B1(new_n478), .B2(G114), .ZN(new_n507));
  OAI22_X1  g082(.A1(new_n492), .A2(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT69), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n504), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n479), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(new_n465), .ZN(new_n513));
  NAND4_X1  g088(.A1(new_n513), .A2(G138), .A3(new_n478), .A4(new_n480), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n502), .B1(new_n514), .B2(KEYINPUT4), .ZN(new_n515));
  OAI21_X1  g090(.A(KEYINPUT69), .B1(new_n515), .B2(new_n508), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n511), .A2(new_n516), .ZN(G164));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(KEYINPUT5), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT5), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G62), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n518), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT70), .B(G651), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n526), .A2(KEYINPUT6), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(KEYINPUT71), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT6), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G651), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT71), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n526), .A2(new_n533), .A3(KEYINPUT6), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n530), .A2(G543), .A3(new_n532), .A4(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(G50), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n528), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n520), .A2(new_n522), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n530), .A2(new_n538), .A3(new_n532), .A4(new_n534), .ZN(new_n539));
  XOR2_X1   g114(.A(KEYINPUT72), .B(G88), .Z(new_n540));
  NOR2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n537), .A2(new_n541), .ZN(G166));
  INV_X1    g117(.A(new_n539), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n543), .A2(G89), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n538), .A2(G63), .A3(G651), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT73), .ZN(new_n546));
  INV_X1    g121(.A(G51), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n547), .B2(new_n535), .ZN(new_n548));
  NAND3_X1  g123(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n549));
  XOR2_X1   g124(.A(new_n549), .B(KEYINPUT7), .Z(new_n550));
  NOR3_X1   g125(.A1(new_n544), .A2(new_n548), .A3(new_n550), .ZN(G168));
  INV_X1    g126(.A(G52), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n538), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n535), .A2(new_n552), .B1(new_n526), .B2(new_n553), .ZN(new_n554));
  XNOR2_X1  g129(.A(KEYINPUT74), .B(G90), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n539), .A2(new_n555), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n554), .A2(new_n556), .ZN(G301));
  INV_X1    g132(.A(G301), .ZN(G171));
  INV_X1    g133(.A(G43), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n538), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n560));
  OAI22_X1  g135(.A1(new_n535), .A2(new_n559), .B1(new_n526), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(G81), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n539), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  AND3_X1   g140(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G36), .ZN(new_n567));
  XOR2_X1   g142(.A(new_n567), .B(KEYINPUT75), .Z(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n566), .A2(new_n570), .ZN(G188));
  INV_X1    g146(.A(new_n535), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n572), .A2(KEYINPUT9), .A3(G53), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n523), .B(KEYINPUT76), .ZN(new_n574));
  INV_X1    g149(.A(G65), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AND2_X1   g151(.A1(G78), .A2(G543), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n543), .A2(G91), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT9), .ZN(new_n580));
  INV_X1    g155(.A(G53), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n535), .B2(new_n581), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n573), .A2(new_n578), .A3(new_n579), .A4(new_n582), .ZN(G299));
  INV_X1    g158(.A(G168), .ZN(G286));
  INV_X1    g159(.A(G166), .ZN(G303));
  NAND2_X1  g160(.A1(new_n572), .A2(G49), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n543), .A2(G87), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n538), .B2(G74), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n586), .A2(new_n587), .A3(KEYINPUT77), .A4(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT77), .ZN(new_n590));
  INV_X1    g165(.A(G87), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n588), .B1(new_n539), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(G49), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n535), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n590), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n589), .A2(new_n595), .ZN(G288));
  NAND3_X1  g171(.A1(new_n538), .A2(KEYINPUT78), .A3(G61), .ZN(new_n597));
  NAND2_X1  g172(.A1(G73), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n599));
  INV_X1    g174(.A(G61), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n523), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n597), .A2(new_n598), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(new_n527), .ZN(new_n603));
  INV_X1    g178(.A(G86), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(new_n539), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G48), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n535), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n606), .A2(new_n609), .ZN(G305));
  NAND2_X1  g185(.A1(new_n543), .A2(G85), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n572), .A2(G47), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n538), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n613));
  OAI211_X1 g188(.A(new_n611), .B(new_n612), .C1(new_n526), .C2(new_n613), .ZN(G290));
  NAND2_X1  g189(.A1(G301), .A2(G868), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n543), .A2(KEYINPUT10), .A3(G92), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT10), .ZN(new_n617));
  INV_X1    g192(.A(G92), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n539), .B2(new_n618), .ZN(new_n619));
  AOI22_X1  g194(.A1(new_n616), .A2(new_n619), .B1(G54), .B2(new_n572), .ZN(new_n620));
  INV_X1    g195(.A(G66), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n574), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(G79), .A2(G543), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT79), .Z(new_n624));
  OAI21_X1  g199(.A(G651), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n615), .B1(new_n627), .B2(G868), .ZN(G284));
  OAI21_X1  g203(.A(new_n615), .B1(new_n627), .B2(G868), .ZN(G321));
  INV_X1    g204(.A(G868), .ZN(new_n630));
  NAND2_X1  g205(.A1(G299), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(G168), .B2(new_n630), .ZN(G297));
  OAI21_X1  g207(.A(new_n631), .B1(G168), .B2(new_n630), .ZN(G280));
  INV_X1    g208(.A(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n627), .B1(new_n634), .B2(G860), .ZN(G148));
  NAND2_X1  g210(.A1(new_n627), .A2(new_n634), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G868), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(G868), .B2(new_n564), .ZN(G323));
  XNOR2_X1  g213(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g214(.A1(new_n484), .A2(G135), .ZN(new_n640));
  OR2_X1    g215(.A1(G99), .A2(G2105), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n641), .B(G2104), .C1(G111), .C2(new_n478), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(new_n492), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n643), .B1(G123), .B2(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2096), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n478), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT12), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2100), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT80), .B(KEYINPUT13), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n646), .A2(new_n651), .ZN(G156));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2438), .ZN(new_n654));
  XOR2_X1   g229(.A(G2427), .B(G2430), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT81), .B(KEYINPUT14), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT82), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  XOR2_X1   g235(.A(G1341), .B(G1348), .Z(new_n661));
  XNOR2_X1  g236(.A(G2451), .B(G2454), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2443), .B(G2446), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n660), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(G14), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(G401));
  XOR2_X1   g243(.A(G2067), .B(G2678), .Z(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G2084), .B(G2090), .Z(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g247(.A1(new_n672), .A2(KEYINPUT17), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n670), .A2(new_n671), .ZN(new_n674));
  AOI21_X1  g249(.A(KEYINPUT18), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2072), .B(G2078), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT83), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(KEYINPUT18), .B2(new_n672), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n675), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G2096), .B(G2100), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(G227));
  XNOR2_X1  g256(.A(G1981), .B(G1986), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1971), .B(G1976), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT84), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT19), .ZN(new_n686));
  XOR2_X1   g261(.A(G1956), .B(G2474), .Z(new_n687));
  XOR2_X1   g262(.A(G1961), .B(G1966), .Z(new_n688));
  AND2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT86), .Z(new_n691));
  XOR2_X1   g266(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n692));
  NOR2_X1   g267(.A1(new_n687), .A2(new_n688), .ZN(new_n693));
  AOI22_X1  g268(.A1(new_n691), .A2(new_n692), .B1(new_n686), .B2(new_n693), .ZN(new_n694));
  OR3_X1    g269(.A1(new_n686), .A2(new_n689), .A3(new_n693), .ZN(new_n695));
  OAI211_X1 g270(.A(new_n694), .B(new_n695), .C1(new_n691), .C2(new_n692), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT87), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n696), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(G1991), .B(G1996), .Z(new_n700));
  AND2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n699), .A2(new_n700), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n683), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n699), .A2(new_n700), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n699), .A2(new_n700), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n704), .A2(new_n682), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n703), .A2(new_n706), .ZN(G229));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G22), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G166), .B2(new_n708), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(G1971), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n708), .A2(G23), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT88), .ZN(new_n713));
  NAND4_X1  g288(.A1(new_n586), .A2(new_n587), .A3(new_n713), .A4(new_n588), .ZN(new_n714));
  OAI21_X1  g289(.A(KEYINPUT88), .B1(new_n592), .B2(new_n594), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n712), .B1(new_n716), .B2(new_n708), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT89), .B(KEYINPUT33), .ZN(new_n718));
  INV_X1    g293(.A(G1976), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n711), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n708), .A2(G6), .ZN(new_n722));
  INV_X1    g297(.A(G305), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n723), .B2(new_n708), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT32), .B(G1981), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n721), .B(new_n726), .C1(new_n720), .C2(new_n717), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n727), .A2(KEYINPUT34), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n708), .A2(G24), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G290), .B2(G16), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(G1986), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n727), .A2(KEYINPUT34), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n644), .A2(G119), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n484), .A2(G131), .ZN(new_n735));
  NOR2_X1   g310(.A1(G95), .A2(G2105), .ZN(new_n736));
  OAI21_X1  g311(.A(G2104), .B1(new_n478), .B2(G107), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n734), .B(new_n735), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  MUX2_X1   g313(.A(G25), .B(new_n738), .S(G29), .Z(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT35), .B(G1991), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G1986), .B2(new_n731), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n728), .A2(new_n732), .A3(new_n733), .A4(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(KEYINPUT36), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n733), .A2(new_n742), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT36), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n745), .A2(new_n746), .A3(new_n732), .A4(new_n728), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT99), .ZN(new_n749));
  INV_X1    g324(.A(G29), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(G35), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G162), .B2(new_n750), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT98), .Z(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(KEYINPUT29), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n752), .B(KEYINPUT98), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT29), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G2090), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n749), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n708), .A2(G19), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n564), .B2(new_n708), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G1341), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n758), .B2(new_n759), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n754), .A2(new_n757), .A3(KEYINPUT99), .A4(G2090), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n486), .A2(G29), .ZN(new_n766));
  OR2_X1    g341(.A1(KEYINPUT24), .A2(G34), .ZN(new_n767));
  NAND2_X1  g342(.A1(KEYINPUT24), .A2(G34), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n767), .A2(new_n750), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n770), .A2(G2084), .ZN(new_n771));
  INV_X1    g346(.A(G2072), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n750), .A2(G33), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n484), .A2(G139), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n478), .A2(G103), .A3(G2104), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT25), .Z(new_n776));
  INV_X1    g351(.A(new_n499), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n777), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n774), .B(new_n776), .C1(new_n478), .C2(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n773), .B1(new_n779), .B2(G29), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n771), .B1(new_n772), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n645), .A2(G29), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT94), .ZN(new_n783));
  INV_X1    g358(.A(G28), .ZN(new_n784));
  NOR3_X1   g359(.A1(new_n784), .A2(KEYINPUT95), .A3(KEYINPUT30), .ZN(new_n785));
  OAI21_X1  g360(.A(KEYINPUT95), .B1(new_n784), .B2(KEYINPUT30), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(new_n750), .ZN(new_n787));
  AOI211_X1 g362(.A(new_n785), .B(new_n787), .C1(KEYINPUT30), .C2(new_n784), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT93), .B(KEYINPUT31), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G11), .ZN(new_n790));
  NOR4_X1   g365(.A1(new_n781), .A2(new_n783), .A3(new_n788), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n708), .A2(G21), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G168), .B2(new_n708), .ZN(new_n793));
  INV_X1    g368(.A(G1966), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(G129), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n492), .A2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT91), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n478), .A2(G105), .A3(G2104), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT92), .ZN(new_n801));
  NAND3_X1  g376(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT26), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(new_n484), .B2(G141), .ZN(new_n804));
  AND3_X1   g379(.A1(new_n799), .A2(new_n801), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n805), .A2(G29), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G29), .B2(G32), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT27), .B(G1996), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n791), .A2(new_n795), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n708), .A2(G4), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n627), .B2(new_n708), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT90), .B(G1348), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n780), .A2(new_n772), .ZN(new_n815));
  NOR3_X1   g390(.A1(new_n810), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n760), .A2(new_n764), .A3(new_n765), .A4(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(G2084), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n766), .A2(new_n818), .A3(new_n769), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n708), .A2(G5), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G171), .B2(new_n708), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT96), .ZN(new_n822));
  OAI221_X1 g397(.A(new_n819), .B1(new_n807), .B2(new_n808), .C1(new_n822), .C2(G1961), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT97), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(G1961), .ZN(new_n825));
  NOR2_X1   g400(.A1(G27), .A2(G29), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(G164), .B2(G29), .ZN(new_n827));
  INV_X1    g402(.A(G2078), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n708), .A2(G20), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT100), .Z(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT23), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(G299), .B2(G16), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(G1956), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n825), .A2(new_n829), .A3(new_n834), .ZN(new_n835));
  NOR3_X1   g410(.A1(new_n817), .A2(new_n824), .A3(new_n835), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n750), .A2(G26), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n644), .A2(G128), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n484), .A2(G140), .ZN(new_n839));
  NOR2_X1   g414(.A1(G104), .A2(G2105), .ZN(new_n840));
  OAI21_X1  g415(.A(G2104), .B1(new_n478), .B2(G116), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n838), .B(new_n839), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n837), .B1(new_n842), .B2(G29), .ZN(new_n843));
  MUX2_X1   g418(.A(new_n837), .B(new_n843), .S(KEYINPUT28), .Z(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(G2067), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n748), .A2(new_n836), .A3(new_n845), .ZN(G150));
  INV_X1    g421(.A(KEYINPUT101), .ZN(new_n847));
  NAND2_X1  g422(.A1(G150), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n748), .A2(new_n836), .A3(KEYINPUT101), .A4(new_n845), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(G311));
  AOI22_X1  g425(.A1(new_n538), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n851), .A2(new_n526), .ZN(new_n852));
  INV_X1    g427(.A(G55), .ZN(new_n853));
  INV_X1    g428(.A(G93), .ZN(new_n854));
  OAI221_X1 g429(.A(new_n852), .B1(new_n535), .B2(new_n853), .C1(new_n854), .C2(new_n539), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT102), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n543), .A2(G93), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n572), .A2(G55), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n858), .A2(new_n859), .A3(KEYINPUT102), .A4(new_n852), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(G860), .ZN(new_n863));
  XOR2_X1   g438(.A(KEYINPUT103), .B(KEYINPUT37), .Z(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n626), .A2(new_n634), .ZN(new_n866));
  XOR2_X1   g441(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n564), .B1(new_n857), .B2(new_n860), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n855), .A2(new_n564), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n868), .B(new_n872), .Z(new_n873));
  OAI21_X1  g448(.A(new_n865), .B1(new_n873), .B2(G860), .ZN(G145));
  NAND2_X1  g449(.A1(new_n644), .A2(G130), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n484), .A2(G142), .ZN(new_n876));
  NOR2_X1   g451(.A1(G106), .A2(G2105), .ZN(new_n877));
  OAI21_X1  g452(.A(G2104), .B1(new_n478), .B2(G118), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n875), .B(new_n876), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(new_n648), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT104), .ZN(new_n882));
  AOI211_X1 g457(.A(new_n882), .B(new_n502), .C1(new_n514), .C2(KEYINPUT4), .ZN(new_n883));
  AOI21_X1  g458(.A(KEYINPUT104), .B1(new_n498), .B2(new_n503), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n509), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n779), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n738), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n805), .B(new_n842), .ZN(new_n888));
  AND2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n887), .A2(new_n888), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n881), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n887), .A2(new_n888), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n887), .A2(new_n888), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n892), .A2(new_n880), .A3(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n891), .A2(new_n894), .A3(KEYINPUT105), .ZN(new_n895));
  XNOR2_X1  g470(.A(G160), .B(new_n645), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n891), .A2(new_n894), .A3(KEYINPUT105), .A4(new_n896), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(G162), .ZN(new_n901));
  INV_X1    g476(.A(G37), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n898), .A2(new_n495), .A3(new_n899), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g480(.A(G299), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n626), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n620), .A2(G299), .A3(new_n625), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(KEYINPUT41), .ZN(new_n911));
  AOI21_X1  g486(.A(KEYINPUT107), .B1(new_n626), .B2(new_n906), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n912), .B1(new_n909), .B2(KEYINPUT107), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n911), .B1(new_n913), .B2(KEYINPUT41), .ZN(new_n914));
  XOR2_X1   g489(.A(new_n872), .B(new_n636), .Z(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT108), .ZN(new_n917));
  XOR2_X1   g492(.A(new_n909), .B(KEYINPUT106), .Z(new_n918));
  OR2_X1    g493(.A1(new_n918), .A2(new_n915), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT108), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n914), .A2(new_n915), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n917), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT109), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n923), .A2(KEYINPUT42), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(G290), .B(G166), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n926), .A2(new_n723), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n723), .ZN(new_n928));
  OR3_X1    g503(.A1(new_n927), .A2(new_n928), .A3(new_n716), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n716), .B1(new_n927), .B2(new_n928), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n932), .B1(new_n923), .B2(KEYINPUT42), .ZN(new_n933));
  INV_X1    g508(.A(new_n924), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n917), .A2(new_n919), .A3(new_n934), .A4(new_n921), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n925), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n933), .B1(new_n925), .B2(new_n935), .ZN(new_n937));
  OAI21_X1  g512(.A(G868), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n938), .B1(G868), .B2(new_n861), .ZN(G295));
  OAI21_X1  g514(.A(new_n938), .B1(G868), .B2(new_n861), .ZN(G331));
  INV_X1    g515(.A(KEYINPUT111), .ZN(new_n941));
  XNOR2_X1  g516(.A(G301), .B(KEYINPUT110), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n564), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n861), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n945), .A2(G286), .A3(new_n870), .ZN(new_n946));
  OAI21_X1  g521(.A(G168), .B1(new_n869), .B2(new_n871), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n946), .A2(new_n943), .A3(new_n947), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(new_n910), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n950), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n952), .A2(new_n948), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n951), .B1(new_n953), .B2(new_n914), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n932), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT43), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n931), .B(new_n951), .C1(new_n953), .C2(new_n914), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n955), .A2(new_n956), .A3(new_n902), .A4(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT44), .ZN(new_n959));
  AOI21_X1  g534(.A(G37), .B1(new_n954), .B2(new_n932), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n918), .A2(new_n950), .A3(new_n949), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n913), .A2(KEYINPUT41), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n962), .B1(KEYINPUT41), .B2(new_n910), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n961), .B(new_n931), .C1(new_n953), .C2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n956), .B1(new_n960), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n941), .B1(new_n959), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n955), .A2(new_n902), .A3(new_n964), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n968), .A2(KEYINPUT111), .A3(KEYINPUT44), .A4(new_n958), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n956), .B1(new_n960), .B2(new_n957), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n971), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n970), .A2(new_n974), .ZN(G397));
  XOR2_X1   g550(.A(KEYINPUT112), .B(G1384), .Z(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT45), .B1(new_n885), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n473), .B1(new_n470), .B2(G2105), .ZN(new_n979));
  AOI211_X1 g554(.A(KEYINPUT66), .B(new_n478), .C1(new_n468), .C2(new_n469), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n485), .B(G40), .C1(new_n979), .C2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT113), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n475), .A2(KEYINPUT113), .A3(G40), .A4(new_n485), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n978), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n986), .A2(G1996), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n987), .B(KEYINPUT114), .ZN(new_n988));
  INV_X1    g563(.A(new_n986), .ZN(new_n989));
  XOR2_X1   g564(.A(new_n842), .B(G2067), .Z(new_n990));
  INV_X1    g565(.A(G1996), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n990), .B1(new_n805), .B2(new_n991), .ZN(new_n992));
  AOI22_X1  g567(.A1(new_n988), .A2(new_n805), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n738), .A2(new_n740), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n738), .A2(new_n740), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n989), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  XNOR2_X1  g572(.A(G290), .B(G1986), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n997), .B1(new_n989), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n504), .A2(new_n882), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n515), .A2(KEYINPUT104), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n508), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1000), .B1(new_n1003), .B2(new_n976), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n885), .A2(KEYINPUT45), .A3(new_n977), .ZN(new_n1005));
  AND4_X1   g580(.A1(KEYINPUT53), .A2(new_n471), .A3(G40), .A4(new_n828), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1004), .A2(new_n485), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT126), .ZN(new_n1008));
  INV_X1    g583(.A(new_n485), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n885), .A2(new_n977), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1009), .B1(new_n1010), .B2(new_n1000), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT126), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1011), .A2(new_n1012), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1008), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n1015));
  INV_X1    g590(.A(G1384), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n511), .A2(new_n516), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n1000), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1018), .A2(new_n1005), .A3(new_n985), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1015), .B1(new_n1019), .B2(G2078), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1014), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G1961), .ZN(new_n1022));
  AOI22_X1  g597(.A1(KEYINPUT50), .A2(new_n1017), .B1(new_n983), .B2(new_n984), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT50), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n885), .A2(new_n1024), .A3(new_n1016), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT122), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1017), .A2(KEYINPUT50), .ZN(new_n1027));
  AND4_X1   g602(.A1(KEYINPUT122), .A2(new_n1027), .A3(new_n1025), .A4(new_n985), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1022), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT125), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1027), .A2(new_n1025), .A3(new_n985), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT122), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1023), .A2(KEYINPUT122), .A3(new_n1025), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT125), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(new_n1036), .A3(new_n1022), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1021), .B1(new_n1030), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT127), .B1(new_n1038), .B2(G301), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n828), .A2(KEYINPUT53), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1000), .B1(new_n1003), .B2(G1384), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1041), .B(new_n985), .C1(new_n1000), .C2(new_n1017), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1029), .B(new_n1020), .C1(new_n1040), .C2(new_n1042), .ZN(new_n1043));
  OR2_X1    g618(.A1(new_n1043), .A2(G171), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1018), .A2(new_n1005), .A3(new_n985), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT53), .B1(new_n1045), .B2(new_n828), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1046), .B1(new_n1008), .B2(new_n1013), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1036), .B1(new_n1035), .B2(new_n1022), .ZN(new_n1048));
  AOI211_X1 g623(.A(KEYINPUT125), .B(G1961), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1047), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT127), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1050), .A2(new_n1051), .A3(G171), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1039), .A2(KEYINPUT54), .A3(new_n1044), .A4(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT51), .ZN(new_n1054));
  INV_X1    g629(.A(G8), .ZN(new_n1055));
  NOR2_X1   g630(.A1(G168), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1042), .A2(new_n1058), .A3(new_n794), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1058), .B1(new_n1042), .B2(new_n794), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1031), .A2(G2084), .ZN(new_n1061));
  NOR3_X1   g636(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1054), .B(new_n1057), .C1(new_n1062), .C2(new_n1055), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1042), .A2(new_n794), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT117), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1061), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1042), .A2(new_n1058), .A3(new_n794), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  OAI211_X1 g643(.A(KEYINPUT51), .B(G8), .C1(new_n1068), .C2(G286), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1063), .A2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1062), .A2(new_n1057), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1003), .A2(G1384), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1055), .B1(new_n1074), .B2(new_n985), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n716), .A2(G1976), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT52), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT49), .ZN(new_n1079));
  OAI21_X1  g654(.A(G1981), .B1(new_n605), .B2(new_n608), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n605), .A2(G1981), .A3(new_n608), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1079), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1082), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1084), .A2(new_n1080), .A3(KEYINPUT49), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1083), .A2(new_n1085), .A3(new_n1075), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT52), .B1(G288), .B2(new_n719), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1087), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1078), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(G8), .B1(new_n537), .B2(new_n541), .ZN(new_n1090));
  XNOR2_X1  g665(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n1090), .B(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G1971), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1019), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1023), .A2(new_n759), .A3(new_n1025), .ZN(new_n1095));
  AOI211_X1 g670(.A(new_n1055), .B(new_n1092), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1089), .A2(new_n1096), .ZN(new_n1097));
  OR2_X1    g672(.A1(new_n1017), .A2(KEYINPUT50), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT50), .B1(new_n1003), .B2(G1384), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1098), .A2(new_n1099), .A3(new_n759), .A4(new_n985), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1055), .B1(new_n1094), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1092), .ZN(new_n1102));
  OR3_X1    g677(.A1(new_n1101), .A2(KEYINPUT116), .A3(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(KEYINPUT116), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1097), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1047), .B(G301), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1043), .A2(G171), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT54), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1105), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1053), .A2(new_n1073), .A3(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(G299), .B(KEYINPUT57), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT56), .B(G2072), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1045), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1098), .A2(new_n1099), .A3(new_n985), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n1117));
  INV_X1    g692(.A(G1956), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1117), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1113), .B(new_n1115), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1121), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n1119), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1126), .A2(KEYINPUT120), .A3(new_n1113), .A4(new_n1115), .ZN(new_n1127));
  INV_X1    g702(.A(new_n813), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1035), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1074), .A2(new_n985), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1130), .A2(G2067), .ZN(new_n1131));
  OR2_X1    g706(.A1(new_n1131), .A2(KEYINPUT121), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(KEYINPUT121), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1129), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(new_n627), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1135), .A2(KEYINPUT123), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1115), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(new_n1112), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1138), .B1(new_n1135), .B2(KEYINPUT123), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1124), .B(new_n1127), .C1(new_n1136), .C2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1124), .A2(new_n1127), .A3(new_n1138), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT61), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  OR2_X1    g718(.A1(new_n627), .A2(KEYINPUT60), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1129), .A2(new_n1132), .A3(new_n1133), .A4(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n627), .A2(KEYINPUT60), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1145), .B(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1138), .A2(KEYINPUT61), .A3(new_n1122), .ZN(new_n1148));
  XOR2_X1   g723(.A(KEYINPUT124), .B(G1996), .Z(new_n1149));
  NAND2_X1  g724(.A1(new_n1045), .A2(new_n1149), .ZN(new_n1150));
  XOR2_X1   g725(.A(KEYINPUT58), .B(G1341), .Z(new_n1151));
  NAND2_X1  g726(.A1(new_n1130), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n944), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  XOR2_X1   g728(.A(new_n1153), .B(KEYINPUT59), .Z(new_n1154));
  NAND4_X1  g729(.A1(new_n1143), .A2(new_n1147), .A3(new_n1148), .A4(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1111), .B1(new_n1140), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT63), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1097), .A2(G8), .A3(G168), .A4(new_n1068), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1157), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT118), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(G8), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1157), .B1(new_n1163), .B2(new_n1092), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1161), .B1(new_n1158), .B2(new_n1165), .ZN(new_n1166));
  NOR4_X1   g741(.A1(new_n1062), .A2(new_n1089), .A3(new_n1096), .A4(new_n1055), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1167), .A2(KEYINPUT118), .A3(G168), .A4(new_n1164), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1160), .A2(new_n1166), .A3(new_n1168), .ZN(new_n1169));
  NOR3_X1   g744(.A1(new_n1089), .A2(new_n1163), .A3(new_n1092), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1086), .A2(new_n719), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1084), .B1(new_n1171), .B2(G288), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1170), .B1(new_n1075), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT62), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1070), .A2(new_n1174), .A3(new_n1072), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1105), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1107), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1071), .B1(new_n1063), .B2(new_n1069), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1178), .B1(new_n1179), .B2(new_n1174), .ZN(new_n1180));
  OAI211_X1 g755(.A(new_n1169), .B(new_n1173), .C1(new_n1177), .C2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n999), .B1(new_n1156), .B2(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n988), .B(KEYINPUT46), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n986), .B1(new_n805), .B2(new_n990), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n1185), .B(KEYINPUT47), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n842), .A2(G2067), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1187), .B1(new_n993), .B2(new_n994), .ZN(new_n1188));
  NOR3_X1   g763(.A1(new_n986), .A2(G1986), .A3(G290), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n1189), .B(KEYINPUT48), .ZN(new_n1190));
  OAI22_X1  g765(.A1(new_n1188), .A2(new_n986), .B1(new_n997), .B2(new_n1190), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n1186), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1182), .A2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  AND3_X1   g768(.A1(new_n703), .A2(new_n706), .A3(new_n667), .ZN(new_n1195));
  NAND2_X1  g769(.A1(new_n1195), .A2(new_n904), .ZN(new_n1196));
  NOR2_X1   g770(.A1(G227), .A2(new_n462), .ZN(new_n1197));
  OAI21_X1  g771(.A(new_n1197), .B1(new_n972), .B2(new_n973), .ZN(new_n1198));
  NOR2_X1   g772(.A1(new_n1196), .A2(new_n1198), .ZN(G308));
  OR2_X1    g773(.A1(new_n972), .A2(new_n973), .ZN(new_n1200));
  NAND4_X1  g774(.A1(new_n1200), .A2(new_n904), .A3(new_n1197), .A4(new_n1195), .ZN(G225));
endmodule


