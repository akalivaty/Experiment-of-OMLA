//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 0 0 0 0 0 0 0 1 1 0 1 0 0 0 0 0 0 0 0 1 1 0 1 0 0 0 1 1 0 0 1 0 1 1 1 0 1 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT73), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT73), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G953), .ZN(new_n193));
  AND2_X1   g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G227), .ZN(new_n195));
  XOR2_X1   g009(.A(G110), .B(G140), .Z(new_n196));
  XNOR2_X1  g010(.A(new_n195), .B(new_n196), .ZN(new_n197));
  OR2_X1    g011(.A1(KEYINPUT66), .A2(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(KEYINPUT66), .A2(G146), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(G143), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(G143), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(KEYINPUT1), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n200), .A2(new_n203), .A3(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT90), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n200), .A2(KEYINPUT90), .A3(new_n203), .A4(new_n205), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n200), .A2(new_n203), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(G146), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT1), .ZN(new_n213));
  OAI21_X1  g027(.A(G128), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n210), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n208), .A2(new_n209), .A3(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G104), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(G107), .ZN(new_n218));
  AND2_X1   g032(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n219));
  NOR2_X1   g033(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT87), .ZN(new_n222));
  INV_X1    g036(.A(G107), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n222), .B1(new_n223), .B2(G104), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n217), .A2(KEYINPUT87), .A3(G107), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G101), .ZN(new_n227));
  OAI22_X1  g041(.A1(new_n217), .A2(G107), .B1(KEYINPUT86), .B2(KEYINPUT3), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n221), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n223), .A2(G104), .ZN(new_n230));
  OAI21_X1  g044(.A(G101), .B1(new_n230), .B2(new_n218), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n216), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT10), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  AND2_X1   g050(.A1(KEYINPUT68), .A2(G128), .ZN(new_n237));
  NOR2_X1   g051(.A1(KEYINPUT68), .A2(G128), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n239), .B1(new_n200), .B2(KEYINPUT1), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n198), .A2(new_n199), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n212), .B1(new_n241), .B2(new_n211), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n206), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n233), .A2(KEYINPUT10), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n236), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT64), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT0), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n247), .A3(new_n204), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(KEYINPUT0), .A2(G128), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT65), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT65), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(KEYINPUT0), .A3(G128), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n250), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT67), .B1(new_n242), .B2(new_n256), .ZN(new_n257));
  AND2_X1   g071(.A1(KEYINPUT66), .A2(G146), .ZN(new_n258));
  NOR2_X1   g072(.A1(KEYINPUT66), .A2(G146), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n211), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n212), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT67), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n262), .A2(new_n263), .A3(new_n250), .A4(new_n255), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n258), .A2(new_n259), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n202), .B1(new_n265), .B2(G143), .ZN(new_n266));
  INV_X1    g080(.A(new_n251), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n257), .A2(new_n264), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT86), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT3), .ZN(new_n271));
  AOI22_X1  g085(.A1(new_n270), .A2(new_n271), .B1(new_n223), .B2(G104), .ZN(new_n272));
  XNOR2_X1  g086(.A(KEYINPUT86), .B(KEYINPUT3), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n272), .B1(new_n218), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n227), .B1(new_n274), .B2(new_n226), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n229), .A2(KEYINPUT4), .ZN(new_n276));
  OAI21_X1  g090(.A(KEYINPUT88), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n221), .A2(new_n226), .A3(new_n228), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G101), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT88), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n279), .A2(new_n280), .A3(KEYINPUT4), .A4(new_n229), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT4), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n275), .A2(new_n282), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n269), .A2(new_n277), .A3(new_n281), .A4(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT89), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n279), .A2(KEYINPUT4), .A3(new_n229), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n287), .A2(KEYINPUT88), .B1(new_n282), .B2(new_n275), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n288), .A2(KEYINPUT89), .A3(new_n269), .A4(new_n281), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n245), .B1(new_n286), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT11), .ZN(new_n291));
  INV_X1    g105(.A(G134), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n291), .B1(new_n292), .B2(G137), .ZN(new_n293));
  INV_X1    g107(.A(G137), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n294), .A2(KEYINPUT11), .A3(G134), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n294), .A2(G134), .ZN(new_n297));
  OAI21_X1  g111(.A(G131), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(G131), .B1(new_n292), .B2(G137), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n293), .A2(new_n299), .A3(new_n295), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n197), .B1(new_n290), .B2(new_n302), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n233), .A2(new_n243), .ZN(new_n304));
  AOI22_X1  g118(.A1(new_n206), .A2(new_n207), .B1(new_n210), .B2(new_n214), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n232), .B1(new_n305), .B2(new_n209), .ZN(new_n306));
  OAI211_X1 g120(.A(KEYINPUT12), .B(new_n301), .C1(new_n304), .C2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT91), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OR2_X1    g123(.A1(new_n237), .A2(new_n238), .ZN(new_n310));
  NOR3_X1   g124(.A1(new_n258), .A2(new_n259), .A3(new_n211), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n310), .B1(new_n311), .B2(new_n213), .ZN(new_n312));
  AOI22_X1  g126(.A1(new_n312), .A2(new_n262), .B1(new_n266), .B2(new_n205), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n232), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n302), .B1(new_n234), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(KEYINPUT91), .A3(KEYINPUT12), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n301), .B1(new_n304), .B2(new_n306), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT12), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n309), .A2(new_n316), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT92), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n320), .A2(new_n321), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n303), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT93), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI211_X1 g140(.A(KEYINPUT93), .B(new_n303), .C1(new_n322), .C2(new_n323), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n290), .B(new_n302), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n197), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n326), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G469), .ZN(new_n331));
  INV_X1    g145(.A(G902), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n290), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n320), .B1(new_n334), .B2(new_n301), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n197), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n303), .B1(new_n302), .B2(new_n290), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n331), .B1(new_n338), .B2(new_n332), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n189), .B1(new_n333), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G237), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n194), .A2(G143), .A3(G214), .A4(new_n342), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n191), .A2(new_n193), .A3(G214), .A4(new_n342), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n211), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT95), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(KEYINPUT18), .A3(G131), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n343), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(G125), .B(G140), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n265), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(G125), .ZN(new_n351));
  NOR3_X1   g165(.A1(new_n351), .A2(KEYINPUT79), .A3(G140), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G140), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G125), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n351), .A2(G140), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n355), .A2(new_n356), .A3(KEYINPUT79), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n350), .B1(new_n358), .B2(new_n201), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n348), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n343), .A2(new_n345), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n361), .A2(new_n346), .A3(KEYINPUT18), .A4(G131), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n355), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT16), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n365), .B1(new_n353), .B2(new_n357), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT80), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n358), .A2(new_n368), .A3(KEYINPUT16), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n370), .A2(KEYINPUT81), .A3(G146), .A4(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n352), .B1(new_n349), .B2(KEYINPUT79), .ZN(new_n373));
  OAI21_X1  g187(.A(KEYINPUT80), .B1(new_n373), .B2(new_n365), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n374), .A2(new_n371), .A3(G146), .A4(new_n366), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT81), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n371), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n201), .B1(new_n369), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n372), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G131), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n381), .B1(new_n343), .B2(new_n345), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT17), .ZN(new_n383));
  INV_X1    g197(.A(new_n382), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n343), .A2(new_n381), .A3(new_n345), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n383), .B1(new_n386), .B2(KEYINPUT17), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n363), .B1(new_n380), .B2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(G113), .B(G122), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n389), .B(new_n217), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  AND2_X1   g205(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n390), .B(new_n363), .C1(new_n380), .C2(new_n387), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n332), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G475), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n358), .A2(KEYINPUT19), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n397), .B1(KEYINPUT19), .B2(new_n349), .ZN(new_n398));
  AOI22_X1  g212(.A1(new_n384), .A2(new_n385), .B1(new_n398), .B2(new_n265), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n375), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n363), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT96), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(new_n402), .A3(new_n391), .ZN(new_n403));
  AOI22_X1  g217(.A1(new_n399), .A2(new_n375), .B1(new_n362), .B2(new_n360), .ZN(new_n404));
  OAI21_X1  g218(.A(KEYINPUT96), .B1(new_n404), .B2(new_n390), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n403), .A2(new_n405), .A3(new_n393), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT20), .ZN(new_n407));
  NOR2_X1   g221(.A1(G475), .A2(G902), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n407), .B1(new_n406), .B2(new_n408), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n396), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n211), .A2(G128), .ZN(new_n412));
  XOR2_X1   g226(.A(new_n412), .B(KEYINPUT13), .Z(new_n413));
  NOR2_X1   g227(.A1(new_n310), .A2(new_n211), .ZN(new_n414));
  OAI21_X1  g228(.A(G134), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n412), .B1(new_n310), .B2(new_n211), .ZN(new_n416));
  INV_X1    g230(.A(G122), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n417), .A2(G116), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n417), .A2(G116), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n223), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n421), .A2(new_n223), .ZN(new_n424));
  OAI221_X1 g238(.A(new_n415), .B1(G134), .B2(new_n416), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n416), .B(G134), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n422), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT14), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n420), .B1(new_n418), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(KEYINPUT97), .B1(new_n418), .B2(new_n428), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n418), .A2(KEYINPUT97), .A3(new_n428), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n223), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n425), .B1(new_n427), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(G217), .ZN(new_n435));
  NOR3_X1   g249(.A1(new_n187), .A2(new_n435), .A3(G953), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  OR2_X1    g251(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n434), .A2(new_n437), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n332), .ZN(new_n441));
  INV_X1    g255(.A(G478), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(KEYINPUT15), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n441), .B(new_n443), .ZN(new_n444));
  OR2_X1    g258(.A1(new_n411), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n190), .A2(G952), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n446), .B1(G234), .B2(G237), .ZN(new_n447));
  AOI211_X1 g261(.A(new_n332), .B(new_n194), .C1(G234), .C2(G237), .ZN(new_n448));
  XNOR2_X1  g262(.A(KEYINPUT21), .B(G898), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n445), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(G214), .B1(G237), .B2(G902), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  XOR2_X1   g267(.A(G116), .B(G119), .Z(new_n454));
  XNOR2_X1  g268(.A(KEYINPUT2), .B(G113), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XOR2_X1   g270(.A(KEYINPUT2), .B(G113), .Z(new_n457));
  XNOR2_X1  g271(.A(G116), .B(G119), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n277), .A2(new_n281), .A3(new_n460), .A4(new_n283), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT5), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n454), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(G116), .ZN(new_n464));
  OAI21_X1  g278(.A(G113), .B1(new_n464), .B2(G119), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n459), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  OR2_X1    g280(.A1(new_n466), .A2(new_n232), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n461), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(G110), .B(G122), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n461), .A2(new_n469), .A3(new_n467), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(KEYINPUT6), .A3(new_n472), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n351), .B(new_n206), .C1(new_n240), .C2(new_n242), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n257), .A2(new_n264), .A3(new_n268), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n475), .B1(new_n476), .B2(G125), .ZN(new_n477));
  INV_X1    g291(.A(G224), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n478), .A2(G953), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n477), .B(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT6), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n468), .A2(new_n482), .A3(new_n470), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n473), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  XOR2_X1   g298(.A(new_n469), .B(KEYINPUT8), .Z(new_n485));
  NAND2_X1  g299(.A1(new_n466), .A2(new_n232), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n485), .B1(new_n467), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n480), .A2(KEYINPUT94), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT7), .ZN(new_n490));
  OAI22_X1  g304(.A1(new_n477), .A2(new_n489), .B1(new_n490), .B2(new_n479), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n479), .A2(new_n490), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n262), .A2(new_n250), .A3(new_n255), .ZN(new_n493));
  AOI22_X1  g307(.A1(new_n493), .A2(KEYINPUT67), .B1(new_n266), .B2(new_n267), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n351), .B1(new_n494), .B2(new_n264), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n492), .B(new_n488), .C1(new_n495), .C2(new_n475), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n487), .B1(new_n491), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(G902), .B1(new_n497), .B2(new_n472), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n484), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(G210), .B1(G237), .B2(G902), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n484), .A2(new_n498), .A3(new_n500), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n453), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n341), .A2(new_n451), .A3(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT98), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n505), .B(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(G472), .ZN(new_n508));
  AOI21_X1  g322(.A(KEYINPUT72), .B1(new_n456), .B2(new_n459), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n456), .A2(new_n459), .A3(KEYINPUT72), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n292), .A2(G137), .ZN(new_n513));
  OAI21_X1  g327(.A(G131), .B1(new_n513), .B2(new_n297), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n514), .A2(new_n300), .A3(KEYINPUT69), .ZN(new_n515));
  AOI21_X1  g329(.A(KEYINPUT69), .B1(new_n514), .B2(new_n300), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n512), .B1(new_n243), .B2(new_n518), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n257), .A2(new_n301), .A3(new_n264), .A4(new_n268), .ZN(new_n520));
  AOI21_X1  g334(.A(KEYINPUT28), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT70), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n522), .B1(new_n517), .B2(new_n313), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n243), .B(KEYINPUT70), .C1(new_n516), .C2(new_n515), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(new_n520), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n512), .ZN(new_n526));
  INV_X1    g340(.A(new_n511), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n527), .A2(new_n509), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n523), .A2(new_n520), .A3(new_n524), .A4(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT28), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT77), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n530), .A2(KEYINPUT77), .A3(KEYINPUT28), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n521), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n191), .A2(new_n193), .A3(G210), .A4(new_n342), .ZN(new_n536));
  OR2_X1    g350(.A1(new_n536), .A2(KEYINPUT27), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT26), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(KEYINPUT27), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n538), .B1(new_n537), .B2(new_n539), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n227), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n537), .A2(new_n539), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT26), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n545), .A2(G101), .A3(new_n540), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n547), .A2(KEYINPUT29), .ZN(new_n548));
  AOI21_X1  g362(.A(G902), .B1(new_n535), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n460), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n514), .A2(new_n300), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n243), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n520), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT30), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n550), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n523), .A2(KEYINPUT30), .A3(new_n520), .A4(new_n524), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT71), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n555), .A2(new_n556), .A3(KEYINPUT71), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n529), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT76), .ZN(new_n563));
  INV_X1    g377(.A(new_n547), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n529), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n566), .B1(new_n559), .B2(new_n560), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT76), .B1(new_n567), .B2(new_n547), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT28), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n553), .A2(new_n460), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n569), .B1(new_n529), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(new_n521), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT29), .B1(new_n572), .B2(new_n547), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n565), .A2(new_n568), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n508), .B1(new_n549), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(G472), .A2(G902), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT31), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n547), .A2(new_n529), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n577), .B1(new_n561), .B2(new_n578), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n555), .A2(new_n556), .A3(KEYINPUT71), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT71), .B1(new_n555), .B2(new_n556), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n577), .B(new_n578), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n564), .B1(new_n571), .B2(new_n521), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT74), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI211_X1 g401(.A(KEYINPUT74), .B(new_n564), .C1(new_n571), .C2(new_n521), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(KEYINPUT75), .B1(new_n584), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n578), .B1(new_n580), .B2(new_n581), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT31), .ZN(new_n592));
  AND4_X1   g406(.A1(KEYINPUT75), .A2(new_n589), .A3(new_n592), .A4(new_n582), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n576), .B1(new_n590), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT32), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n575), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI211_X1 g410(.A(KEYINPUT32), .B(new_n576), .C1(new_n590), .C2(new_n593), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT78), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n576), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT75), .ZN(new_n601));
  INV_X1    g415(.A(new_n589), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n592), .A2(new_n582), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n589), .A2(KEYINPUT75), .A3(new_n592), .A4(new_n582), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n600), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n606), .A2(KEYINPUT78), .A3(KEYINPUT32), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n596), .A2(new_n599), .A3(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n239), .A2(KEYINPUT23), .A3(G119), .ZN(new_n609));
  AOI21_X1  g423(.A(KEYINPUT23), .B1(new_n204), .B2(G119), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n204), .A2(G119), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n611), .B1(new_n239), .B2(G119), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT24), .B(G110), .Z(new_n615));
  AOI22_X1  g429(.A1(new_n613), .A2(G110), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n380), .A2(new_n616), .ZN(new_n617));
  OAI22_X1  g431(.A1(new_n613), .A2(G110), .B1(new_n614), .B2(new_n615), .ZN(new_n618));
  OR2_X1    g432(.A1(new_n618), .A2(KEYINPUT82), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(KEYINPUT82), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n619), .A2(new_n375), .A3(new_n620), .A4(new_n350), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n194), .A2(G221), .A3(G234), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT22), .B(G137), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT83), .B(KEYINPUT84), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n622), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n617), .A2(new_n621), .A3(new_n627), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n435), .B1(G234), .B2(new_n332), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(G902), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(new_n634), .B(KEYINPUT85), .Z(new_n635));
  NAND3_X1  g449(.A1(new_n629), .A2(new_n332), .A3(new_n630), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(KEYINPUT25), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT25), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n629), .A2(new_n638), .A3(new_n332), .A4(new_n630), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n637), .A2(new_n639), .A3(new_n632), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n635), .A2(new_n640), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n608), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n507), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G101), .ZN(G3));
  NAND2_X1  g458(.A1(new_n604), .A2(new_n605), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n508), .B1(new_n645), .B2(new_n332), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n646), .A2(new_n606), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n647), .A2(new_n641), .A3(new_n341), .ZN(new_n648));
  INV_X1    g462(.A(new_n450), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT33), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n650), .A2(KEYINPUT99), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n440), .A2(new_n652), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n650), .A2(KEYINPUT99), .ZN(new_n654));
  OAI211_X1 g468(.A(new_n438), .B(new_n439), .C1(new_n654), .C2(new_n651), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n442), .A2(G902), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n653), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(KEYINPUT100), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT100), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n653), .A2(new_n659), .A3(new_n655), .A4(new_n656), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n441), .A2(new_n442), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n658), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n662), .A2(new_n411), .A3(KEYINPUT101), .ZN(new_n663));
  AOI21_X1  g477(.A(KEYINPUT101), .B1(new_n662), .B2(new_n411), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n649), .B(new_n504), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n648), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT102), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT34), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G104), .ZN(G6));
  XOR2_X1   g484(.A(new_n450), .B(KEYINPUT103), .Z(new_n671));
  NAND2_X1  g485(.A1(new_n504), .A2(new_n671), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n444), .B(new_n396), .C1(new_n410), .C2(new_n409), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n648), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT35), .B(G107), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G9));
  NOR2_X1   g491(.A1(new_n628), .A2(KEYINPUT36), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n622), .B(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n633), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n640), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n647), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n507), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(new_n684), .B(KEYINPUT37), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT104), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G110), .ZN(G12));
  INV_X1    g501(.A(G900), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n447), .B1(new_n448), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(KEYINPUT105), .B1(new_n673), .B2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n411), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n692));
  INV_X1    g506(.A(new_n689), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n691), .A2(new_n692), .A3(new_n444), .A4(new_n693), .ZN(new_n694));
  AND2_X1   g508(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n681), .A2(new_n504), .ZN(new_n696));
  AOI211_X1 g510(.A(new_n189), .B(new_n696), .C1(new_n333), .C2(new_n340), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n608), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G128), .ZN(G30));
  XOR2_X1   g513(.A(new_n689), .B(KEYINPUT39), .Z(new_n700));
  NAND2_X1  g514(.A1(new_n341), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(new_n701), .B(KEYINPUT40), .Z(new_n702));
  NAND2_X1  g516(.A1(new_n599), .A2(new_n607), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n562), .A2(new_n547), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n564), .A2(new_n529), .A3(new_n526), .ZN(new_n705));
  AOI21_X1  g519(.A(KEYINPUT106), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OAI211_X1 g520(.A(KEYINPUT106), .B(new_n705), .C1(new_n567), .C2(new_n564), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n332), .ZN(new_n708));
  OAI21_X1  g522(.A(G472), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT107), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OAI211_X1 g525(.A(KEYINPUT107), .B(G472), .C1(new_n706), .C2(new_n708), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n711), .B(new_n712), .C1(KEYINPUT32), .C2(new_n606), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n703), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n714), .A2(new_n681), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n502), .A2(new_n503), .ZN(new_n716));
  XOR2_X1   g530(.A(new_n716), .B(KEYINPUT38), .Z(new_n717));
  NAND2_X1  g531(.A1(new_n411), .A2(new_n444), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n717), .A2(new_n453), .A3(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n702), .A2(new_n715), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G143), .ZN(G45));
  NAND2_X1  g535(.A1(new_n662), .A2(new_n411), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n722), .A2(new_n689), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n608), .A2(new_n697), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G146), .ZN(G48));
  NAND2_X1  g539(.A1(new_n330), .A2(new_n332), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(G469), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n727), .A2(new_n188), .A3(new_n333), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n666), .A2(new_n608), .A3(new_n641), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(KEYINPUT41), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G113), .ZN(G15));
  NAND4_X1  g545(.A1(new_n608), .A2(new_n641), .A3(new_n674), .A4(new_n728), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(KEYINPUT108), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G116), .ZN(G18));
  INV_X1    g548(.A(new_n696), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n608), .A2(new_n451), .A3(new_n735), .A4(new_n728), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G119), .ZN(G21));
  NAND2_X1  g551(.A1(new_n533), .A2(new_n534), .ZN(new_n738));
  INV_X1    g552(.A(new_n521), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n547), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n576), .B1(new_n740), .B2(new_n603), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT109), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT109), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n743), .B(new_n576), .C1(new_n740), .C2(new_n603), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n646), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n672), .A2(new_n718), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n728), .A2(new_n746), .A3(new_n641), .A4(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G122), .ZN(G24));
  NAND4_X1  g563(.A1(new_n728), .A2(new_n746), .A3(new_n735), .A4(new_n723), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G125), .ZN(G27));
  AOI22_X1  g565(.A1(new_n324), .A2(new_n325), .B1(new_n328), .B2(new_n197), .ZN(new_n752));
  AOI21_X1  g566(.A(G902), .B1(new_n752), .B2(new_n327), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n339), .B1(new_n753), .B2(new_n331), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n716), .A2(new_n453), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n754), .A2(new_n189), .A3(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(KEYINPUT42), .A3(new_n723), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n759), .B1(new_n606), .B2(KEYINPUT32), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n575), .B1(new_n606), .B2(KEYINPUT32), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n594), .A2(KEYINPUT110), .A3(new_n595), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n641), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(KEYINPUT111), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT111), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n763), .A2(new_n766), .A3(new_n641), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n758), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n608), .A2(new_n757), .A3(new_n641), .A4(new_n723), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT42), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT112), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n768), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n758), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n763), .A2(new_n766), .A3(new_n641), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n766), .B1(new_n763), .B2(new_n641), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n769), .A2(new_n770), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT112), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n773), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G131), .ZN(G33));
  AND4_X1   g595(.A1(new_n608), .A2(new_n757), .A3(new_n641), .A4(new_n695), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(new_n292), .ZN(G36));
  INV_X1    g597(.A(new_n681), .ZN(new_n784));
  OR3_X1    g598(.A1(new_n647), .A2(KEYINPUT114), .A3(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(KEYINPUT114), .B1(new_n647), .B2(new_n784), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n691), .A2(new_n662), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT113), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT43), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(KEYINPUT113), .A2(KEYINPUT43), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n788), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n787), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT44), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n787), .B(KEYINPUT44), .C1(new_n794), .C2(new_n796), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT46), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT45), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n331), .B1(new_n338), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n336), .A2(KEYINPUT45), .A3(new_n337), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n331), .A2(new_n332), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n801), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n333), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n805), .A2(new_n801), .A3(new_n806), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n188), .B(new_n700), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n799), .A2(new_n755), .A3(new_n800), .A4(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT115), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(new_n294), .ZN(G39));
  OAI21_X1  g628(.A(new_n188), .B1(new_n808), .B2(new_n809), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT47), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT47), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n817), .B(new_n188), .C1(new_n808), .C2(new_n809), .ZN(new_n818));
  INV_X1    g632(.A(new_n723), .ZN(new_n819));
  NOR4_X1   g633(.A1(new_n608), .A2(new_n641), .A3(new_n819), .A4(new_n756), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n816), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(G140), .ZN(G42));
  INV_X1    g636(.A(new_n788), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n641), .A2(new_n188), .A3(new_n452), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(KEYINPUT116), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n825), .A2(new_n717), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n727), .A2(new_n333), .ZN(new_n827));
  XOR2_X1   g641(.A(new_n827), .B(KEYINPUT49), .Z(new_n828));
  OR2_X1    g642(.A1(new_n824), .A2(KEYINPUT116), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n826), .A2(new_n714), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n698), .A2(new_n750), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n504), .A2(new_n411), .A3(new_n444), .A4(new_n693), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n754), .A2(new_n189), .A3(new_n833), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n834), .B(new_n784), .C1(new_n703), .C2(new_n713), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n832), .A2(KEYINPUT52), .A3(new_n724), .A4(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n835), .A2(new_n698), .A3(new_n724), .A4(new_n750), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT52), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n772), .B1(new_n768), .B2(new_n771), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n777), .A2(KEYINPUT112), .A3(new_n778), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n445), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n608), .A2(new_n844), .A3(new_n693), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n746), .A2(new_n723), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n757), .A2(new_n681), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n782), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n722), .A2(new_n673), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n851), .A2(new_n672), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n852), .A2(new_n647), .A3(new_n641), .A4(new_n341), .ZN(new_n853));
  AND4_X1   g667(.A1(new_n729), .A2(new_n736), .A3(new_n748), .A4(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n507), .B1(new_n642), .B2(new_n683), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n733), .A2(new_n849), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n831), .B1(new_n843), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT54), .ZN(new_n858));
  AND4_X1   g672(.A1(new_n733), .A2(new_n849), .A3(new_n854), .A4(new_n855), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n831), .B1(new_n777), .B2(new_n778), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n859), .A2(new_n840), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n857), .A2(new_n858), .A3(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n780), .A2(new_n859), .A3(KEYINPUT53), .A4(new_n840), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n858), .B1(new_n857), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT117), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n862), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI211_X1 g680(.A(KEYINPUT117), .B(new_n858), .C1(new_n857), .C2(new_n863), .ZN(new_n867));
  INV_X1    g681(.A(new_n447), .ZN(new_n868));
  INV_X1    g682(.A(new_n794), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n868), .B1(new_n869), .B2(new_n795), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n827), .A2(new_n189), .A3(new_n756), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT118), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n870), .A2(new_n871), .A3(KEYINPUT118), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n765), .A2(new_n767), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(KEYINPUT121), .A2(KEYINPUT48), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AND2_X1   g694(.A1(KEYINPUT121), .A2(KEYINPUT48), .ZN(new_n881));
  OR3_X1    g695(.A1(new_n878), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n746), .A2(new_n641), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n883), .A2(new_n728), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n884), .A2(new_n504), .A3(new_n870), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT120), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n884), .A2(KEYINPUT120), .A3(new_n504), .A4(new_n870), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n446), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n714), .A2(new_n871), .A3(new_n641), .A4(new_n447), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT119), .ZN(new_n891));
  OR2_X1    g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n890), .A2(new_n891), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n892), .B(new_n893), .C1(new_n664), .C2(new_n663), .ZN(new_n894));
  AND4_X1   g708(.A1(new_n880), .A2(new_n882), .A3(new_n889), .A4(new_n894), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n870), .A2(new_n755), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n816), .A2(new_n818), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n827), .A2(new_n188), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n883), .B(new_n896), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n717), .A2(new_n453), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n883), .A2(new_n728), .A3(new_n870), .A4(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT50), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n901), .A2(new_n902), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n745), .A2(new_n646), .A3(new_n784), .ZN(new_n905));
  AOI22_X1  g719(.A1(new_n903), .A2(new_n904), .B1(new_n876), .B2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(new_n662), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n892), .A2(new_n691), .A3(new_n907), .A4(new_n893), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n899), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n909), .A2(KEYINPUT51), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n909), .A2(KEYINPUT51), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n895), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n866), .A2(new_n867), .A3(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(G952), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n190), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT122), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n830), .B1(new_n913), .B2(new_n916), .ZN(G75));
  INV_X1    g731(.A(new_n194), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n914), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT123), .Z(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT56), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n857), .A2(new_n861), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(G902), .ZN(new_n924));
  INV_X1    g738(.A(G210), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n922), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n473), .A2(new_n483), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(new_n481), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT55), .Z(new_n929));
  NAND2_X1  g743(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n929), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n922), .B(new_n931), .C1(new_n924), .C2(new_n925), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n921), .B1(new_n930), .B2(new_n932), .ZN(G51));
  XNOR2_X1  g747(.A(new_n806), .B(KEYINPUT57), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n857), .A2(new_n858), .A3(new_n861), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n858), .B1(new_n857), .B2(new_n861), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n330), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n332), .B1(new_n857), .B2(new_n861), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n805), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n921), .B1(new_n938), .B2(new_n940), .ZN(G54));
  AND2_X1   g755(.A1(KEYINPUT58), .A2(G475), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n939), .A2(new_n406), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n406), .B1(new_n939), .B2(new_n942), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n943), .A2(new_n944), .A3(new_n921), .ZN(G60));
  NAND2_X1  g759(.A1(new_n653), .A2(new_n655), .ZN(new_n946));
  NAND2_X1  g760(.A1(G478), .A2(G902), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT59), .Z(new_n948));
  NOR2_X1   g762(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n949), .B1(new_n935), .B2(new_n936), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n920), .ZN(new_n951));
  INV_X1    g765(.A(new_n948), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n952), .B1(new_n866), .B2(new_n867), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n951), .B1(new_n953), .B2(new_n946), .ZN(G63));
  INV_X1    g768(.A(KEYINPUT61), .ZN(new_n955));
  NAND2_X1  g769(.A1(G217), .A2(G902), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT60), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n957), .B1(new_n857), .B2(new_n861), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n679), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n920), .B1(new_n958), .B2(new_n631), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n955), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n958), .A2(new_n631), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n963), .A2(KEYINPUT61), .A3(new_n920), .A4(new_n959), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n962), .A2(new_n964), .ZN(G66));
  NAND3_X1  g779(.A1(new_n733), .A2(new_n854), .A3(new_n855), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n194), .ZN(new_n967));
  OAI21_X1  g781(.A(G953), .B1(new_n449), .B2(new_n478), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OR2_X1    g783(.A1(new_n969), .A2(KEYINPUT124), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(KEYINPUT124), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(KEYINPUT125), .ZN(new_n973));
  INV_X1    g787(.A(G898), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n927), .B1(new_n974), .B2(new_n918), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT125), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n970), .A2(new_n976), .A3(new_n971), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n973), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n975), .B1(new_n973), .B2(new_n977), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n978), .A2(new_n979), .ZN(G69));
  AOI21_X1  g794(.A(new_n194), .B1(G227), .B2(G900), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n832), .A2(new_n724), .ZN(new_n982));
  AND3_X1   g796(.A1(new_n504), .A2(new_n444), .A3(new_n411), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n877), .A2(new_n811), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n821), .ZN(new_n986));
  NOR3_X1   g800(.A1(new_n985), .A2(new_n782), .A3(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n987), .A2(new_n780), .A3(new_n812), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n988), .A2(new_n194), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n553), .A2(new_n554), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n556), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(new_n398), .ZN(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n993), .B1(G900), .B2(new_n194), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT62), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n982), .A2(new_n720), .A3(new_n995), .ZN(new_n996));
  NOR3_X1   g810(.A1(new_n701), .A2(new_n756), .A3(new_n851), .ZN(new_n997));
  AOI22_X1  g811(.A1(new_n897), .A2(new_n820), .B1(new_n642), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n812), .A2(new_n996), .A3(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT126), .ZN(new_n1000));
  INV_X1    g814(.A(new_n720), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n832), .A2(new_n724), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n1000), .B(KEYINPUT62), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(KEYINPUT62), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(KEYINPUT126), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n999), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n992), .A2(new_n194), .ZN(new_n1007));
  OAI22_X1  g821(.A1(new_n989), .A2(new_n994), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n981), .B1(new_n1008), .B2(KEYINPUT127), .ZN(new_n1009));
  INV_X1    g823(.A(new_n999), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1005), .A2(new_n1003), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1007), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n994), .B1(new_n988), .B2(new_n194), .ZN(new_n1013));
  OAI211_X1 g827(.A(KEYINPUT127), .B(new_n981), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1014), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n1009), .A2(new_n1015), .ZN(G72));
  NAND2_X1  g830(.A1(G472), .A2(G902), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1017), .B(KEYINPUT63), .Z(new_n1018));
  OAI21_X1  g832(.A(new_n1018), .B1(new_n988), .B2(new_n966), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1019), .A2(new_n564), .A3(new_n567), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1020), .A2(new_n920), .ZN(new_n1021));
  INV_X1    g835(.A(new_n966), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1006), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n704), .B1(new_n1023), .B2(new_n1018), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n565), .A2(new_n591), .A3(new_n568), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1025), .A2(new_n1018), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1026), .B1(new_n857), .B2(new_n863), .ZN(new_n1027));
  NOR3_X1   g841(.A1(new_n1021), .A2(new_n1024), .A3(new_n1027), .ZN(G57));
endmodule


