

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818;

  NOR2_X1 U371 ( .A1(n413), .A2(n410), .ZN(n463) );
  OR2_X1 U372 ( .A1(n660), .A2(KEYINPUT106), .ZN(n360) );
  XNOR2_X1 U373 ( .A(n754), .B(KEYINPUT79), .ZN(n660) );
  INV_X1 U374 ( .A(n621), .ZN(n350) );
  BUF_X1 U375 ( .A(G146), .Z(n349) );
  XNOR2_X2 U376 ( .A(n631), .B(KEYINPUT31), .ZN(n723) );
  XNOR2_X1 U377 ( .A(n526), .B(n525), .ZN(n353) );
  NAND2_X1 U378 ( .A1(n353), .A2(n712), .ZN(n643) );
  NAND2_X1 U379 ( .A1(n643), .A2(KEYINPUT44), .ZN(n477) );
  AND2_X2 U380 ( .A1(n348), .A2(n473), .ZN(n470) );
  AND2_X2 U381 ( .A1(n493), .A2(n516), .ZN(n348) );
  NAND2_X4 U382 ( .A1(G214), .A2(n593), .ZN(n749) );
  XOR2_X2 U383 ( .A(KEYINPUT45), .B(KEYINPUT82), .Z(n384) );
  INV_X2 U384 ( .A(G143), .ZN(n511) );
  NOR2_X2 U385 ( .A1(n752), .A2(n753), .ZN(n676) );
  XNOR2_X2 U386 ( .A(n451), .B(n671), .ZN(n680) );
  OR2_X2 U387 ( .A1(n763), .A2(n677), .ZN(n400) );
  OR2_X1 U388 ( .A1(n418), .A2(KEYINPUT77), .ZN(n416) );
  INV_X2 U389 ( .A(G116), .ZN(n575) );
  XNOR2_X2 U390 ( .A(n616), .B(n615), .ZN(n803) );
  XNOR2_X2 U391 ( .A(n351), .B(n350), .ZN(n630) );
  OR2_X2 U392 ( .A1(n781), .A2(G902), .ZN(n351) );
  AND2_X4 U393 ( .A1(n679), .A2(n672), .ZN(n754) );
  XNOR2_X2 U394 ( .A(n713), .B(KEYINPUT105), .ZN(n679) );
  XOR2_X1 U395 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n558) );
  XNOR2_X1 U396 ( .A(KEYINPUT4), .B(KEYINPUT66), .ZN(n510) );
  XOR2_X1 U397 ( .A(KEYINPUT80), .B(KEYINPUT8), .Z(n543) );
  XNOR2_X1 U398 ( .A(G107), .B(G110), .ZN(n554) );
  XNOR2_X1 U399 ( .A(G902), .B(KEYINPUT15), .ZN(n688) );
  BUF_X1 U400 ( .A(G116), .Z(n475) );
  BUF_X1 U401 ( .A(G143), .Z(n478) );
  AND2_X1 U402 ( .A1(n374), .A2(KEYINPUT85), .ZN(n352) );
  XNOR2_X2 U403 ( .A(n580), .B(KEYINPUT10), .ZN(n615) );
  NAND2_X2 U404 ( .A1(n388), .A2(n377), .ZN(n387) );
  XNOR2_X1 U405 ( .A(n538), .B(n537), .ZN(n664) );
  NOR2_X2 U406 ( .A1(G953), .A2(G237), .ZN(n611) );
  NOR2_X1 U407 ( .A1(n795), .A2(n805), .ZN(n453) );
  NOR2_X1 U408 ( .A1(n815), .A2(n818), .ZN(n678) );
  XNOR2_X1 U409 ( .A(n400), .B(n399), .ZN(n818) );
  NOR2_X1 U410 ( .A1(n817), .A2(n378), .ZN(n536) );
  NOR2_X1 U411 ( .A1(n626), .A2(n664), .ZN(n735) );
  XNOR2_X1 U412 ( .A(n513), .B(KEYINPUT1), .ZN(n734) );
  NOR2_X1 U413 ( .A1(n697), .A2(G902), .ZN(n566) );
  XNOR2_X1 U414 ( .A(n439), .B(n555), .ZN(n779) );
  XNOR2_X1 U415 ( .A(n561), .B(n440), .ZN(n578) );
  XNOR2_X1 U416 ( .A(n491), .B(G122), .ZN(n617) );
  INV_X1 U417 ( .A(G113), .ZN(n441) );
  NOR2_X2 U418 ( .A1(n795), .A2(n449), .ZN(n733) );
  XNOR2_X1 U419 ( .A(n409), .B(n528), .ZN(n527) );
  XNOR2_X1 U420 ( .A(n658), .B(KEYINPUT78), .ZN(n418) );
  AND2_X1 U421 ( .A1(n529), .A2(n727), .ZN(n460) );
  INV_X1 U422 ( .A(n639), .ZN(n641) );
  NAND2_X1 U423 ( .A1(n423), .A2(n419), .ZN(n659) );
  AND2_X1 U424 ( .A1(n424), .A2(n425), .ZN(n423) );
  AND2_X1 U425 ( .A1(n685), .A2(n730), .ZN(n686) );
  NAND2_X1 U426 ( .A1(n396), .A2(n393), .ZN(n815) );
  AND2_X1 U427 ( .A1(n398), .A2(n397), .ZN(n396) );
  NAND2_X1 U428 ( .A1(n395), .A2(n394), .ZN(n393) );
  NAND2_X1 U429 ( .A1(n422), .A2(n420), .ZN(n419) );
  AND2_X1 U430 ( .A1(n536), .A2(KEYINPUT77), .ZN(n415) );
  XNOR2_X1 U431 ( .A(n652), .B(KEYINPUT111), .ZN(n817) );
  INV_X2 U432 ( .A(n391), .ZN(n683) );
  XNOR2_X1 U433 ( .A(n369), .B(KEYINPUT74), .ZN(n635) );
  NAND2_X1 U434 ( .A1(n497), .A2(n380), .ZN(n496) );
  INV_X1 U435 ( .A(n557), .ZN(n354) );
  AND2_X1 U436 ( .A1(n506), .A2(KEYINPUT85), .ZN(n505) );
  XNOR2_X1 U437 ( .A(n371), .B(n454), .ZN(n370) );
  XNOR2_X1 U438 ( .A(n402), .B(n401), .ZN(n670) );
  XNOR2_X1 U439 ( .A(n457), .B(n456), .ZN(n557) );
  NOR2_X1 U440 ( .A1(n654), .A2(n655), .ZN(n484) );
  NAND2_X1 U441 ( .A1(n734), .A2(n735), .ZN(n457) );
  BUF_X1 U442 ( .A(n513), .Z(n512) );
  XNOR2_X1 U443 ( .A(n607), .B(n608), .ZN(n629) );
  XNOR2_X1 U444 ( .A(n372), .B(n539), .ZN(n782) );
  XNOR2_X1 U445 ( .A(n697), .B(KEYINPUT62), .ZN(n698) );
  XNOR2_X1 U446 ( .A(n605), .B(n362), .ZN(n785) );
  XNOR2_X1 U447 ( .A(n604), .B(n606), .ZN(n362) );
  XNOR2_X1 U448 ( .A(n434), .B(n432), .ZN(n788) );
  XNOR2_X1 U449 ( .A(n545), .B(n544), .ZN(n434) );
  XNOR2_X1 U450 ( .A(n441), .B(G119), .ZN(n440) );
  XNOR2_X1 U451 ( .A(n511), .B(G128), .ZN(n390) );
  XNOR2_X1 U452 ( .A(G122), .B(KEYINPUT102), .ZN(n474) );
  XOR2_X1 U453 ( .A(KEYINPUT65), .B(G101), .Z(n584) );
  XNOR2_X1 U454 ( .A(KEYINPUT7), .B(KEYINPUT103), .ZN(n599) );
  INV_X2 U455 ( .A(G953), .ZN(n806) );
  INV_X4 U456 ( .A(G104), .ZN(n491) );
  XNOR2_X1 U457 ( .A(n353), .B(G119), .ZN(G21) );
  NOR2_X2 U458 ( .A1(n700), .A2(n790), .ZN(n703) );
  NOR2_X2 U459 ( .A1(n784), .A2(n790), .ZN(n363) );
  NOR2_X2 U460 ( .A1(n776), .A2(n790), .ZN(n364) );
  NAND2_X1 U461 ( .A1(n356), .A2(n435), .ZN(n355) );
  NAND2_X1 U462 ( .A1(n354), .A2(n518), .ZN(n520) );
  INV_X1 U463 ( .A(G143), .ZN(n368) );
  NAND2_X1 U464 ( .A1(n361), .A2(n360), .ZN(n358) );
  AND2_X1 U465 ( .A1(n359), .A2(n358), .ZN(n357) );
  NAND2_X1 U466 ( .A1(n357), .A2(n355), .ZN(n634) );
  INV_X1 U467 ( .A(n723), .ZN(n356) );
  NAND2_X1 U468 ( .A1(n723), .A2(n381), .ZN(n359) );
  NAND2_X1 U469 ( .A1(n436), .A2(n660), .ZN(n361) );
  NOR2_X1 U470 ( .A1(n352), .A2(n505), .ZN(n388) );
  XNOR2_X1 U471 ( .A(n363), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U472 ( .A(n364), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X2 U473 ( .A(n366), .B(n692), .ZN(n696) );
  NAND2_X2 U474 ( .A1(n691), .A2(n690), .ZN(n366) );
  NAND2_X1 U475 ( .A1(n367), .A2(n627), .ZN(n628) );
  AND2_X1 U476 ( .A1(n367), .A2(n520), .ZN(n519) );
  NAND2_X1 U477 ( .A1(n367), .A2(n633), .ZN(n709) );
  AND2_X1 U478 ( .A1(n367), .A2(n467), .ZN(n631) );
  XNOR2_X2 U479 ( .A(n476), .B(n383), .ZN(n367) );
  NAND2_X1 U480 ( .A1(n370), .A2(n523), .ZN(n369) );
  NAND2_X1 U481 ( .A1(n489), .A2(n386), .ZN(n371) );
  BUF_X1 U482 ( .A(n781), .Z(n372) );
  BUF_X1 U483 ( .A(n798), .Z(n373) );
  XNOR2_X1 U484 ( .A(n628), .B(KEYINPUT22), .ZN(n374) );
  XNOR2_X1 U485 ( .A(n628), .B(KEYINPUT22), .ZN(n636) );
  BUF_X1 U486 ( .A(n704), .Z(n375) );
  AND2_X1 U487 ( .A1(n660), .A2(n437), .ZN(n435) );
  AND2_X1 U488 ( .A1(n634), .A2(KEYINPUT107), .ZN(n492) );
  XOR2_X1 U489 ( .A(G131), .B(G140), .Z(n616) );
  INV_X1 U490 ( .A(G469), .ZN(n524) );
  XNOR2_X1 U491 ( .A(n547), .B(n548), .ZN(n537) );
  NAND2_X1 U492 ( .A1(n412), .A2(n535), .ZN(n411) );
  NAND2_X1 U493 ( .A1(KEYINPUT87), .A2(n640), .ZN(n516) );
  NOR2_X1 U494 ( .A1(n408), .A2(n472), .ZN(n471) );
  OR2_X1 U495 ( .A1(G237), .A2(G902), .ZN(n593) );
  INV_X1 U496 ( .A(KEYINPUT75), .ZN(n426) );
  XOR2_X1 U497 ( .A(KEYINPUT101), .B(KEYINPUT9), .Z(n600) );
  NAND2_X1 U498 ( .A1(n460), .A2(n461), .ZN(n409) );
  INV_X1 U499 ( .A(KEYINPUT69), .ZN(n462) );
  NOR2_X1 U500 ( .A1(n523), .A2(n567), .ZN(n518) );
  NAND2_X1 U501 ( .A1(n455), .A2(n486), .ZN(n746) );
  INV_X1 U502 ( .A(n457), .ZN(n455) );
  NOR2_X1 U503 ( .A1(n664), .A2(n653), .ZN(n404) );
  XNOR2_X1 U504 ( .A(n407), .B(n406), .ZN(n405) );
  INV_X1 U505 ( .A(KEYINPUT30), .ZN(n406) );
  NAND2_X1 U506 ( .A1(n741), .A2(n749), .ZN(n407) );
  NAND2_X1 U507 ( .A1(n504), .A2(n507), .ZN(n503) );
  XNOR2_X1 U508 ( .A(G140), .B(KEYINPUT95), .ZN(n531) );
  XNOR2_X1 U509 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n532) );
  XNOR2_X1 U510 ( .A(n534), .B(n533), .ZN(n433) );
  XNOR2_X1 U511 ( .A(G119), .B(G137), .ZN(n533) );
  XNOR2_X1 U512 ( .A(n483), .B(G110), .ZN(n534) );
  INV_X1 U513 ( .A(G128), .ZN(n483) );
  XNOR2_X1 U514 ( .A(G113), .B(n478), .ZN(n609) );
  XNOR2_X1 U515 ( .A(n613), .B(n612), .ZN(n614) );
  XOR2_X1 U516 ( .A(KEYINPUT98), .B(KEYINPUT100), .Z(n613) );
  XNOR2_X1 U517 ( .A(n674), .B(n673), .ZN(n675) );
  INV_X1 U518 ( .A(KEYINPUT113), .ZN(n673) );
  NAND2_X1 U519 ( .A1(n672), .A2(n382), .ZN(n397) );
  INV_X1 U520 ( .A(KEYINPUT108), .ZN(n454) );
  BUF_X1 U521 ( .A(n779), .Z(n487) );
  NOR2_X1 U522 ( .A1(G952), .A2(n806), .ZN(n790) );
  XNOR2_X1 U523 ( .A(n695), .B(n450), .ZN(n449) );
  INV_X1 U524 ( .A(KEYINPUT83), .ZN(n450) );
  INV_X1 U525 ( .A(KEYINPUT106), .ZN(n437) );
  NOR2_X1 U526 ( .A1(n386), .A2(KEYINPUT107), .ZN(n385) );
  AND2_X1 U527 ( .A1(n517), .A2(KEYINPUT44), .ZN(n515) );
  NAND2_X1 U528 ( .A1(n379), .A2(n411), .ZN(n410) );
  INV_X1 U529 ( .A(KEYINPUT68), .ZN(n446) );
  INV_X1 U530 ( .A(KEYINPUT86), .ZN(n459) );
  INV_X1 U531 ( .A(KEYINPUT109), .ZN(n456) );
  XNOR2_X1 U532 ( .A(n475), .B(G131), .ZN(n562) );
  XOR2_X1 U533 ( .A(G137), .B(G134), .Z(n549) );
  XNOR2_X1 U534 ( .A(n551), .B(n491), .ZN(n552) );
  INV_X1 U535 ( .A(KEYINPUT48), .ZN(n528) );
  NAND2_X1 U536 ( .A1(n501), .A2(n687), .ZN(n499) );
  NAND2_X1 U537 ( .A1(n512), .A2(KEYINPUT75), .ZN(n421) );
  NAND2_X1 U538 ( .A1(n427), .A2(n426), .ZN(n425) );
  INV_X1 U539 ( .A(G472), .ZN(n458) );
  INV_X1 U540 ( .A(G107), .ZN(n574) );
  XOR2_X1 U541 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n587) );
  NAND2_X1 U542 ( .A1(n519), .A2(n376), .ZN(n595) );
  INV_X1 U543 ( .A(n746), .ZN(n467) );
  INV_X1 U544 ( .A(KEYINPUT70), .ZN(n401) );
  NAND2_X1 U545 ( .A1(n405), .A2(n403), .ZN(n402) );
  AND2_X1 U546 ( .A1(n404), .A2(n512), .ZN(n403) );
  BUF_X1 U547 ( .A(n741), .Z(n486) );
  OR2_X1 U548 ( .A1(n508), .A2(n503), .ZN(n502) );
  XNOR2_X1 U549 ( .A(n530), .B(n433), .ZN(n432) );
  XNOR2_X1 U550 ( .A(n532), .B(n531), .ZN(n530) );
  XNOR2_X1 U551 ( .A(n618), .B(n485), .ZN(n781) );
  XNOR2_X1 U552 ( .A(n619), .B(n620), .ZN(n485) );
  INV_X1 U553 ( .A(KEYINPUT42), .ZN(n399) );
  NOR2_X1 U554 ( .A1(n672), .A2(n382), .ZN(n394) );
  NOR2_X1 U555 ( .A1(n683), .A2(n681), .ZN(n668) );
  XNOR2_X1 U556 ( .A(KEYINPUT73), .B(KEYINPUT32), .ZN(n525) );
  XOR2_X1 U557 ( .A(KEYINPUT110), .B(n672), .Z(n718) );
  NAND2_X1 U558 ( .A1(n387), .A2(n737), .ZN(n704) );
  XNOR2_X1 U559 ( .A(n785), .B(KEYINPUT122), .ZN(n465) );
  XNOR2_X1 U560 ( .A(n777), .B(n490), .ZN(n780) );
  XNOR2_X1 U561 ( .A(n487), .B(n778), .ZN(n490) );
  AND2_X1 U562 ( .A1(n522), .A2(n521), .ZN(n376) );
  OR2_X1 U563 ( .A1(n374), .A2(n502), .ZN(n377) );
  AND2_X1 U564 ( .A1(n754), .A2(KEYINPUT47), .ZN(n378) );
  INV_X1 U565 ( .A(n512), .ZN(n429) );
  INV_X1 U566 ( .A(n688), .ZN(n687) );
  OR2_X1 U567 ( .A1(n661), .A2(KEYINPUT47), .ZN(n379) );
  AND2_X1 U568 ( .A1(n592), .A2(n688), .ZN(n380) );
  AND2_X1 U569 ( .A1(n709), .A2(KEYINPUT106), .ZN(n381) );
  XOR2_X1 U570 ( .A(KEYINPUT112), .B(KEYINPUT40), .Z(n382) );
  XOR2_X1 U571 ( .A(KEYINPUT0), .B(KEYINPUT88), .Z(n383) );
  INV_X1 U572 ( .A(KEYINPUT107), .ZN(n495) );
  INV_X1 U573 ( .A(KEYINPUT87), .ZN(n517) );
  NAND2_X1 U574 ( .A1(n387), .A2(n385), .ZN(n468) );
  INV_X1 U575 ( .A(n737), .ZN(n386) );
  BUF_X1 U576 ( .A(n763), .Z(n389) );
  XNOR2_X1 U577 ( .A(n676), .B(n675), .ZN(n763) );
  XNOR2_X1 U578 ( .A(n368), .B(G128), .ZN(n598) );
  AND2_X2 U579 ( .A1(n527), .A2(n686), .ZN(n694) );
  NAND2_X1 U580 ( .A1(n630), .A2(n629), .ZN(n672) );
  BUF_X2 U581 ( .A(n734), .Z(n489) );
  NAND2_X1 U582 ( .A1(n498), .A2(n496), .ZN(n391) );
  NAND2_X1 U583 ( .A1(n498), .A2(n496), .ZN(n662) );
  BUF_X1 U584 ( .A(n597), .Z(n392) );
  NAND2_X1 U585 ( .A1(n694), .A2(n687), .ZN(n452) );
  AND2_X1 U586 ( .A1(n391), .A2(n650), .ZN(n651) );
  NAND2_X1 U587 ( .A1(n680), .A2(n382), .ZN(n398) );
  INV_X1 U588 ( .A(n680), .ZN(n395) );
  NAND2_X1 U589 ( .A1(n477), .A2(n514), .ZN(n408) );
  XNOR2_X1 U590 ( .A(n444), .B(n384), .ZN(n693) );
  INV_X1 U591 ( .A(n536), .ZN(n412) );
  NAND2_X1 U592 ( .A1(n416), .A2(n414), .ZN(n413) );
  NAND2_X1 U593 ( .A1(n418), .A2(n415), .ZN(n414) );
  INV_X1 U594 ( .A(n657), .ZN(n428) );
  OR2_X1 U595 ( .A1(n430), .A2(n429), .ZN(n677) );
  NOR2_X1 U596 ( .A1(n657), .A2(n421), .ZN(n420) );
  INV_X1 U597 ( .A(n430), .ZN(n422) );
  NAND2_X1 U598 ( .A1(n430), .A2(n426), .ZN(n424) );
  NAND2_X1 U599 ( .A1(n428), .A2(n512), .ZN(n427) );
  XNOR2_X1 U600 ( .A(n484), .B(n431), .ZN(n430) );
  INV_X1 U601 ( .A(KEYINPUT28), .ZN(n431) );
  NAND2_X1 U602 ( .A1(n438), .A2(n437), .ZN(n436) );
  INV_X1 U603 ( .A(n709), .ZN(n438) );
  XNOR2_X1 U604 ( .A(n439), .B(n565), .ZN(n697) );
  XNOR2_X2 U605 ( .A(n804), .B(n550), .ZN(n439) );
  XNOR2_X2 U606 ( .A(n442), .B(n578), .ZN(n798) );
  XNOR2_X2 U607 ( .A(n443), .B(n617), .ZN(n442) );
  XNOR2_X2 U608 ( .A(n597), .B(n479), .ZN(n443) );
  NAND2_X2 U609 ( .A1(n577), .A2(n576), .ZN(n597) );
  NAND2_X1 U610 ( .A1(n447), .A2(n445), .ZN(n444) );
  XNOR2_X1 U611 ( .A(n644), .B(n446), .ZN(n445) );
  XNOR2_X1 U612 ( .A(n448), .B(n459), .ZN(n447) );
  NAND2_X1 U613 ( .A1(n471), .A2(n470), .ZN(n448) );
  XNOR2_X1 U614 ( .A(n463), .B(n462), .ZN(n461) );
  INV_X1 U615 ( .A(n741), .ZN(n655) );
  NAND2_X1 U616 ( .A1(n670), .A2(n750), .ZN(n451) );
  OR2_X2 U617 ( .A1(n693), .A2(n452), .ZN(n691) );
  INV_X1 U618 ( .A(n694), .ZN(n805) );
  XNOR2_X1 U619 ( .A(n741), .B(KEYINPUT6), .ZN(n523) );
  XNOR2_X2 U620 ( .A(n566), .B(n458), .ZN(n741) );
  NOR2_X1 U621 ( .A1(n464), .A2(n790), .ZN(G63) );
  XNOR2_X1 U622 ( .A(n466), .B(n465), .ZN(n464) );
  NAND2_X1 U623 ( .A1(n786), .A2(G478), .ZN(n466) );
  NAND2_X1 U624 ( .A1(n469), .A2(n468), .ZN(n472) );
  NAND2_X1 U625 ( .A1(n492), .A2(n704), .ZN(n469) );
  NAND2_X1 U626 ( .A1(n641), .A2(KEYINPUT87), .ZN(n473) );
  XNOR2_X1 U627 ( .A(n598), .B(n474), .ZN(n602) );
  NAND2_X1 U628 ( .A1(n656), .A2(n594), .ZN(n476) );
  XNOR2_X2 U629 ( .A(n624), .B(n623), .ZN(n639) );
  XNOR2_X2 U630 ( .A(n482), .B(KEYINPUT19), .ZN(n656) );
  XNOR2_X2 U631 ( .A(G110), .B(KEYINPUT16), .ZN(n479) );
  BUF_X1 U632 ( .A(n723), .Z(n480) );
  NAND2_X1 U633 ( .A1(n494), .A2(n495), .ZN(n493) );
  XNOR2_X2 U634 ( .A(n481), .B(n591), .ZN(n773) );
  NAND2_X1 U635 ( .A1(n582), .A2(n583), .ZN(n481) );
  NAND2_X1 U636 ( .A1(n662), .A2(n749), .ZN(n482) );
  INV_X1 U637 ( .A(n798), .ZN(n581) );
  NOR2_X1 U638 ( .A1(n788), .A2(G902), .ZN(n538) );
  NOR2_X2 U639 ( .A1(n630), .A2(n629), .ZN(n713) );
  XOR2_X2 U640 ( .A(G146), .B(G125), .Z(n580) );
  NAND2_X1 U641 ( .A1(n488), .A2(n650), .ZN(n624) );
  XNOR2_X1 U642 ( .A(n595), .B(n596), .ZN(n488) );
  INV_X1 U643 ( .A(n634), .ZN(n494) );
  INV_X1 U644 ( .A(n773), .ZN(n497) );
  AND2_X2 U645 ( .A1(n500), .A2(n499), .ZN(n498) );
  NAND2_X1 U646 ( .A1(n773), .A2(n501), .ZN(n500) );
  INV_X1 U647 ( .A(n592), .ZN(n501) );
  OR2_X1 U648 ( .A1(n374), .A2(n489), .ZN(n509) );
  INV_X1 U649 ( .A(n489), .ZN(n504) );
  OR2_X1 U650 ( .A1(n508), .A2(n489), .ZN(n506) );
  INV_X1 U651 ( .A(n509), .ZN(n638) );
  INV_X1 U652 ( .A(KEYINPUT85), .ZN(n507) );
  INV_X1 U653 ( .A(n523), .ZN(n508) );
  XNOR2_X2 U654 ( .A(n585), .B(n549), .ZN(n804) );
  XNOR2_X2 U655 ( .A(n390), .B(n510), .ZN(n585) );
  NAND2_X1 U656 ( .A1(n735), .A2(n512), .ZN(n632) );
  XNOR2_X2 U657 ( .A(n556), .B(n524), .ZN(n513) );
  NAND2_X1 U658 ( .A1(n639), .A2(n515), .ZN(n514) );
  NAND2_X1 U659 ( .A1(n376), .A2(n520), .ZN(n764) );
  NAND2_X1 U660 ( .A1(n523), .A2(n567), .ZN(n521) );
  NAND2_X1 U661 ( .A1(n557), .A2(n567), .ZN(n522) );
  NOR2_X2 U662 ( .A1(n636), .A2(n635), .ZN(n526) );
  XNOR2_X1 U663 ( .A(n678), .B(KEYINPUT46), .ZN(n529) );
  INV_X1 U664 ( .A(KEYINPUT77), .ZN(n535) );
  XNOR2_X1 U665 ( .A(KEYINPUT59), .B(KEYINPUT89), .ZN(n539) );
  NAND2_X1 U666 ( .A1(n641), .A2(n640), .ZN(n642) );
  INV_X1 U667 ( .A(n728), .ZN(n685) );
  INV_X1 U668 ( .A(KEYINPUT33), .ZN(n567) );
  XNOR2_X1 U669 ( .A(n578), .B(n562), .ZN(n563) );
  XNOR2_X1 U670 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U671 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U672 ( .A(n552), .B(n616), .ZN(n553) );
  INV_X1 U673 ( .A(KEYINPUT63), .ZN(n701) );
  XNOR2_X1 U674 ( .A(n701), .B(KEYINPUT90), .ZN(n702) );
  XOR2_X1 U675 ( .A(KEYINPUT34), .B(KEYINPUT72), .Z(n596) );
  NAND2_X1 U676 ( .A1(G234), .A2(n688), .ZN(n540) );
  XNOR2_X1 U677 ( .A(KEYINPUT20), .B(n540), .ZN(n546) );
  NAND2_X1 U678 ( .A1(n546), .A2(G221), .ZN(n541) );
  XOR2_X1 U679 ( .A(KEYINPUT21), .B(n541), .Z(n738) );
  INV_X1 U680 ( .A(n738), .ZN(n626) );
  INV_X1 U681 ( .A(KEYINPUT25), .ZN(n548) );
  INV_X1 U682 ( .A(n615), .ZN(n545) );
  NAND2_X1 U683 ( .A1(G234), .A2(n806), .ZN(n542) );
  XNOR2_X1 U684 ( .A(n543), .B(n542), .ZN(n603) );
  NAND2_X1 U685 ( .A1(G221), .A2(n603), .ZN(n544) );
  NAND2_X1 U686 ( .A1(n546), .A2(G217), .ZN(n547) );
  XOR2_X1 U687 ( .A(n349), .B(n584), .Z(n550) );
  NAND2_X1 U688 ( .A1(G227), .A2(n806), .ZN(n551) );
  XNOR2_X1 U689 ( .A(n554), .B(n553), .ZN(n555) );
  NOR2_X2 U690 ( .A1(n779), .A2(G902), .ZN(n556) );
  NAND2_X1 U691 ( .A1(n611), .A2(G210), .ZN(n559) );
  XNOR2_X1 U692 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U693 ( .A(n560), .B(KEYINPUT5), .Z(n564) );
  XNOR2_X1 U694 ( .A(KEYINPUT91), .B(KEYINPUT3), .ZN(n561) );
  NAND2_X1 U695 ( .A1(G234), .A2(G237), .ZN(n568) );
  XNOR2_X1 U696 ( .A(n568), .B(KEYINPUT14), .ZN(n570) );
  NAND2_X1 U697 ( .A1(G952), .A2(n570), .ZN(n762) );
  NOR2_X1 U698 ( .A1(n762), .A2(G953), .ZN(n569) );
  XNOR2_X1 U699 ( .A(n569), .B(KEYINPUT93), .ZN(n647) );
  NOR2_X1 U700 ( .A1(G898), .A2(n806), .ZN(n800) );
  NAND2_X1 U701 ( .A1(G902), .A2(n570), .ZN(n645) );
  INV_X1 U702 ( .A(n645), .ZN(n571) );
  NAND2_X1 U703 ( .A1(n800), .A2(n571), .ZN(n572) );
  NAND2_X1 U704 ( .A1(n647), .A2(n572), .ZN(n573) );
  XNOR2_X1 U705 ( .A(KEYINPUT94), .B(n573), .ZN(n594) );
  NAND2_X1 U706 ( .A1(n574), .A2(G116), .ZN(n577) );
  NAND2_X1 U707 ( .A1(n575), .A2(G107), .ZN(n576) );
  INV_X1 U708 ( .A(n580), .ZN(n579) );
  NAND2_X1 U709 ( .A1(n798), .A2(n579), .ZN(n583) );
  NAND2_X1 U710 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U711 ( .A(n585), .B(n584), .ZN(n590) );
  NAND2_X1 U712 ( .A1(G224), .A2(n806), .ZN(n586) );
  XNOR2_X1 U713 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U714 ( .A(KEYINPUT92), .B(n588), .ZN(n589) );
  NAND2_X1 U715 ( .A1(G210), .A2(n593), .ZN(n592) );
  XNOR2_X1 U716 ( .A(KEYINPUT104), .B(G478), .ZN(n608) );
  XNOR2_X1 U717 ( .A(n392), .B(G134), .ZN(n606) );
  XNOR2_X1 U718 ( .A(n600), .B(n599), .ZN(n601) );
  XOR2_X1 U719 ( .A(n602), .B(n601), .Z(n605) );
  NAND2_X1 U720 ( .A1(G217), .A2(n603), .ZN(n604) );
  NOR2_X1 U721 ( .A1(G902), .A2(n785), .ZN(n607) );
  XOR2_X1 U722 ( .A(KEYINPUT11), .B(KEYINPUT99), .Z(n610) );
  XNOR2_X1 U723 ( .A(n610), .B(n609), .ZN(n620) );
  NAND2_X1 U724 ( .A1(G214), .A2(n611), .ZN(n612) );
  XOR2_X1 U725 ( .A(n614), .B(KEYINPUT12), .Z(n619) );
  XNOR2_X1 U726 ( .A(n803), .B(n617), .ZN(n618) );
  XNOR2_X1 U727 ( .A(KEYINPUT13), .B(G475), .ZN(n621) );
  INV_X1 U728 ( .A(n630), .ZN(n625) );
  NOR2_X1 U729 ( .A1(n629), .A2(n625), .ZN(n650) );
  XOR2_X1 U730 ( .A(KEYINPUT35), .B(KEYINPUT71), .Z(n623) );
  NAND2_X1 U731 ( .A1(n629), .A2(n625), .ZN(n752) );
  NOR2_X1 U732 ( .A1(n752), .A2(n626), .ZN(n627) );
  INV_X1 U733 ( .A(n664), .ZN(n737) );
  NOR2_X1 U734 ( .A1(n486), .A2(n632), .ZN(n633) );
  NOR2_X1 U735 ( .A1(n486), .A2(n737), .ZN(n637) );
  NAND2_X1 U736 ( .A1(n638), .A2(n637), .ZN(n712) );
  INV_X1 U737 ( .A(KEYINPUT44), .ZN(n640) );
  NOR2_X1 U738 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U739 ( .A1(G900), .A2(n645), .ZN(n646) );
  NAND2_X1 U740 ( .A1(G953), .A2(n646), .ZN(n648) );
  NAND2_X1 U741 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U742 ( .A1(n649), .A2(n738), .ZN(n653) );
  NAND2_X1 U743 ( .A1(n670), .A2(n651), .ZN(n652) );
  XNOR2_X1 U744 ( .A(KEYINPUT67), .B(n653), .ZN(n663) );
  NAND2_X1 U745 ( .A1(n664), .A2(n663), .ZN(n654) );
  INV_X1 U746 ( .A(n656), .ZN(n657) );
  NAND2_X1 U747 ( .A1(n659), .A2(KEYINPUT47), .ZN(n658) );
  INV_X1 U748 ( .A(n659), .ZN(n717) );
  NAND2_X1 U749 ( .A1(n717), .A2(n660), .ZN(n661) );
  NAND2_X1 U750 ( .A1(n663), .A2(n749), .ZN(n666) );
  NAND2_X1 U751 ( .A1(n664), .A2(n718), .ZN(n665) );
  NOR2_X1 U752 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U753 ( .A1(n508), .A2(n667), .ZN(n681) );
  XNOR2_X1 U754 ( .A(n668), .B(KEYINPUT36), .ZN(n669) );
  NAND2_X1 U755 ( .A1(n669), .A2(n489), .ZN(n727) );
  XNOR2_X2 U756 ( .A(n683), .B(KEYINPUT38), .ZN(n750) );
  XOR2_X1 U757 ( .A(KEYINPUT84), .B(KEYINPUT39), .Z(n671) );
  NAND2_X1 U758 ( .A1(n750), .A2(n749), .ZN(n753) );
  XNOR2_X1 U759 ( .A(KEYINPUT114), .B(KEYINPUT41), .ZN(n674) );
  NOR2_X1 U760 ( .A1(n680), .A2(n679), .ZN(n728) );
  OR2_X1 U761 ( .A1(n489), .A2(n681), .ZN(n682) );
  XNOR2_X1 U762 ( .A(n682), .B(KEYINPUT43), .ZN(n684) );
  NAND2_X1 U763 ( .A1(n684), .A2(n683), .ZN(n730) );
  XNOR2_X1 U764 ( .A(n688), .B(KEYINPUT81), .ZN(n689) );
  NAND2_X1 U765 ( .A1(n689), .A2(KEYINPUT2), .ZN(n690) );
  INV_X1 U766 ( .A(KEYINPUT64), .ZN(n692) );
  BUF_X1 U767 ( .A(n693), .Z(n795) );
  NAND2_X1 U768 ( .A1(n694), .A2(KEYINPUT2), .ZN(n695) );
  NOR2_X4 U769 ( .A1(n696), .A2(n733), .ZN(n786) );
  NAND2_X1 U770 ( .A1(n786), .A2(G472), .ZN(n699) );
  XNOR2_X1 U771 ( .A(n699), .B(n698), .ZN(n700) );
  XNOR2_X1 U772 ( .A(n703), .B(n702), .ZN(G57) );
  XNOR2_X1 U773 ( .A(n375), .B(G101), .ZN(G3) );
  INV_X1 U774 ( .A(n718), .ZN(n720) );
  NOR2_X1 U775 ( .A1(n720), .A2(n709), .ZN(n706) );
  XNOR2_X1 U776 ( .A(G104), .B(KEYINPUT115), .ZN(n705) );
  XNOR2_X1 U777 ( .A(n706), .B(n705), .ZN(G6) );
  XOR2_X1 U778 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n708) );
  XNOR2_X1 U779 ( .A(G107), .B(KEYINPUT116), .ZN(n707) );
  XNOR2_X1 U780 ( .A(n708), .B(n707), .ZN(n711) );
  INV_X1 U781 ( .A(n713), .ZN(n724) );
  NOR2_X1 U782 ( .A1(n724), .A2(n709), .ZN(n710) );
  XOR2_X1 U783 ( .A(n711), .B(n710), .Z(G9) );
  XNOR2_X1 U784 ( .A(G110), .B(n712), .ZN(G12) );
  XOR2_X1 U785 ( .A(KEYINPUT117), .B(KEYINPUT29), .Z(n715) );
  NAND2_X1 U786 ( .A1(n717), .A2(n713), .ZN(n714) );
  XNOR2_X1 U787 ( .A(n715), .B(n714), .ZN(n716) );
  XOR2_X1 U788 ( .A(G128), .B(n716), .Z(G30) );
  NAND2_X1 U789 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U790 ( .A(n719), .B(n349), .ZN(G48) );
  NOR2_X1 U791 ( .A1(n720), .A2(n480), .ZN(n721) );
  XOR2_X1 U792 ( .A(KEYINPUT118), .B(n721), .Z(n722) );
  XNOR2_X1 U793 ( .A(G113), .B(n722), .ZN(G15) );
  NOR2_X1 U794 ( .A1(n724), .A2(n480), .ZN(n725) );
  XOR2_X1 U795 ( .A(n475), .B(n725), .Z(G18) );
  XOR2_X1 U796 ( .A(G125), .B(KEYINPUT37), .Z(n726) );
  XNOR2_X1 U797 ( .A(n727), .B(n726), .ZN(G27) );
  XOR2_X1 U798 ( .A(G134), .B(n728), .Z(G36) );
  XOR2_X1 U799 ( .A(G140), .B(KEYINPUT119), .Z(n729) );
  XNOR2_X1 U800 ( .A(n730), .B(n729), .ZN(G42) );
  XNOR2_X1 U801 ( .A(KEYINPUT76), .B(KEYINPUT2), .ZN(n731) );
  NOR2_X1 U802 ( .A1(n453), .A2(n731), .ZN(n732) );
  NOR2_X1 U803 ( .A1(n733), .A2(n732), .ZN(n770) );
  NOR2_X1 U804 ( .A1(n735), .A2(n489), .ZN(n736) );
  XOR2_X1 U805 ( .A(KEYINPUT50), .B(n736), .Z(n744) );
  NOR2_X1 U806 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U807 ( .A(KEYINPUT49), .B(n739), .Z(n740) );
  NOR2_X1 U808 ( .A1(n486), .A2(n740), .ZN(n742) );
  XNOR2_X1 U809 ( .A(KEYINPUT120), .B(n742), .ZN(n743) );
  NAND2_X1 U810 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U811 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U812 ( .A(KEYINPUT51), .B(n747), .ZN(n748) );
  NOR2_X1 U813 ( .A1(n389), .A2(n748), .ZN(n759) );
  NOR2_X1 U814 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U815 ( .A1(n752), .A2(n751), .ZN(n756) );
  NOR2_X1 U816 ( .A1(n754), .A2(n753), .ZN(n755) );
  NOR2_X1 U817 ( .A1(n756), .A2(n755), .ZN(n757) );
  NOR2_X1 U818 ( .A1(n757), .A2(n764), .ZN(n758) );
  NOR2_X1 U819 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U820 ( .A(n760), .B(KEYINPUT52), .ZN(n761) );
  NOR2_X1 U821 ( .A1(n762), .A2(n761), .ZN(n766) );
  NOR2_X1 U822 ( .A1(n764), .A2(n389), .ZN(n765) );
  NOR2_X1 U823 ( .A1(n766), .A2(n765), .ZN(n767) );
  XOR2_X1 U824 ( .A(KEYINPUT121), .B(n767), .Z(n768) );
  NAND2_X1 U825 ( .A1(n768), .A2(n806), .ZN(n769) );
  NOR2_X1 U826 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U827 ( .A(KEYINPUT53), .B(n771), .ZN(G75) );
  NAND2_X1 U828 ( .A1(n786), .A2(G210), .ZN(n775) );
  XOR2_X1 U829 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n772) );
  XNOR2_X1 U830 ( .A(n773), .B(n772), .ZN(n774) );
  XNOR2_X1 U831 ( .A(n775), .B(n774), .ZN(n776) );
  XOR2_X1 U832 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n778) );
  NAND2_X1 U833 ( .A1(n786), .A2(G469), .ZN(n777) );
  NOR2_X1 U834 ( .A1(n790), .A2(n780), .ZN(G54) );
  NAND2_X1 U835 ( .A1(n786), .A2(G475), .ZN(n783) );
  XNOR2_X1 U836 ( .A(n783), .B(n782), .ZN(n784) );
  NAND2_X1 U837 ( .A1(G217), .A2(n786), .ZN(n787) );
  XNOR2_X1 U838 ( .A(n788), .B(n787), .ZN(n789) );
  NOR2_X1 U839 ( .A1(n790), .A2(n789), .ZN(G66) );
  XOR2_X1 U840 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n792) );
  NAND2_X1 U841 ( .A1(G224), .A2(G953), .ZN(n791) );
  XNOR2_X1 U842 ( .A(n792), .B(n791), .ZN(n793) );
  NAND2_X1 U843 ( .A1(G898), .A2(n793), .ZN(n794) );
  XOR2_X1 U844 ( .A(KEYINPUT124), .B(n794), .Z(n797) );
  NOR2_X1 U845 ( .A1(G953), .A2(n795), .ZN(n796) );
  NOR2_X1 U846 ( .A1(n797), .A2(n796), .ZN(n802) );
  XNOR2_X1 U847 ( .A(G101), .B(n373), .ZN(n799) );
  NOR2_X1 U848 ( .A1(n800), .A2(n799), .ZN(n801) );
  XOR2_X1 U849 ( .A(n802), .B(n801), .Z(G69) );
  XOR2_X1 U850 ( .A(n804), .B(n803), .Z(n808) );
  XNOR2_X1 U851 ( .A(n805), .B(n808), .ZN(n807) );
  NAND2_X1 U852 ( .A1(n807), .A2(n806), .ZN(n813) );
  XNOR2_X1 U853 ( .A(G227), .B(n808), .ZN(n809) );
  NAND2_X1 U854 ( .A1(n809), .A2(G900), .ZN(n810) );
  NAND2_X1 U855 ( .A1(G953), .A2(n810), .ZN(n811) );
  XOR2_X1 U856 ( .A(KEYINPUT125), .B(n811), .Z(n812) );
  NAND2_X1 U857 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U858 ( .A(KEYINPUT126), .B(n814), .ZN(G72) );
  XOR2_X1 U859 ( .A(n815), .B(G131), .Z(G33) );
  XNOR2_X1 U860 ( .A(n639), .B(G122), .ZN(n816) );
  XNOR2_X1 U861 ( .A(n816), .B(KEYINPUT127), .ZN(G24) );
  XOR2_X1 U862 ( .A(n817), .B(n478), .Z(G45) );
  XOR2_X1 U863 ( .A(n818), .B(G137), .Z(G39) );
endmodule

