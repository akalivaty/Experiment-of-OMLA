//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 0 0 1 1 1 1 1 0 0 0 1 0 1 1 1 1 0 1 0 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT64), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT65), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n209), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n212), .B(new_n219), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT67), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n240), .B(KEYINPUT68), .Z(new_n241));
  XOR2_X1   g0041(.A(G50), .B(G58), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT66), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G68), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G351));
  OR2_X1    g0046(.A1(KEYINPUT3), .A2(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  AOI21_X1  g0048(.A(G1698), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G222), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n247), .A2(new_n248), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G223), .A3(G1698), .ZN(new_n252));
  AND2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G77), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n250), .A2(new_n252), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(KEYINPUT70), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT70), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n250), .A2(new_n252), .A3(new_n259), .A4(new_n256), .ZN(new_n260));
  AND2_X1   g0060(.A1(G1), .A2(G13), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT71), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G33), .A2(G41), .ZN(new_n263));
  AND3_X1   g0063(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n262), .B1(new_n261), .B2(new_n263), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n258), .A2(new_n260), .A3(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n263), .A2(G1), .A3(G13), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n269), .A2(new_n270), .A3(G274), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT69), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n273), .B1(new_n270), .B2(new_n268), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n270), .A2(new_n273), .A3(new_n268), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n272), .B1(new_n277), .B2(G226), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n267), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(G169), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n213), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n207), .A2(G33), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT8), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G58), .ZN(new_n286));
  XNOR2_X1  g0086(.A(new_n286), .B(KEYINPUT73), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT72), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n202), .A2(KEYINPUT72), .A3(KEYINPUT8), .ZN(new_n291));
  AND2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n284), .B1(new_n287), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n294));
  INV_X1    g0094(.A(G33), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n207), .A2(new_n295), .A3(KEYINPUT74), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT74), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n297), .B1(G20), .B2(G33), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G150), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n294), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n283), .B1(new_n293), .B2(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n207), .A2(G1), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT75), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n304), .B1(new_n306), .B2(new_n283), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n305), .A2(KEYINPUT75), .A3(new_n213), .A4(new_n282), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n303), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G50), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n306), .A2(new_n201), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n302), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n279), .A2(G179), .ZN(new_n314));
  NOR3_X1   g0114(.A1(new_n281), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G200), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(new_n267), .B2(new_n278), .ZN(new_n317));
  OAI21_X1  g0117(.A(KEYINPUT10), .B1(new_n317), .B2(KEYINPUT79), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n302), .A2(KEYINPUT9), .A3(new_n310), .A4(new_n311), .ZN(new_n320));
  XNOR2_X1  g0120(.A(new_n320), .B(KEYINPUT78), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT9), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n312), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n267), .A2(G190), .A3(new_n278), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n323), .B(new_n324), .C1(new_n280), .C2(new_n316), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n319), .B1(new_n321), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT78), .ZN(new_n327));
  XNOR2_X1  g0127(.A(new_n320), .B(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n317), .B1(new_n322), .B2(new_n312), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n328), .A2(new_n318), .A3(new_n324), .A4(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n315), .B1(new_n326), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n277), .A2(G244), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n332), .A2(KEYINPUT76), .A3(new_n271), .ZN(new_n333));
  INV_X1    g0133(.A(G1698), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n251), .A2(G232), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n251), .A2(G238), .A3(G1698), .ZN(new_n336));
  INV_X1    g0136(.A(G107), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n335), .B(new_n336), .C1(new_n337), .C2(new_n251), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n266), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT76), .ZN(new_n340));
  INV_X1    g0140(.A(G244), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n341), .B1(new_n275), .B2(new_n276), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n340), .B1(new_n342), .B2(new_n272), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n333), .A2(new_n339), .A3(new_n343), .ZN(new_n344));
  OR2_X1    g0144(.A1(new_n344), .A2(G179), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n296), .A2(new_n298), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n286), .A2(new_n288), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g0148(.A(KEYINPUT15), .B(G87), .ZN(new_n349));
  INV_X1    g0149(.A(G77), .ZN(new_n350));
  OAI22_X1  g0150(.A1(new_n349), .A2(new_n284), .B1(new_n207), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n283), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n306), .A2(new_n283), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n303), .A2(new_n350), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n353), .A2(new_n354), .B1(new_n350), .B2(new_n306), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G169), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n344), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n345), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n356), .B1(new_n344), .B2(G200), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n361), .A2(KEYINPUT77), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G190), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n344), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n365), .B1(new_n361), .B2(KEYINPUT77), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n360), .B1(new_n363), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n331), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT80), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT80), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n331), .A2(new_n367), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT87), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT16), .ZN(new_n373));
  INV_X1    g0173(.A(G68), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n247), .A2(new_n207), .A3(new_n248), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT7), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n247), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n248), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n374), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  XNOR2_X1  g0179(.A(G58), .B(G68), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(G20), .ZN(new_n381));
  INV_X1    g0181(.A(G159), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n381), .B1(new_n299), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n373), .B1(new_n379), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT7), .B1(new_n255), .B2(new_n207), .ZN(new_n385));
  NOR4_X1   g0185(.A1(new_n253), .A2(new_n254), .A3(new_n376), .A4(G20), .ZN(new_n386));
  OAI21_X1  g0186(.A(G68), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n346), .A2(G159), .B1(new_n380), .B2(G20), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n387), .A2(KEYINPUT16), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n384), .A2(new_n389), .A3(new_n283), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT85), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n287), .A2(new_n292), .A3(new_n305), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT73), .ZN(new_n393));
  XNOR2_X1  g0193(.A(new_n286), .B(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n290), .A2(new_n291), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n392), .B1(new_n309), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT86), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT86), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n399), .B(new_n392), .C1(new_n309), .C2(new_n396), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT85), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n384), .A2(new_n389), .A3(new_n402), .A4(new_n283), .ZN(new_n403));
  INV_X1    g0203(.A(G232), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n270), .A2(new_n268), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n271), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  OR2_X1    g0207(.A1(G223), .A2(G1698), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(G226), .B2(new_n334), .ZN(new_n409));
  INV_X1    g0209(.A(G87), .ZN(new_n410));
  OAI22_X1  g0210(.A1(new_n409), .A2(new_n255), .B1(new_n295), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n266), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n407), .A2(new_n364), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n406), .B1(new_n411), .B2(new_n266), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n413), .B1(new_n414), .B2(G200), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n391), .A2(new_n401), .A3(new_n403), .A4(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT17), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n416), .A2(new_n417), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n372), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n391), .A2(new_n401), .A3(new_n403), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT18), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n414), .A2(G179), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(new_n357), .B2(new_n414), .ZN(new_n424));
  AND3_X1   g0224(.A1(new_n421), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n422), .B1(new_n421), .B2(new_n424), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n391), .A2(new_n403), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n428), .A2(KEYINPUT17), .A3(new_n401), .A4(new_n415), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n416), .A2(new_n417), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n429), .A2(KEYINPUT87), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n420), .A2(new_n427), .A3(new_n431), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n369), .A2(new_n371), .B1(KEYINPUT88), .B2(new_n432), .ZN(new_n433));
  OR2_X1    g0233(.A1(new_n432), .A2(KEYINPUT88), .ZN(new_n434));
  OAI211_X1 g0234(.A(G232), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n435));
  OAI211_X1 g0235(.A(G226), .B(new_n334), .C1(new_n253), .C2(new_n254), .ZN(new_n436));
  NAND2_X1  g0236(.A1(G33), .A2(G97), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n266), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n270), .A2(new_n273), .A3(new_n268), .ZN(new_n440));
  OAI21_X1  g0240(.A(G238), .B1(new_n440), .B2(new_n274), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT13), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n439), .A2(new_n441), .A3(new_n442), .A4(new_n271), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(G179), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n439), .A2(new_n441), .A3(new_n271), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT81), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n442), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT82), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n439), .A2(new_n441), .A3(KEYINPUT81), .A4(new_n271), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n450), .B1(new_n449), .B2(new_n451), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n446), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT14), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n447), .A2(KEYINPUT13), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n443), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n455), .B1(new_n457), .B2(G169), .ZN(new_n458));
  AOI211_X1 g0258(.A(KEYINPUT14), .B(new_n357), .C1(new_n456), .C2(new_n443), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n454), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n299), .A2(new_n201), .ZN(new_n462));
  OAI22_X1  g0262(.A1(new_n284), .A2(new_n350), .B1(new_n207), .B2(G68), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n283), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT11), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT12), .B1(new_n305), .B2(G68), .ZN(new_n467));
  OR3_X1    g0267(.A1(new_n305), .A2(KEYINPUT12), .A3(G68), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n303), .A2(new_n374), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n467), .A2(new_n468), .B1(new_n353), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n470), .B1(new_n464), .B2(new_n465), .ZN(new_n471));
  OR2_X1    g0271(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n461), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n444), .A2(new_n364), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n447), .A2(new_n448), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n476), .A2(KEYINPUT13), .A3(new_n451), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(KEYINPUT82), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n475), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n457), .A2(G200), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n466), .A2(new_n471), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR3_X1   g0283(.A1(new_n480), .A2(KEYINPUT83), .A3(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT83), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n474), .B1(new_n452), .B2(new_n453), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n472), .B1(G200), .B2(new_n457), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n473), .B1(new_n484), .B2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT84), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n473), .B(KEYINPUT84), .C1(new_n488), .C2(new_n484), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n433), .A2(new_n434), .A3(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(G107), .B1(new_n385), .B2(new_n386), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT91), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g0297(.A(KEYINPUT91), .B(G107), .C1(new_n385), .C2(new_n386), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n337), .A2(KEYINPUT6), .A3(G97), .ZN(new_n499));
  OR2_X1    g0299(.A1(new_n499), .A2(KEYINPUT90), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(KEYINPUT90), .ZN(new_n501));
  INV_X1    g0301(.A(G97), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n502), .A2(new_n337), .ZN(new_n503));
  NOR2_X1   g0303(.A1(G97), .A2(G107), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n500), .B(new_n501), .C1(KEYINPUT6), .C2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G20), .ZN(new_n507));
  AND3_X1   g0307(.A1(new_n346), .A2(KEYINPUT89), .A3(G77), .ZN(new_n508));
  AOI21_X1  g0308(.A(KEYINPUT89), .B1(new_n346), .B2(G77), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n497), .A2(new_n498), .A3(new_n507), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n283), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n305), .A2(G97), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n206), .A2(G33), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n353), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n513), .B1(new_n516), .B2(G97), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT92), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT5), .ZN(new_n520));
  INV_X1    g0320(.A(G41), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(KEYINPUT5), .A2(G41), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(G45), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n525), .A2(G1), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n524), .A2(new_n526), .B1(new_n261), .B2(new_n263), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G257), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n206), .A2(G45), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n529), .B1(new_n522), .B2(new_n523), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n530), .A2(G274), .A3(new_n270), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(G250), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT94), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n251), .A2(KEYINPUT94), .A3(G250), .A4(G1698), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(G244), .B(new_n334), .C1(new_n253), .C2(new_n254), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT4), .ZN(new_n539));
  OAI21_X1  g0339(.A(KEYINPUT93), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n538), .A2(new_n539), .B1(G33), .B2(G283), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT93), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n249), .A2(new_n542), .A3(KEYINPUT4), .A4(G244), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n537), .A2(new_n540), .A3(new_n541), .A4(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n532), .B1(new_n544), .B2(new_n266), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n364), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(G200), .B2(new_n545), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT92), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n512), .A2(new_n548), .A3(new_n517), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n519), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  AND2_X1   g0350(.A1(new_n545), .A2(G179), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n545), .A2(new_n357), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n518), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n283), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n251), .A2(new_n207), .A3(G68), .ZN(new_n555));
  XNOR2_X1  g0355(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(new_n502), .B2(new_n284), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n207), .B1(new_n556), .B2(new_n437), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n504), .A2(new_n410), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n554), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n515), .A2(new_n410), .ZN(new_n563));
  INV_X1    g0363(.A(new_n349), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n564), .A2(new_n305), .ZN(new_n565));
  NOR3_X1   g0365(.A1(new_n562), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n251), .A2(G244), .A3(G1698), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n251), .A2(G238), .A3(new_n334), .ZN(new_n568));
  INV_X1    g0368(.A(G116), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n295), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n567), .A2(new_n568), .A3(new_n571), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n572), .A2(new_n266), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n270), .A2(G274), .A3(new_n526), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n270), .A2(G250), .A3(new_n529), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n574), .A2(new_n575), .A3(KEYINPUT95), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(KEYINPUT95), .B1(new_n574), .B2(new_n575), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(G200), .B1(new_n573), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n578), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n581), .A2(new_n576), .B1(new_n572), .B2(new_n266), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(G190), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n566), .A2(new_n580), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n516), .A2(new_n564), .ZN(new_n585));
  INV_X1    g0385(.A(new_n565), .ZN(new_n586));
  AND3_X1   g0386(.A1(new_n561), .A2(new_n557), .A3(new_n555), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n585), .B(new_n586), .C1(new_n587), .C2(new_n554), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n357), .B1(new_n573), .B2(new_n579), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n582), .A2(new_n445), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n584), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n550), .A2(new_n553), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n270), .A2(G274), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n527), .A2(G270), .B1(new_n595), .B2(new_n530), .ZN(new_n596));
  OAI211_X1 g0396(.A(G264), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n597));
  OAI211_X1 g0397(.A(G257), .B(new_n334), .C1(new_n253), .C2(new_n254), .ZN(new_n598));
  INV_X1    g0398(.A(G303), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n597), .B(new_n598), .C1(new_n599), .C2(new_n251), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n266), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n596), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n353), .A2(G116), .A3(new_n514), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n306), .A2(new_n569), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n282), .A2(new_n213), .B1(G20), .B2(new_n569), .ZN(new_n605));
  AOI21_X1  g0405(.A(G20), .B1(G33), .B2(G283), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(G33), .B2(new_n502), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n605), .A2(new_n607), .A3(KEYINPUT20), .ZN(new_n608));
  AOI21_X1  g0408(.A(KEYINPUT20), .B1(new_n605), .B2(new_n607), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n603), .B(new_n604), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n602), .A2(KEYINPUT21), .A3(new_n610), .A4(G169), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT97), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n357), .B1(new_n596), .B2(new_n601), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n614), .A2(KEYINPUT97), .A3(KEYINPUT21), .A4(new_n610), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n614), .A2(new_n610), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT21), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n602), .A2(new_n445), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n617), .A2(new_n618), .B1(new_n619), .B2(new_n610), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n610), .B1(new_n602), .B2(G200), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n364), .B2(new_n602), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n616), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n306), .A2(KEYINPUT25), .A3(new_n337), .ZN(new_n624));
  AOI21_X1  g0424(.A(KEYINPUT25), .B1(new_n306), .B2(new_n337), .ZN(new_n625));
  OAI22_X1  g0425(.A1(new_n515), .A2(new_n337), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n410), .A2(KEYINPUT98), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n251), .A2(new_n207), .A3(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT22), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n251), .A2(KEYINPUT22), .A3(new_n207), .A4(new_n627), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT23), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(new_n207), .B2(G107), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n337), .A2(KEYINPUT23), .A3(G20), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n633), .A2(new_n634), .B1(new_n570), .B2(new_n207), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n630), .A2(new_n631), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT24), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT24), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n630), .A2(new_n638), .A3(new_n631), .A4(new_n635), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n626), .B1(new_n640), .B2(new_n283), .ZN(new_n641));
  OAI211_X1 g0441(.A(G257), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n642));
  OAI211_X1 g0442(.A(G250), .B(new_n334), .C1(new_n253), .C2(new_n254), .ZN(new_n643));
  INV_X1    g0443(.A(G294), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n642), .B(new_n643), .C1(new_n295), .C2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n266), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT99), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n645), .A2(KEYINPUT99), .A3(new_n266), .ZN(new_n649));
  INV_X1    g0449(.A(new_n523), .ZN(new_n650));
  NOR2_X1   g0450(.A1(KEYINPUT5), .A2(G41), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n526), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n652), .A2(G264), .A3(new_n270), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n531), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n648), .A2(new_n364), .A3(new_n649), .A4(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n646), .A2(new_n531), .A3(new_n653), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n316), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n641), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n654), .B1(new_n646), .B2(new_n647), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n357), .B1(new_n661), .B2(new_n649), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n657), .A2(new_n445), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n554), .B1(new_n637), .B2(new_n639), .ZN(new_n664));
  OAI22_X1  g0464(.A1(new_n662), .A2(new_n663), .B1(new_n664), .B2(new_n626), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n623), .A2(new_n666), .ZN(new_n667));
  NOR3_X1   g0467(.A1(new_n494), .A2(new_n593), .A3(new_n667), .ZN(G372));
  AND2_X1   g0468(.A1(new_n420), .A2(new_n431), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n360), .B1(new_n480), .B2(new_n483), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n473), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n427), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n326), .A2(new_n330), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n315), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n665), .A2(new_n616), .A3(new_n620), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n660), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n591), .B1(new_n593), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n584), .A2(new_n591), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT26), .ZN(new_n681));
  NOR3_X1   g0481(.A1(new_n553), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n551), .A2(new_n552), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n548), .B1(new_n512), .B2(new_n517), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n512), .A2(new_n548), .A3(new_n517), .ZN(new_n685));
  OAI211_X1 g0485(.A(new_n592), .B(new_n683), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n682), .B1(new_n686), .B2(new_n681), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n679), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n676), .B1(new_n494), .B2(new_n689), .ZN(G369));
  NAND3_X1  g0490(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n691), .A2(KEYINPUT27), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(KEYINPUT27), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(G213), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(G343), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n610), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n623), .A2(new_n697), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n616), .A2(new_n620), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n698), .B1(new_n699), .B2(new_n697), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(G330), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n696), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n666), .B1(new_n641), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n665), .B2(new_n703), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n699), .A2(new_n696), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n666), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n665), .B2(new_n696), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n707), .A2(new_n710), .ZN(G399));
  INV_X1    g0511(.A(new_n210), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(G41), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n560), .A2(G116), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n714), .A2(G1), .A3(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT100), .ZN(new_n717));
  OAI22_X1  g0517(.A1(new_n716), .A2(new_n717), .B1(new_n217), .B2(new_n714), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n718), .B1(new_n717), .B2(new_n716), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT101), .ZN(new_n720));
  XOR2_X1   g0520(.A(new_n720), .B(KEYINPUT28), .Z(new_n721));
  NAND2_X1  g0521(.A1(new_n686), .A2(KEYINPUT26), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n592), .A2(new_n683), .A3(new_n681), .A4(new_n518), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n703), .B1(new_n724), .B2(new_n679), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(KEYINPUT29), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT29), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n727), .B(new_n703), .C1(new_n679), .C2(new_n687), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(G330), .ZN(new_n731));
  OR3_X1    g0531(.A1(new_n593), .A2(new_n667), .A3(new_n696), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT30), .ZN(new_n733));
  INV_X1    g0533(.A(new_n602), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n646), .A2(new_n653), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n734), .A2(new_n735), .A3(new_n582), .A4(G179), .ZN(new_n736));
  INV_X1    g0536(.A(new_n545), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n733), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n734), .A2(new_n582), .A3(G179), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n739), .A2(new_n737), .A3(new_n657), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n735), .A2(new_n582), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n741), .A2(KEYINPUT30), .A3(new_n545), .A4(new_n619), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n738), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n696), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT31), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n743), .A2(KEYINPUT31), .A3(new_n696), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n731), .B1(new_n732), .B2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n730), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n721), .B1(new_n753), .B2(G1), .ZN(G364));
  INV_X1    g0554(.A(G13), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n206), .B1(new_n756), .B2(G45), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n713), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n712), .A2(new_n255), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT102), .ZN(new_n761));
  NAND2_X1  g0561(.A1(G355), .A2(new_n761), .ZN(new_n762));
  OR2_X1    g0562(.A1(G355), .A2(new_n761), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n760), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n764), .B1(G116), .B2(new_n210), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n245), .A2(new_n525), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n712), .A2(new_n251), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n768), .B1(new_n218), .B2(new_n525), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n765), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(G20), .B1(KEYINPUT103), .B2(G169), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(KEYINPUT103), .B2(G169), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n213), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n773), .A2(KEYINPUT104), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(KEYINPUT104), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G13), .A2(G33), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G20), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n759), .B1(new_n770), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n776), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n445), .A2(new_n316), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT105), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n207), .A2(G190), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n382), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT32), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n207), .A2(G179), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n791), .A2(new_n364), .A3(G200), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n337), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n791), .A2(G190), .A3(G200), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n255), .B(new_n793), .C1(G87), .C2(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT106), .ZN(new_n797));
  NAND2_X1  g0597(.A1(G20), .A2(G179), .ZN(new_n798));
  NOR3_X1   g0598(.A1(new_n798), .A2(new_n316), .A3(G190), .ZN(new_n799));
  NOR3_X1   g0599(.A1(new_n798), .A2(G190), .A3(G200), .ZN(new_n800));
  AOI22_X1  g0600(.A1(G68), .A2(new_n799), .B1(new_n800), .B2(G77), .ZN(new_n801));
  NOR3_X1   g0601(.A1(new_n798), .A2(new_n364), .A3(new_n316), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n798), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n804), .A2(G190), .A3(new_n316), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n801), .B1(new_n201), .B2(new_n803), .C1(new_n202), .C2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n207), .B1(new_n786), .B2(G190), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n806), .B1(new_n808), .B2(G97), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n790), .A2(new_n797), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n808), .A2(G294), .ZN(new_n811));
  INV_X1    g0611(.A(G283), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n792), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n799), .ZN(new_n814));
  INV_X1    g0614(.A(G317), .ZN(new_n815));
  AND2_X1   g0615(.A1(new_n815), .A2(KEYINPUT33), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n815), .A2(KEYINPUT33), .ZN(new_n817));
  NOR3_X1   g0617(.A1(new_n814), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n813), .B(new_n818), .C1(G326), .C2(new_n802), .ZN(new_n819));
  INV_X1    g0619(.A(new_n788), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(G329), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n255), .B1(new_n794), .B2(new_n599), .ZN(new_n822));
  INV_X1    g0622(.A(new_n800), .ZN(new_n823));
  INV_X1    g0623(.A(G311), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n805), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n822), .B(new_n825), .C1(G322), .C2(new_n826), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n811), .A2(new_n819), .A3(new_n821), .A4(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n783), .B1(new_n810), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n782), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n779), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n830), .B1(new_n700), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n759), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n701), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n700), .A2(G330), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n832), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT107), .ZN(G396));
  NAND2_X1  g0637(.A1(new_n356), .A2(new_n696), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n361), .A2(KEYINPUT77), .ZN(new_n839));
  INV_X1    g0639(.A(new_n365), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n838), .B1(new_n841), .B2(new_n362), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n359), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n359), .A2(new_n696), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n689), .B2(new_n696), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n844), .B1(new_n842), .B2(new_n359), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n848), .B(new_n703), .C1(new_n679), .C2(new_n687), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n759), .B1(new_n850), .B2(new_n751), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n751), .B2(new_n850), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n776), .A2(new_n777), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n759), .B1(new_n854), .B2(G77), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n808), .A2(G97), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n820), .A2(G311), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n792), .A2(new_n410), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n255), .B1(new_n803), .B2(new_n599), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n858), .B(new_n859), .C1(G116), .C2(new_n800), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n794), .A2(new_n337), .B1(new_n805), .B2(new_n644), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(G283), .B2(new_n799), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n856), .A2(new_n857), .A3(new_n860), .A4(new_n862), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n826), .A2(G143), .B1(G137), .B2(new_n802), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n864), .B1(new_n300), .B2(new_n814), .C1(new_n382), .C2(new_n823), .ZN(new_n865));
  XOR2_X1   g0665(.A(new_n865), .B(KEYINPUT34), .Z(new_n866));
  NOR2_X1   g0666(.A1(new_n792), .A2(new_n374), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n255), .B(new_n867), .C1(G50), .C2(new_n795), .ZN(new_n868));
  INV_X1    g0668(.A(G132), .ZN(new_n869));
  OAI221_X1 g0669(.A(new_n868), .B1(new_n869), .B2(new_n788), .C1(new_n202), .C2(new_n807), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n863), .B1(new_n866), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n855), .B1(new_n871), .B2(new_n776), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n848), .B2(new_n778), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n852), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(G384));
  NOR2_X1   g0675(.A1(new_n756), .A2(new_n206), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT40), .ZN(new_n877));
  NOR3_X1   g0677(.A1(new_n593), .A2(new_n667), .A3(new_n696), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n848), .B1(new_n878), .B2(new_n748), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n461), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n484), .B2(new_n488), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n482), .A2(new_n703), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n883), .B1(new_n486), .B2(new_n487), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n473), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT108), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT83), .B1(new_n480), .B2(new_n483), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n486), .A2(new_n487), .A3(new_n485), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n461), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n883), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n886), .B(KEYINPUT108), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n880), .B1(new_n887), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n421), .A2(new_n424), .ZN(new_n895));
  INV_X1    g0695(.A(new_n694), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n421), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT37), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n895), .A2(new_n897), .A3(new_n898), .A4(new_n416), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n390), .A2(new_n397), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n424), .B2(new_n896), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n416), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT37), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT38), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n694), .B1(new_n390), .B2(new_n397), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n905), .B1(new_n432), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n432), .A2(new_n906), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n904), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT38), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n907), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n877), .B1(new_n894), .B2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT110), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n886), .B1(new_n890), .B2(new_n891), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT108), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n879), .B1(new_n917), .B2(new_n892), .ZN(new_n918));
  INV_X1    g0718(.A(new_n905), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n908), .A2(new_n919), .ZN(new_n920));
  AND2_X1   g0720(.A1(new_n899), .A2(new_n903), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(new_n432), .B2(new_n906), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n920), .B1(KEYINPUT38), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n918), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n924), .A2(KEYINPUT110), .A3(new_n877), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n914), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n895), .A2(new_n897), .A3(new_n416), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(KEYINPUT37), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n928), .A2(new_n899), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n418), .A2(new_n419), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n897), .B1(new_n427), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n910), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n877), .B1(new_n920), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n918), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n926), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n369), .A2(new_n371), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n432), .A2(KEYINPUT88), .ZN(new_n937));
  AND4_X1   g0737(.A1(new_n936), .A2(new_n937), .A3(new_n434), .A4(new_n493), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n878), .B2(new_n748), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n935), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(G330), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n935), .B2(new_n939), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n473), .A2(new_n696), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT109), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT39), .ZN(new_n947));
  INV_X1    g0747(.A(new_n426), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n421), .A2(new_n422), .A3(new_n424), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n948), .A2(new_n429), .A3(new_n949), .A4(new_n430), .ZN(new_n950));
  INV_X1    g0750(.A(new_n897), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n950), .A2(new_n951), .B1(new_n928), .B2(new_n899), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n947), .B1(new_n952), .B2(KEYINPUT38), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n946), .B1(new_n953), .B2(new_n907), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n920), .A2(new_n932), .A3(KEYINPUT109), .A4(new_n947), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n923), .A2(KEYINPUT39), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n945), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n917), .A2(new_n892), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n849), .A2(new_n845), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n961), .A2(new_n911), .B1(new_n427), .B2(new_n896), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n958), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n673), .A2(new_n675), .ZN(new_n964));
  INV_X1    g0764(.A(new_n315), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(new_n938), .B2(new_n729), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n963), .B(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n876), .B1(new_n943), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n968), .B2(new_n943), .ZN(new_n970));
  AOI211_X1 g0770(.A(new_n569), .B(new_n215), .C1(new_n506), .C2(KEYINPUT35), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(KEYINPUT35), .B2(new_n506), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT36), .ZN(new_n973));
  OAI21_X1  g0773(.A(G77), .B1(new_n202), .B2(new_n374), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n974), .A2(new_n217), .B1(G50), .B2(new_n374), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n975), .A2(G1), .A3(new_n755), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n970), .A2(new_n973), .A3(new_n976), .ZN(G367));
  OAI22_X1  g0777(.A1(new_n768), .A2(new_n235), .B1(new_n210), .B2(new_n349), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n759), .B1(new_n781), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n802), .A2(G143), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n300), .B2(new_n805), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n807), .A2(new_n374), .ZN(new_n982));
  INV_X1    g0782(.A(new_n792), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n981), .B(new_n982), .C1(G77), .C2(new_n983), .ZN(new_n984));
  AOI22_X1  g0784(.A1(G50), .A2(new_n800), .B1(new_n799), .B2(G159), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n985), .B(new_n251), .C1(new_n202), .C2(new_n794), .ZN(new_n986));
  XNOR2_X1  g0786(.A(KEYINPUT114), .B(G137), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n986), .B1(new_n820), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n255), .B1(new_n792), .B2(new_n502), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n794), .A2(new_n569), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT46), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n990), .B(new_n992), .C1(G317), .C2(new_n820), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n823), .A2(new_n812), .B1(new_n805), .B2(new_n599), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n803), .A2(new_n824), .B1(new_n814), .B2(new_n644), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n994), .B(new_n995), .C1(new_n808), .C2(G107), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n984), .A2(new_n989), .B1(new_n993), .B2(new_n996), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n997), .A2(KEYINPUT47), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n783), .B1(new_n997), .B2(KEYINPUT47), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n979), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n566), .A2(new_n703), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n680), .A2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n1001), .A2(new_n590), .A3(new_n588), .A4(new_n589), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1000), .B1(new_n831), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n696), .B1(new_n685), .B2(new_n684), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n550), .A2(new_n1006), .A3(new_n553), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n683), .B(new_n696), .C1(new_n684), .C2(new_n685), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n710), .A2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT112), .Z(new_n1012));
  OR2_X1    g0812(.A1(new_n1012), .A2(KEYINPUT44), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(KEYINPUT44), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n710), .A2(new_n1010), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT45), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1013), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n707), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n702), .A2(KEYINPUT113), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n709), .B1(new_n705), .B2(new_n708), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1019), .B(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n753), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1013), .A2(new_n1014), .A3(new_n706), .A4(new_n1016), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1018), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n753), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n713), .B(KEYINPUT41), .Z(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n758), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n553), .B1(new_n1010), .B2(new_n665), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n703), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1009), .A2(new_n666), .A3(new_n708), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT42), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1031), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1004), .A2(KEYINPUT43), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1004), .A2(KEYINPUT43), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1039), .A2(KEYINPUT111), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(KEYINPUT111), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n706), .A2(new_n1010), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1043), .B(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1005), .B1(new_n1029), .B2(new_n1046), .ZN(G387));
  INV_X1    g0847(.A(new_n1021), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n752), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1049), .A2(new_n1022), .A3(new_n713), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1021), .A2(new_n758), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n715), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n760), .A2(new_n1052), .B1(new_n337), .B2(new_n712), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n232), .A2(new_n525), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n347), .A2(new_n201), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT50), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n715), .B(new_n525), .C1(new_n374), .C2(new_n350), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n767), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1053), .B1(new_n1054), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n833), .B1(new_n1059), .B2(new_n780), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n396), .A2(new_n814), .B1(new_n374), .B2(new_n823), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT116), .Z(new_n1062));
  NAND2_X1  g0862(.A1(new_n808), .A2(new_n564), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n794), .A2(new_n350), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n251), .B1(new_n792), .B2(new_n502), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1064), .B(new_n1065), .C1(G50), .C2(new_n826), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n820), .A2(G150), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n802), .A2(G159), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT115), .Z(new_n1069));
  NAND4_X1  g0869(.A1(new_n1063), .A2(new_n1066), .A3(new_n1067), .A4(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1062), .A2(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT117), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n820), .A2(G326), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n255), .B1(new_n792), .B2(new_n569), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n823), .A2(new_n599), .B1(new_n805), .B2(new_n815), .ZN(new_n1075));
  OR2_X1    g0875(.A1(new_n1075), .A2(KEYINPUT118), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(KEYINPUT118), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(G322), .A2(new_n802), .B1(new_n799), .B2(G311), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT119), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n1081), .A2(KEYINPUT48), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1081), .A2(KEYINPUT48), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n807), .A2(new_n812), .B1(new_n644), .B2(new_n794), .ZN(new_n1084));
  NOR3_X1   g0884(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n1073), .B(new_n1074), .C1(new_n1085), .C2(KEYINPUT49), .ZN(new_n1086));
  OR2_X1    g0886(.A1(new_n1085), .A2(KEYINPUT49), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1072), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1060), .B1(new_n705), .B2(new_n831), .C1(new_n1088), .C2(new_n783), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n1051), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1050), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT120), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1050), .A2(KEYINPUT120), .A3(new_n1090), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(new_n1094), .ZN(G393));
  AND2_X1   g0895(.A1(new_n1018), .A2(new_n1024), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n758), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n780), .B1(new_n502), .B2(new_n210), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n240), .A2(new_n767), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n759), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n255), .B(new_n858), .C1(new_n820), .C2(G143), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n347), .A2(new_n800), .B1(new_n799), .B2(G50), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1101), .B(new_n1102), .C1(new_n374), .C2(new_n794), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n826), .A2(G159), .B1(G150), .B2(new_n802), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n808), .A2(G77), .B1(KEYINPUT51), .B2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(KEYINPUT51), .B2(new_n1104), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n251), .B(new_n793), .C1(new_n820), .C2(G322), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n644), .A2(new_n823), .B1(new_n814), .B2(new_n599), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(G283), .B2(new_n795), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1107), .B(new_n1109), .C1(new_n569), .C2(new_n807), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n826), .A2(G311), .B1(G317), .B2(new_n802), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT52), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n1103), .A2(new_n1106), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1100), .B1(new_n1113), .B2(new_n776), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n1009), .B2(new_n831), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1096), .A2(new_n1023), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1025), .A2(new_n713), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1097), .B(new_n1115), .C1(new_n1116), .C2(new_n1117), .ZN(G390));
  NAND2_X1  g0918(.A1(new_n961), .A2(new_n945), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1119), .A2(new_n956), .A3(new_n957), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n944), .B1(new_n920), .B2(new_n932), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n959), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n703), .B(new_n843), .C1(new_n724), .C2(new_n679), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n1123), .A2(new_n845), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1121), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1120), .A2(new_n1125), .ZN(new_n1126));
  OAI211_X1 g0926(.A(G330), .B(new_n848), .C1(new_n878), .C2(new_n748), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n959), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1126), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1120), .A2(new_n1129), .A3(new_n1125), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n433), .A2(new_n434), .A3(new_n493), .A4(new_n750), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1127), .A2(new_n917), .A3(new_n892), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1129), .A2(new_n1124), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n1129), .A2(new_n1135), .B1(new_n845), .B2(new_n849), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n967), .B(new_n1134), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n714), .B1(new_n1133), .B2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n676), .B(new_n1134), .C1(new_n730), .C2(new_n494), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1129), .A2(new_n1135), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n960), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n1136), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1131), .A2(new_n1132), .A3(new_n1142), .A4(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1140), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1131), .A2(new_n758), .A3(new_n1132), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT124), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n956), .A2(new_n777), .A3(new_n957), .ZN(new_n1150));
  XOR2_X1   g0950(.A(KEYINPUT54), .B(G143), .Z(new_n1151));
  AOI22_X1  g0951(.A1(new_n988), .A2(new_n799), .B1(new_n1151), .B2(new_n800), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n807), .B2(new_n382), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT121), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n255), .B1(new_n802), .B2(G128), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(G50), .A2(new_n983), .B1(new_n826), .B2(G132), .ZN(new_n1156));
  OR3_X1    g0956(.A1(new_n794), .A2(KEYINPUT53), .A3(new_n300), .ZN(new_n1157));
  OAI21_X1  g0957(.A(KEYINPUT53), .B1(new_n794), .B2(new_n300), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n820), .B2(G125), .ZN(new_n1160));
  AND4_X1   g0960(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .A4(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n867), .B1(G283), .B2(new_n802), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1162), .B1(new_n569), .B2(new_n805), .C1(new_n788), .C2(new_n644), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n502), .A2(new_n823), .B1(new_n814), .B2(new_n337), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(KEYINPUT122), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n807), .B2(new_n350), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1164), .A2(KEYINPUT122), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n255), .B1(new_n794), .B2(new_n410), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT123), .ZN(new_n1169));
  NOR4_X1   g0969(.A1(new_n1163), .A2(new_n1166), .A3(new_n1167), .A4(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n776), .B1(new_n1161), .B2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n833), .B1(new_n853), .B2(new_n396), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1150), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1148), .A2(new_n1149), .A3(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1149), .B1(new_n1148), .B2(new_n1173), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1147), .B1(new_n1175), .B2(new_n1176), .ZN(G378));
  OAI21_X1  g0977(.A(new_n759), .B1(new_n854), .B2(G50), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n201), .B1(G33), .B2(G41), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n255), .B2(new_n521), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n803), .A2(new_n569), .B1(new_n814), .B2(new_n502), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1181), .B(new_n982), .C1(new_n564), .C2(new_n800), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n792), .A2(new_n202), .B1(new_n805), .B2(new_n337), .ZN(new_n1183));
  NOR4_X1   g0983(.A1(new_n1183), .A2(new_n1064), .A3(G41), .A4(new_n251), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1182), .B(new_n1184), .C1(new_n812), .C2(new_n788), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT58), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1180), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n826), .A2(G128), .B1(G125), .B2(new_n802), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(G137), .B2(new_n800), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n795), .A2(new_n1151), .B1(G132), .B2(new_n799), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1190), .B(new_n1191), .C1(new_n300), .C2(new_n807), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1192), .A2(KEYINPUT59), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(KEYINPUT59), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n295), .B(new_n521), .C1(new_n792), .C2(new_n382), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(new_n820), .B2(G124), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1187), .B1(new_n1186), .B2(new_n1185), .C1(new_n1193), .C2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1178), .B1(new_n1198), .B2(new_n776), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n313), .A2(new_n694), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n331), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n331), .A2(new_n1201), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  OR3_X1    g1006(.A1(new_n1203), .A2(new_n1204), .A3(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1206), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1199), .B1(new_n1209), .B2(new_n778), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT125), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n963), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n731), .B1(new_n933), .B2(new_n918), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1209), .B1(new_n926), .B2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(KEYINPUT110), .B1(new_n924), .B2(new_n877), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n913), .B(KEYINPUT40), .C1(new_n918), .C2(new_n923), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1209), .B(new_n1213), .C1(new_n1215), .C2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1212), .B1(new_n1214), .B2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1213), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1209), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1222), .A2(new_n963), .A3(new_n1217), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1219), .A2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1211), .B1(new_n1224), .B2(new_n758), .ZN(new_n1225));
  AND3_X1   g1025(.A1(new_n1222), .A2(new_n963), .A3(new_n1217), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n963), .B1(new_n1222), .B2(new_n1217), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n1120), .A2(new_n1129), .A3(new_n1125), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1129), .B1(new_n1120), .B2(new_n1125), .ZN(new_n1230));
  NOR3_X1   g1030(.A1(new_n1229), .A2(new_n1230), .A3(new_n1139), .ZN(new_n1231));
  OAI21_X1  g1031(.A(KEYINPUT57), .B1(new_n1231), .B2(new_n1141), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n713), .B1(new_n1228), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1146), .A2(new_n1142), .ZN(new_n1234));
  AOI21_X1  g1034(.A(KEYINPUT57), .B1(new_n1224), .B2(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1225), .B1(new_n1233), .B2(new_n1235), .ZN(G375));
  NAND2_X1  g1036(.A1(new_n1145), .A2(new_n758), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n759), .B1(new_n854), .B2(G68), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n808), .A2(G50), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n803), .A2(new_n869), .B1(new_n823), .B2(new_n300), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n255), .B(new_n1240), .C1(G58), .C2(new_n983), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n820), .A2(G128), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n794), .A2(new_n382), .B1(new_n805), .B2(new_n987), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n799), .B2(new_n1151), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1239), .A2(new_n1241), .A3(new_n1242), .A4(new_n1244), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n803), .A2(new_n644), .B1(new_n823), .B2(new_n337), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(G116), .B2(new_n799), .ZN(new_n1247));
  XOR2_X1   g1047(.A(new_n1247), .B(KEYINPUT126), .Z(new_n1248));
  NAND2_X1  g1048(.A1(new_n820), .A2(G303), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n251), .B1(new_n983), .B2(G77), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(G97), .A2(new_n795), .B1(new_n826), .B2(G283), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1063), .A2(new_n1249), .A3(new_n1250), .A4(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1245), .B1(new_n1248), .B2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1238), .B1(new_n1253), .B2(new_n776), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1254), .B1(new_n959), .B2(new_n778), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1237), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1141), .A2(new_n1144), .A3(new_n1136), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1139), .A2(new_n1258), .A3(new_n1028), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1257), .A2(new_n1259), .ZN(G381));
  INV_X1    g1060(.A(G390), .ZN(new_n1261));
  INV_X1    g1061(.A(G381), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(G393), .A2(G396), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1261), .A2(new_n874), .A3(new_n1262), .A4(new_n1263), .ZN(new_n1264));
  OR4_X1    g1064(.A1(G387), .A2(new_n1264), .A3(G378), .A4(G375), .ZN(G407));
  INV_X1    g1065(.A(new_n1176), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n1266), .A2(new_n1174), .B1(new_n1140), .B2(new_n1146), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n695), .A2(G213), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1267), .A2(new_n1269), .ZN(new_n1270));
  OAI211_X1 g1070(.A(G407), .B(G213), .C1(G375), .C2(new_n1270), .ZN(G409));
  OAI211_X1 g1071(.A(G378), .B(new_n1225), .C1(new_n1233), .C2(new_n1235), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1234), .B(new_n1028), .C1(new_n1226), .C2(new_n1227), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1211), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n758), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1273), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1267), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1272), .A2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n1268), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1269), .A2(G2897), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1141), .A2(new_n1144), .A3(KEYINPUT60), .A4(new_n1136), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n713), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT60), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1258), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n1139), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(KEYINPUT127), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT127), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1285), .A2(new_n1288), .A3(new_n1139), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1283), .B1(new_n1287), .B2(new_n1289), .ZN(new_n1290));
  NOR3_X1   g1090(.A1(new_n1290), .A2(new_n874), .A3(new_n1256), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1283), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1285), .A2(new_n1288), .A3(new_n1139), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1288), .B1(new_n1285), .B2(new_n1139), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1292), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(G384), .B1(new_n1295), .B2(new_n1257), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1281), .B1(new_n1291), .B2(new_n1296), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n874), .B1(new_n1290), .B2(new_n1256), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1295), .A2(G384), .A3(new_n1257), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1298), .A2(new_n1299), .A3(new_n1280), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1297), .A2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(KEYINPUT61), .B1(new_n1279), .B2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT63), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1291), .A2(new_n1296), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1303), .B1(new_n1279), .B2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1261), .A2(G387), .ZN(new_n1307));
  OAI211_X1 g1107(.A(G390), .B(new_n1005), .C1(new_n1029), .C2(new_n1046), .ZN(new_n1308));
  XOR2_X1   g1108(.A(G393), .B(G396), .Z(new_n1309));
  AND3_X1   g1109(.A1(new_n1307), .A2(new_n1308), .A3(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1309), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1269), .B1(new_n1272), .B2(new_n1277), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1313), .A2(KEYINPUT63), .A3(new_n1304), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1302), .A2(new_n1306), .A3(new_n1312), .A4(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT62), .ZN(new_n1316));
  AND3_X1   g1116(.A1(new_n1313), .A2(new_n1316), .A3(new_n1304), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT61), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1297), .A2(new_n1300), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1318), .B1(new_n1313), .B2(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1316), .B1(new_n1313), .B2(new_n1304), .ZN(new_n1321));
  NOR3_X1   g1121(.A1(new_n1317), .A2(new_n1320), .A3(new_n1321), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1315), .B1(new_n1322), .B2(new_n1312), .ZN(G405));
  AND2_X1   g1123(.A1(G375), .A2(new_n1267), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1272), .ZN(new_n1325));
  OR3_X1    g1125(.A1(new_n1324), .A2(new_n1325), .A3(new_n1304), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1304), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1312), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1326), .A2(new_n1312), .A3(new_n1327), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(G402));
endmodule


