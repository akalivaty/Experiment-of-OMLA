//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 1 0 0 0 0 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1273,
    new_n1274, new_n1275, new_n1276, new_n1277, new_n1278, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  INV_X1    g0007(.A(G77), .ZN(new_n208));
  NAND3_X1  g0008(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT65), .ZN(G353));
  OAI21_X1  g0010(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NOR2_X1   g0011(.A1(new_n206), .A2(new_n207), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G1), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n214), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(G13), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT0), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  XOR2_X1   g0023(.A(KEYINPUT66), .B(G238), .Z(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT67), .B(G77), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n203), .C1(new_n225), .C2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(KEYINPUT68), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n228), .A2(KEYINPUT68), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n219), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n216), .B(new_n222), .C1(new_n234), .C2(KEYINPUT1), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n235), .B1(KEYINPUT1), .B2(new_n234), .ZN(G361));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT69), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  INV_X1    g0041(.A(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT2), .B(G226), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n240), .B(new_n245), .ZN(G358));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n207), .A2(G68), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n203), .A2(G50), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G58), .B(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n249), .B(new_n254), .ZN(G351));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1698), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n260), .A2(G222), .A3(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G223), .ZN(new_n263));
  AND2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  OAI21_X1  g0065(.A(G1698), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OAI221_X1 g0066(.A(new_n262), .B1(new_n263), .B2(new_n266), .C1(new_n227), .C2(new_n260), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G41), .ZN(new_n270));
  INV_X1    g0070(.A(G45), .ZN(new_n271));
  AOI21_X1  g0071(.A(G1), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(G1), .A3(G13), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n272), .A2(new_n274), .A3(G274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n268), .A2(new_n272), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n276), .B1(G226), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n269), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G200), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n213), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n214), .B1(new_n206), .B2(new_n207), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT8), .B(G58), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n214), .A2(G33), .ZN(new_n285));
  INV_X1    g0085(.A(G150), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  OAI22_X1  g0088(.A1(new_n284), .A2(new_n285), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n282), .B1(new_n283), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n217), .A2(G13), .A3(G20), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(new_n213), .A3(new_n281), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n207), .B1(new_n217), .B2(G20), .ZN(new_n294));
  INV_X1    g0094(.A(new_n291), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n293), .A2(new_n294), .B1(new_n207), .B2(new_n295), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n290), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G190), .ZN(new_n298));
  OAI221_X1 g0098(.A(new_n280), .B1(KEYINPUT9), .B2(new_n297), .C1(new_n298), .C2(new_n279), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(KEYINPUT9), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT71), .ZN(new_n301));
  OR3_X1    g0101(.A1(new_n299), .A2(new_n301), .A3(KEYINPUT10), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT10), .B1(new_n299), .B2(new_n301), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G169), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n297), .B1(new_n279), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(G179), .B2(new_n279), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  OAI22_X1  g0108(.A1(new_n285), .A2(new_n208), .B1(new_n214), .B2(G68), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT72), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(new_n288), .B2(new_n207), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n287), .A2(KEYINPUT72), .A3(G50), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n309), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT11), .ZN(new_n314));
  INV_X1    g0114(.A(new_n282), .ZN(new_n315));
  OR3_X1    g0115(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n314), .B1(new_n313), .B2(new_n315), .ZN(new_n317));
  OAI21_X1  g0117(.A(KEYINPUT12), .B1(new_n291), .B2(G68), .ZN(new_n318));
  OR3_X1    g0118(.A1(new_n291), .A2(KEYINPUT12), .A3(G68), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n203), .B1(new_n217), .B2(G20), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n318), .A2(new_n319), .B1(new_n293), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n316), .A2(new_n317), .A3(new_n321), .ZN(new_n322));
  OAI211_X1 g0122(.A(G232), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n323));
  OAI211_X1 g0123(.A(G226), .B(new_n261), .C1(new_n264), .C2(new_n265), .ZN(new_n324));
  NAND2_X1  g0124(.A1(G33), .A2(G97), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n268), .ZN(new_n327));
  INV_X1    g0127(.A(G274), .ZN(new_n328));
  INV_X1    g0128(.A(new_n213), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n328), .B1(new_n329), .B2(new_n273), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n277), .A2(G238), .B1(new_n330), .B2(new_n272), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT13), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT13), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n327), .A2(new_n331), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n333), .A2(G179), .A3(new_n335), .ZN(new_n336));
  AND3_X1   g0136(.A1(new_n327), .A2(new_n331), .A3(new_n334), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n334), .B1(new_n327), .B2(new_n331), .ZN(new_n338));
  OAI21_X1  g0138(.A(G169), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n336), .B1(new_n339), .B2(KEYINPUT14), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT14), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n333), .A2(new_n335), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n341), .B1(new_n342), .B2(G169), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n322), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n322), .ZN(new_n345));
  OAI21_X1  g0145(.A(G200), .B1(new_n337), .B2(new_n338), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n333), .A2(G190), .A3(new_n335), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n284), .B1(new_n217), .B2(G20), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n350), .A2(new_n293), .B1(new_n295), .B2(new_n284), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n258), .A2(new_n214), .A3(new_n259), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT7), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT73), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n258), .A2(KEYINPUT7), .A3(new_n214), .A4(new_n259), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n357), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(KEYINPUT73), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n358), .A2(G68), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(G58), .A2(G68), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n204), .A2(new_n205), .A3(new_n362), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n363), .A2(G20), .B1(G159), .B2(new_n287), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT16), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n203), .B1(new_n355), .B2(new_n357), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n363), .A2(G20), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n287), .A2(G159), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n315), .B1(new_n372), .B2(KEYINPUT16), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n352), .B1(new_n367), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(G226), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G1698), .ZN(new_n376));
  OAI221_X1 g0176(.A(new_n376), .B1(G223), .B2(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n377));
  NAND2_X1  g0177(.A1(G33), .A2(G87), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n274), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n217), .B1(G41), .B2(G45), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n274), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n275), .B1(new_n242), .B2(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G179), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n305), .B2(new_n383), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(KEYINPUT18), .B1(new_n374), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n383), .A2(new_n298), .ZN(new_n388));
  INV_X1    g0188(.A(G200), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n379), .B2(new_n382), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n374), .A2(KEYINPUT17), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(KEYINPUT16), .B1(new_n361), .B2(new_n364), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n264), .A2(new_n265), .ZN(new_n394));
  AOI21_X1  g0194(.A(KEYINPUT7), .B1(new_n394), .B2(new_n214), .ZN(new_n395));
  OAI21_X1  g0195(.A(G68), .B1(new_n395), .B2(new_n359), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n396), .A2(KEYINPUT16), .A3(new_n364), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n282), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n391), .B(new_n351), .C1(new_n393), .C2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT17), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n351), .B1(new_n393), .B2(new_n398), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT18), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(new_n403), .A3(new_n385), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n387), .A2(new_n392), .A3(new_n401), .A4(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(G77), .B1(new_n214), .B2(G1), .ZN(new_n406));
  OAI22_X1  g0206(.A1(new_n292), .A2(new_n406), .B1(new_n226), .B2(new_n291), .ZN(new_n407));
  INV_X1    g0207(.A(new_n285), .ZN(new_n408));
  INV_X1    g0208(.A(G87), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(KEYINPUT15), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT15), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(G87), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n408), .A2(new_n413), .B1(new_n226), .B2(G20), .ZN(new_n414));
  INV_X1    g0214(.A(new_n284), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT70), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n287), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n288), .A2(KEYINPUT70), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n415), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n414), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n407), .B1(new_n420), .B2(new_n282), .ZN(new_n421));
  OAI211_X1 g0221(.A(G232), .B(new_n261), .C1(new_n264), .C2(new_n265), .ZN(new_n422));
  INV_X1    g0222(.A(G107), .ZN(new_n423));
  OAI221_X1 g0223(.A(new_n422), .B1(new_n260), .B2(new_n423), .C1(new_n224), .C2(new_n266), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n268), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n275), .B1(new_n225), .B2(new_n381), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n421), .B1(new_n428), .B2(new_n305), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n426), .B1(new_n424), .B2(new_n268), .ZN(new_n430));
  INV_X1    g0230(.A(G179), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n425), .A2(new_n427), .A3(G190), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n434), .B(new_n421), .C1(new_n389), .C2(new_n430), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NOR4_X1   g0236(.A1(new_n308), .A2(new_n349), .A3(new_n405), .A4(new_n436), .ZN(new_n437));
  AND3_X1   g0237(.A1(new_n358), .A2(G107), .A3(new_n360), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n287), .A2(G77), .ZN(new_n439));
  XOR2_X1   g0239(.A(new_n439), .B(KEYINPUT74), .Z(new_n440));
  XNOR2_X1  g0240(.A(KEYINPUT75), .B(G107), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(G97), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n443), .A2(new_n423), .A3(KEYINPUT6), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(KEYINPUT6), .B2(new_n443), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n441), .B(new_n444), .C1(KEYINPUT6), .C2(new_n443), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n440), .B1(new_n448), .B2(new_n214), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n282), .B1(new_n438), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n291), .A2(new_n443), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n217), .A2(G33), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n291), .A2(new_n452), .A3(new_n213), .A4(new_n281), .ZN(new_n453));
  OR2_X1    g0253(.A1(new_n453), .A2(KEYINPUT76), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(KEYINPUT76), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n451), .B1(new_n456), .B2(new_n443), .ZN(new_n457));
  OR2_X1    g0257(.A1(KEYINPUT5), .A2(G41), .ZN(new_n458));
  NAND2_X1  g0258(.A1(KEYINPUT5), .A2(G41), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n217), .A2(G45), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n463), .A2(G257), .A3(new_n274), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n461), .B1(new_n458), .B2(new_n459), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n330), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(G250), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n468), .B1(new_n258), .B2(new_n259), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT4), .ZN(new_n470));
  OAI21_X1  g0270(.A(G1698), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n470), .B1(new_n394), .B2(new_n225), .ZN(new_n472));
  NAND2_X1  g0272(.A1(G33), .A2(G283), .ZN(new_n473));
  AND2_X1   g0273(.A1(KEYINPUT4), .A2(G244), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n261), .B(new_n474), .C1(new_n264), .C2(new_n265), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n471), .A2(new_n472), .A3(new_n473), .A4(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n467), .B1(new_n476), .B2(new_n268), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n477), .A2(G200), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n464), .A2(new_n466), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n225), .B1(new_n258), .B2(new_n259), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n475), .B(new_n473), .C1(new_n480), .C2(KEYINPUT4), .ZN(new_n481));
  OAI21_X1  g0281(.A(G250), .B1(new_n264), .B2(new_n265), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n261), .B1(new_n482), .B2(KEYINPUT4), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n268), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n479), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(G190), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n450), .B(new_n457), .C1(new_n478), .C2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n450), .A2(new_n457), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n479), .A2(new_n484), .A3(G179), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n489), .B1(new_n477), .B2(new_n305), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n468), .B1(new_n271), .B2(G1), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n217), .A2(new_n328), .A3(G45), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n274), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT77), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n274), .A2(new_n493), .A3(new_n494), .A4(KEYINPUT77), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(G238), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n261), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n225), .A2(G1698), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n501), .B(new_n502), .C1(new_n264), .C2(new_n265), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G33), .A2(G116), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n268), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n389), .B1(new_n499), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n497), .A2(new_n498), .B1(new_n505), .B2(new_n268), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G190), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n454), .A2(new_n455), .A3(G87), .ZN(new_n511));
  OR2_X1    g0311(.A1(KEYINPUT79), .A2(G87), .ZN(new_n512));
  NAND2_X1  g0312(.A1(KEYINPUT79), .A2(G87), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n512), .A2(new_n443), .A3(new_n423), .A4(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT19), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n214), .B1(new_n325), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n260), .A2(new_n214), .A3(G68), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n515), .B1(new_n285), .B2(new_n443), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n413), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n520), .A2(new_n282), .B1(new_n295), .B2(new_n521), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n508), .A2(new_n510), .A3(new_n511), .A4(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n499), .A2(new_n506), .A3(new_n431), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT78), .ZN(new_n525));
  AOI21_X1  g0325(.A(G169), .B1(new_n499), .B2(new_n506), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n520), .A2(new_n282), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n454), .A2(new_n455), .A3(new_n413), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n521), .A2(new_n295), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT78), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n509), .A2(new_n532), .A3(new_n431), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n525), .A2(new_n527), .A3(new_n531), .A4(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n492), .A2(KEYINPUT80), .A3(new_n523), .A4(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT80), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n487), .A2(new_n491), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n534), .A2(new_n523), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n465), .A2(new_n268), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(G264), .ZN(new_n541));
  OAI211_X1 g0341(.A(G257), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n542));
  INV_X1    g0342(.A(G294), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n542), .B1(new_n257), .B2(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(G250), .B(new_n261), .C1(new_n264), .C2(new_n265), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT83), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n469), .A2(KEYINPUT83), .A3(new_n261), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n544), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n466), .B(new_n541), .C1(new_n549), .C2(new_n274), .ZN(new_n550));
  OR2_X1    g0350(.A1(new_n550), .A2(G179), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n305), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT24), .ZN(new_n553));
  AND2_X1   g0353(.A1(KEYINPUT81), .A2(G87), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n214), .B(new_n554), .C1(new_n264), .C2(new_n265), .ZN(new_n555));
  XNOR2_X1  g0355(.A(new_n555), .B(KEYINPUT22), .ZN(new_n556));
  OAI21_X1  g0356(.A(KEYINPUT23), .B1(new_n214), .B2(G107), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT23), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n558), .A2(new_n423), .A3(G20), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n214), .A2(G33), .A3(G116), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n557), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT82), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n557), .A2(new_n559), .A3(new_n560), .A4(KEYINPUT82), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n553), .B1(new_n556), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n556), .A2(new_n553), .A3(new_n565), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n315), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n456), .A2(G107), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n295), .A2(new_n423), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT25), .ZN(new_n572));
  XNOR2_X1  g0372(.A(new_n571), .B(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n551), .B(new_n552), .C1(new_n569), .C2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(G116), .ZN(new_n576));
  OR2_X1    g0376(.A1(new_n453), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n295), .A2(new_n576), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n281), .A2(new_n213), .B1(G20), .B2(new_n576), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n473), .B(new_n214), .C1(G33), .C2(new_n443), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n579), .A2(KEYINPUT20), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(KEYINPUT20), .B1(new_n579), .B2(new_n580), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n577), .B(new_n578), .C1(new_n581), .C2(new_n582), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n540), .A2(G270), .B1(new_n330), .B2(new_n465), .ZN(new_n584));
  OAI211_X1 g0384(.A(G264), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n585));
  OAI211_X1 g0385(.A(G257), .B(new_n261), .C1(new_n264), .C2(new_n265), .ZN(new_n586));
  INV_X1    g0386(.A(G303), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n585), .B(new_n586), .C1(new_n587), .C2(new_n260), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n268), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n583), .B1(new_n590), .B2(G200), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(new_n298), .B2(new_n590), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n590), .A2(G169), .A3(new_n583), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT21), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n590), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n596), .A2(G179), .A3(new_n583), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n590), .A2(KEYINPUT21), .A3(new_n583), .A4(G169), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n595), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n556), .A2(new_n553), .A3(new_n565), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n282), .B1(new_n600), .B2(new_n566), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n570), .A2(new_n573), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n550), .A2(G200), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n548), .A2(new_n547), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n268), .B1(new_n604), .B2(new_n544), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n605), .A2(G190), .A3(new_n466), .A4(new_n541), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n601), .A2(new_n602), .A3(new_n603), .A4(new_n606), .ZN(new_n607));
  AND4_X1   g0407(.A1(new_n575), .A2(new_n592), .A3(new_n599), .A4(new_n607), .ZN(new_n608));
  AND4_X1   g0408(.A1(new_n437), .A2(new_n535), .A3(new_n539), .A4(new_n608), .ZN(G372));
  INV_X1    g0409(.A(new_n307), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n387), .A2(new_n404), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n339), .A2(KEYINPUT14), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n342), .A2(new_n341), .A3(G169), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n612), .A2(new_n613), .A3(new_n336), .ZN(new_n614));
  INV_X1    g0414(.A(new_n433), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n614), .A2(new_n322), .B1(new_n615), .B2(new_n348), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n392), .A2(new_n401), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n611), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n610), .B1(new_n304), .B2(new_n618), .ZN(new_n619));
  NOR3_X1   g0419(.A1(new_n308), .A2(new_n405), .A3(new_n436), .ZN(new_n620));
  INV_X1    g0420(.A(new_n349), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n528), .A2(new_n511), .A3(new_n530), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n499), .A2(new_n506), .A3(G190), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n623), .A2(new_n624), .A3(new_n507), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n499), .A2(new_n506), .A3(new_n431), .ZN(new_n626));
  OAI21_X1  g0426(.A(KEYINPUT84), .B1(new_n626), .B2(new_n526), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT84), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n524), .B(new_n628), .C1(G169), .C2(new_n509), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n625), .B1(new_n630), .B2(new_n531), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n490), .A2(KEYINPUT85), .B1(new_n450), .B2(new_n457), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT26), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT85), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n489), .B(new_n634), .C1(new_n477), .C2(new_n305), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n631), .A2(new_n632), .A3(new_n633), .A4(new_n635), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n627), .A2(new_n629), .B1(new_n522), .B2(new_n529), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n488), .A2(new_n534), .A3(new_n490), .A4(new_n523), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n637), .B1(new_n638), .B2(KEYINPUT26), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n631), .A2(new_n491), .A3(new_n487), .A4(new_n607), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n595), .A2(new_n597), .A3(new_n598), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n602), .A2(new_n601), .B1(new_n305), .B2(new_n550), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n641), .B1(new_n642), .B2(new_n551), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n636), .B(new_n639), .C1(new_n640), .C2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n619), .B1(new_n622), .B2(new_n645), .ZN(G369));
  INV_X1    g0446(.A(G13), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n647), .A2(G1), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n214), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT27), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n648), .A2(new_n651), .A3(new_n214), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n650), .A2(G213), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(KEYINPUT86), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT86), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n650), .A2(new_n655), .A3(G213), .A4(new_n652), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n654), .A2(G343), .A3(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n575), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n657), .ZN(new_n659));
  OR3_X1    g0459(.A1(new_n575), .A2(KEYINPUT87), .A3(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(KEYINPUT87), .B1(new_n575), .B2(new_n659), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n657), .B1(new_n569), .B2(new_n574), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n575), .A2(new_n607), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(KEYINPUT88), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n662), .A2(KEYINPUT88), .A3(new_n664), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n599), .A2(new_n657), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n658), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n657), .A2(new_n583), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n641), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n599), .A2(new_n592), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n672), .B1(new_n673), .B2(new_n671), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(G330), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n668), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n670), .A2(new_n678), .ZN(G399));
  INV_X1    g0479(.A(new_n220), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(G41), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G1), .ZN(new_n683));
  OR2_X1    g0483(.A1(new_n514), .A2(G116), .ZN(new_n684));
  INV_X1    g0484(.A(new_n212), .ZN(new_n685));
  OAI22_X1  g0485(.A1(new_n683), .A2(new_n684), .B1(new_n685), .B2(new_n682), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT89), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT28), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n645), .A2(KEYINPUT29), .A3(new_n657), .ZN(new_n689));
  INV_X1    g0489(.A(new_n489), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n305), .B1(new_n479), .B2(new_n484), .ZN(new_n691));
  OAI21_X1  g0491(.A(KEYINPUT85), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  AND3_X1   g0492(.A1(new_n692), .A2(new_n635), .A3(new_n488), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n633), .B1(new_n693), .B2(new_n631), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n630), .A2(new_n531), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n638), .B2(KEYINPUT26), .ZN(new_n696));
  OAI21_X1  g0496(.A(KEYINPUT90), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n695), .A2(new_n523), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n692), .A2(new_n635), .A3(new_n488), .ZN(new_n699));
  OAI21_X1  g0499(.A(KEYINPUT26), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  AND4_X1   g0500(.A1(new_n488), .A2(new_n534), .A3(new_n490), .A4(new_n523), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n637), .B1(new_n701), .B2(new_n633), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT90), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n700), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n640), .A2(new_n643), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n697), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n659), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n689), .B1(new_n707), .B2(KEYINPUT29), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n535), .A2(new_n608), .A3(new_n539), .A4(new_n659), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n605), .A2(new_n509), .A3(new_n541), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n485), .A2(new_n590), .A3(new_n431), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(KEYINPUT30), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n596), .A2(new_n477), .A3(G179), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n714), .B1(new_n715), .B2(new_n710), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n509), .A2(G179), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n550), .A2(new_n485), .A3(new_n590), .A4(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n713), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n657), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(KEYINPUT31), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT31), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n719), .A2(new_n722), .A3(new_n657), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n709), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G330), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n708), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n688), .B1(new_n728), .B2(G1), .ZN(G364));
  NOR2_X1   g0529(.A1(new_n647), .A2(G20), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n217), .B1(new_n730), .B2(G45), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n681), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n677), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(G330), .B2(new_n674), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n213), .B1(G20), .B2(new_n305), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(G179), .A2(G200), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n214), .B1(new_n738), .B2(G190), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n443), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n214), .A2(new_n298), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n389), .A2(G179), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n743), .B1(new_n512), .B2(new_n513), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n214), .A2(G190), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n431), .A2(G200), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n744), .B1(new_n226), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n745), .A2(new_n742), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G107), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n749), .A2(new_n260), .A3(new_n752), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n214), .A2(new_n431), .A3(new_n389), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n298), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI211_X1 g0556(.A(new_n740), .B(new_n753), .C1(G68), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n745), .A2(new_n738), .ZN(new_n758));
  INV_X1    g0558(.A(G159), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XOR2_X1   g0560(.A(KEYINPUT96), .B(KEYINPUT32), .Z(new_n761));
  XNOR2_X1  g0561(.A(new_n760), .B(new_n761), .ZN(new_n762));
  AND2_X1   g0562(.A1(new_n741), .A2(new_n746), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n763), .A2(KEYINPUT94), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(KEYINPUT94), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n762), .B1(G58), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n754), .A2(G190), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(KEYINPUT95), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n768), .A2(KEYINPUT95), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n757), .B(new_n767), .C1(new_n207), .C2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n758), .ZN(new_n774));
  AOI22_X1  g0574(.A1(G283), .A2(new_n751), .B1(new_n774), .B2(G329), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n775), .B1(new_n587), .B2(new_n743), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n776), .B1(G322), .B2(new_n766), .ZN(new_n777));
  INV_X1    g0577(.A(G311), .ZN(new_n778));
  XOR2_X1   g0578(.A(KEYINPUT33), .B(G317), .Z(new_n779));
  OAI221_X1 g0579(.A(new_n394), .B1(new_n747), .B2(new_n778), .C1(new_n755), .C2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n739), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n780), .B1(G294), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G326), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n777), .B(new_n782), .C1(new_n783), .C2(new_n772), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n737), .B1(new_n773), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n733), .B(KEYINPUT91), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n680), .A2(new_n394), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n788), .A2(G355), .B1(new_n576), .B2(new_n680), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n680), .A2(new_n260), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n790), .B1(new_n685), .B2(G45), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n254), .A2(new_n271), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n789), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(G13), .A2(G33), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(G20), .ZN(new_n796));
  XOR2_X1   g0596(.A(new_n796), .B(KEYINPUT92), .Z(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n736), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n787), .B1(new_n793), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(KEYINPUT93), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n785), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n800), .A2(KEYINPUT93), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n802), .B(new_n803), .C1(new_n674), .C2(new_n797), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n735), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(G396));
  INV_X1    g0606(.A(KEYINPUT99), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n429), .A2(new_n432), .A3(new_n659), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n315), .B1(new_n414), .B2(new_n419), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n657), .B1(new_n809), .B2(new_n407), .ZN(new_n810));
  AND2_X1   g0610(.A1(new_n435), .A2(new_n810), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n807), .B(new_n808), .C1(new_n811), .C2(new_n615), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n435), .A2(new_n810), .B1(new_n429), .B2(new_n432), .ZN(new_n813));
  AND3_X1   g0613(.A1(new_n429), .A2(new_n432), .A3(new_n659), .ZN(new_n814));
  OAI21_X1  g0614(.A(KEYINPUT99), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n645), .B2(new_n657), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n657), .B1(new_n812), .B2(new_n815), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n644), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n733), .B1(new_n821), .B2(new_n726), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n726), .B2(new_n821), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n736), .A2(new_n794), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT97), .Z(new_n825));
  OAI21_X1  g0625(.A(new_n786), .B1(G77), .B2(new_n825), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n755), .B(KEYINPUT98), .Z(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n772), .ZN(new_n829));
  AOI22_X1  g0629(.A1(G283), .A2(new_n828), .B1(new_n829), .B2(G303), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n766), .A2(G294), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n750), .A2(new_n409), .B1(new_n758), .B2(new_n778), .ZN(new_n832));
  INV_X1    g0632(.A(new_n743), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n832), .B1(G107), .B2(new_n833), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n260), .B(new_n740), .C1(G116), .C2(new_n748), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n830), .A2(new_n831), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n755), .A2(new_n286), .B1(new_n759), .B2(new_n747), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(new_n766), .B2(G143), .ZN(new_n838));
  INV_X1    g0638(.A(G137), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n838), .B1(new_n772), .B2(new_n839), .ZN(new_n840));
  XOR2_X1   g0640(.A(new_n840), .B(KEYINPUT34), .Z(new_n841));
  AOI22_X1  g0641(.A1(G68), .A2(new_n751), .B1(new_n774), .B2(G132), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n394), .B1(new_n833), .B2(G50), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n842), .B(new_n843), .C1(new_n202), .C2(new_n739), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n836), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n826), .B1(new_n845), .B2(new_n736), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n795), .B2(new_n816), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n823), .A2(new_n847), .ZN(G384));
  INV_X1    g0648(.A(KEYINPUT35), .ZN(new_n849));
  OAI211_X1 g0649(.A(G116), .B(new_n215), .C1(new_n448), .C2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(new_n849), .B2(new_n448), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n851), .B(KEYINPUT36), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n212), .A2(new_n226), .A3(new_n362), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n217), .B(G13), .C1(new_n853), .C2(new_n250), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n614), .A2(new_n322), .A3(new_n659), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT104), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n366), .B1(new_n368), .B2(new_n371), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n858), .A2(new_n397), .A3(new_n282), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n351), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(KEYINPUT101), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n654), .A2(new_n656), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT101), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n859), .A2(new_n864), .A3(new_n351), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n861), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n405), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT38), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n399), .B1(new_n374), .B2(new_n386), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT37), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n374), .B2(new_n862), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n861), .A2(new_n385), .A3(new_n865), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n866), .A2(new_n874), .A3(new_n399), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n873), .B1(new_n875), .B2(KEYINPUT37), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n857), .B1(new_n869), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT39), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n875), .A2(KEYINPUT37), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT37), .B1(new_n402), .B2(new_n863), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n402), .A2(new_n385), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n880), .A2(new_n881), .A3(new_n399), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT38), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(new_n405), .B2(new_n867), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n883), .A2(KEYINPUT104), .A3(new_n885), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n877), .A2(new_n878), .A3(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT102), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n402), .A2(new_n863), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n881), .A2(new_n889), .A3(new_n399), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n882), .A2(new_n888), .B1(new_n890), .B2(KEYINPUT37), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n880), .A2(KEYINPUT102), .A3(new_n881), .A4(new_n399), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n374), .A2(new_n862), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n891), .A2(new_n892), .B1(new_n405), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(KEYINPUT103), .B1(new_n894), .B2(KEYINPUT38), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n888), .B1(new_n870), .B2(new_n872), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n896), .A2(new_n897), .A3(new_n892), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n405), .A2(new_n893), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT103), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n900), .A2(new_n901), .A3(new_n884), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n895), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n887), .A2(new_n903), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n405), .A2(new_n867), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n884), .B1(new_n876), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n883), .A2(new_n885), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT39), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n856), .B1(new_n904), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT105), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n322), .A2(new_n657), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n344), .A2(new_n348), .A3(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n348), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n322), .B(new_n657), .C1(new_n614), .C2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT100), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n917), .B1(new_n820), .B2(new_n808), .ZN(new_n918));
  AOI211_X1 g0718(.A(KEYINPUT100), .B(new_n814), .C1(new_n644), .C2(new_n819), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n916), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AND2_X1   g0720(.A1(new_n906), .A2(new_n907), .ZN(new_n921));
  OAI22_X1  g0721(.A1(new_n920), .A2(new_n921), .B1(new_n611), .B2(new_n863), .ZN(new_n922));
  NOR3_X1   g0722(.A1(new_n910), .A2(new_n911), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n901), .B1(new_n900), .B2(new_n884), .ZN(new_n924));
  AOI211_X1 g0724(.A(KEYINPUT103), .B(KEYINPUT38), .C1(new_n898), .C2(new_n899), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n877), .A2(new_n886), .A3(new_n878), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n909), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n856), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n611), .A2(new_n863), .ZN(new_n931));
  INV_X1    g0731(.A(new_n916), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n820), .A2(new_n808), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT100), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n820), .A2(new_n917), .A3(new_n808), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n931), .B1(new_n936), .B2(new_n908), .ZN(new_n937));
  AOI21_X1  g0737(.A(KEYINPUT105), .B1(new_n930), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n923), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n619), .B1(new_n708), .B2(new_n622), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n939), .B(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n916), .A2(new_n816), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(new_n709), .B2(new_n724), .ZN(new_n943));
  AOI21_X1  g0743(.A(KEYINPUT40), .B1(new_n908), .B2(new_n943), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n877), .B(new_n886), .C1(new_n924), .C2(new_n925), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n943), .A2(KEYINPUT40), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n944), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n437), .A2(new_n725), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n676), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n948), .B2(new_n949), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n941), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n217), .B2(new_n730), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n941), .A2(new_n951), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n855), .B1(new_n953), .B2(new_n954), .ZN(G367));
  INV_X1    g0755(.A(KEYINPUT108), .ZN(new_n956));
  AND3_X1   g0756(.A1(new_n662), .A2(KEYINPUT88), .A3(new_n664), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n669), .B1(new_n957), .B2(new_n665), .ZN(new_n958));
  INV_X1    g0758(.A(new_n658), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n488), .A2(new_n657), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n492), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n693), .A2(new_n657), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n958), .A2(new_n959), .A3(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT45), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n964), .A2(new_n965), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n958), .A2(new_n959), .ZN(new_n968));
  INV_X1    g0768(.A(new_n963), .ZN(new_n969));
  AOI21_X1  g0769(.A(KEYINPUT44), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT44), .ZN(new_n971));
  AOI211_X1 g0771(.A(new_n971), .B(new_n963), .C1(new_n958), .C2(new_n959), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n966), .A2(new_n967), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n678), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n666), .B(new_n667), .C1(new_n599), .C2(new_n657), .ZN(new_n976));
  AND3_X1   g0776(.A1(new_n976), .A2(new_n677), .A3(new_n958), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n677), .B1(new_n976), .B2(new_n958), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n728), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n971), .B1(new_n670), .B2(new_n963), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n968), .A2(KEYINPUT44), .A3(new_n969), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n964), .B(new_n965), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n984), .A2(new_n985), .A3(new_n678), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n975), .A2(new_n981), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(KEYINPUT106), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT106), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n975), .A2(new_n981), .A3(new_n986), .A4(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n727), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n681), .B(KEYINPUT41), .Z(new_n992));
  OAI21_X1  g0792(.A(new_n731), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n657), .A2(new_n623), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n695), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(new_n631), .B2(new_n994), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT43), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n668), .A2(new_n669), .A3(new_n963), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n999), .A2(KEYINPUT42), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n963), .A2(new_n551), .A3(new_n642), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n657), .B1(new_n1001), .B2(new_n491), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(new_n999), .B2(KEYINPUT42), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n998), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n996), .A2(new_n997), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n974), .A2(new_n963), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1006), .B(new_n1007), .Z(new_n1008));
  NAND2_X1  g0808(.A1(new_n993), .A2(new_n1008), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n240), .A2(new_n790), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n799), .B1(new_n220), .B2(new_n521), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(G159), .A2(new_n828), .B1(new_n829), .B2(G143), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n766), .A2(G150), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n743), .A2(new_n202), .B1(new_n747), .B2(new_n207), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(G137), .B2(new_n774), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n739), .A2(new_n203), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n394), .B(new_n1016), .C1(new_n226), .C2(new_n751), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1012), .A2(new_n1013), .A3(new_n1015), .A4(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n833), .A2(G116), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT46), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n1019), .A2(new_n1020), .B1(new_n423), .B2(new_n739), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(new_n1020), .B2(new_n1019), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(G283), .A2(new_n748), .B1(new_n774), .B2(G317), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n751), .A2(G97), .ZN(new_n1024));
  AND3_X1   g0824(.A1(new_n1023), .A2(new_n394), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n766), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1022), .B(new_n1025), .C1(new_n587), .C2(new_n1026), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n827), .A2(new_n543), .B1(new_n772), .B2(new_n778), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1018), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT47), .Z(new_n1030));
  OAI221_X1 g0830(.A(new_n786), .B1(new_n1010), .B2(new_n1011), .C1(new_n1030), .C2(new_n737), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT107), .Z(new_n1032));
  AND2_X1   g0832(.A1(new_n996), .A2(new_n798), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n956), .B1(new_n1009), .B2(new_n1035), .ZN(new_n1036));
  AOI211_X1 g0836(.A(KEYINPUT108), .B(new_n1034), .C1(new_n993), .C2(new_n1008), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1036), .A2(new_n1037), .ZN(G387));
  NAND2_X1  g0838(.A1(new_n979), .A2(new_n732), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n790), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n245), .B2(G45), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n684), .B2(new_n788), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n284), .A2(G50), .ZN(new_n1043));
  XOR2_X1   g0843(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n1044));
  XNOR2_X1  g0844(.A(new_n1043), .B(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n271), .B1(new_n203), .B2(new_n208), .ZN(new_n1046));
  NOR3_X1   g0846(.A1(new_n1045), .A2(new_n684), .A3(new_n1046), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n1042), .A2(new_n1047), .B1(G107), .B2(new_n220), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n787), .B1(new_n1048), .B2(new_n799), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1026), .A2(new_n207), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n772), .A2(new_n759), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n756), .A2(new_n415), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n521), .A2(new_n739), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1052), .A2(new_n1054), .A3(new_n260), .A4(new_n1024), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n833), .A2(new_n226), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(KEYINPUT110), .B(G150), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1056), .B1(new_n203), .B2(new_n747), .C1(new_n758), .C2(new_n1057), .ZN(new_n1058));
  NOR4_X1   g0858(.A1(new_n1050), .A2(new_n1051), .A3(new_n1055), .A4(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n829), .A2(G322), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n766), .A2(G317), .B1(G303), .B2(new_n748), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1060), .B(new_n1061), .C1(new_n778), .C2(new_n827), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT48), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n833), .A2(G294), .B1(new_n781), .B2(G283), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT49), .Z(new_n1068));
  OR2_X1    g0868(.A1(new_n1068), .A2(KEYINPUT111), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n394), .B1(new_n758), .B2(new_n783), .C1(new_n576), .C2(new_n750), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n1068), .B2(KEYINPUT111), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1059), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1049), .B1(new_n668), .B2(new_n797), .C1(new_n1072), .C2(new_n737), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n980), .A2(new_n681), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n979), .A2(new_n728), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1039), .B(new_n1073), .C1(new_n1074), .C2(new_n1075), .ZN(G393));
  NAND2_X1  g0876(.A1(new_n988), .A2(new_n990), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n975), .A2(new_n986), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1077), .B(new_n681), .C1(new_n981), .C2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(KEYINPUT112), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT112), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n731), .B1(new_n1078), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n969), .A2(new_n798), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n799), .B1(new_n443), .B2(new_n220), .C1(new_n249), .C2(new_n1040), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n786), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n1026), .A2(new_n759), .B1(new_n772), .B2(new_n286), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT51), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(G68), .A2(new_n833), .B1(new_n774), .B2(G143), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1089), .B(new_n260), .C1(new_n409), .C2(new_n750), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT113), .Z(new_n1091));
  OAI22_X1  g0891(.A1(new_n747), .A2(new_n284), .B1(new_n739), .B2(new_n208), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n828), .B2(G50), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1088), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1094));
  OR2_X1    g0894(.A1(new_n1094), .A2(KEYINPUT114), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n829), .A2(G317), .B1(G311), .B2(new_n766), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT52), .Z(new_n1097));
  AOI22_X1  g0897(.A1(G294), .A2(new_n748), .B1(new_n774), .B2(G322), .ZN(new_n1098));
  INV_X1    g0898(.A(G283), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1098), .B1(new_n1099), .B2(new_n743), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n752), .B(new_n394), .C1(new_n576), .C2(new_n739), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n1100), .B(new_n1101), .C1(new_n828), .C2(G303), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1097), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1094), .A2(KEYINPUT114), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1095), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1086), .B1(new_n1105), .B2(new_n736), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1081), .A2(new_n1083), .B1(new_n1084), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1080), .A2(new_n1107), .ZN(G390));
  NAND2_X1  g0908(.A1(new_n920), .A2(new_n856), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1109), .A2(new_n909), .A3(new_n904), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n706), .A2(new_n659), .A3(new_n816), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n808), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n916), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1113), .A2(new_n856), .A3(new_n945), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1110), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n676), .B1(new_n709), .B2(new_n724), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1116), .A2(new_n816), .A3(new_n916), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1110), .A2(new_n1114), .A3(new_n1117), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n932), .B1(new_n726), .B2(new_n817), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n1117), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n919), .B2(new_n918), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1122), .A2(new_n808), .A3(new_n1117), .A4(new_n1111), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n437), .A2(new_n1116), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1127), .B(new_n619), .C1(new_n708), .C2(new_n622), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n682), .B1(new_n1121), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT115), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n1110), .A2(new_n1117), .A3(new_n1114), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1117), .B1(new_n1110), .B2(new_n1114), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1128), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1132), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1119), .A2(new_n1136), .A3(new_n1132), .A4(new_n1120), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1131), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT116), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1119), .A2(new_n732), .A3(new_n1120), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n825), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n787), .B1(new_n284), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(G132), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1026), .A2(new_n1146), .ZN(new_n1147));
  OR3_X1    g0947(.A1(new_n743), .A2(new_n1057), .A3(KEYINPUT53), .ZN(new_n1148));
  OAI21_X1  g0948(.A(KEYINPUT53), .B1(new_n743), .B2(new_n1057), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1148), .B(new_n1149), .C1(new_n759), .C2(new_n739), .ZN(new_n1150));
  INV_X1    g0950(.A(G125), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n260), .B1(new_n758), .B2(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(KEYINPUT54), .B(G143), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n1153), .A2(new_n747), .B1(new_n750), .B2(new_n207), .ZN(new_n1154));
  NOR4_X1   g0954(.A1(new_n1147), .A2(new_n1150), .A3(new_n1152), .A4(new_n1154), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(G137), .A2(new_n828), .B1(new_n829), .B2(G128), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n394), .B1(new_n739), .B2(new_n208), .C1(new_n203), .C2(new_n750), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(G87), .A2(new_n833), .B1(new_n748), .B2(G97), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n543), .B2(new_n758), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n1157), .B(new_n1159), .C1(G116), .C2(new_n766), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G107), .A2(new_n828), .B1(new_n829), .B2(G283), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n1155), .A2(new_n1156), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1145), .B1(new_n737), .B2(new_n1162), .C1(new_n928), .C2(new_n795), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1143), .A2(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT117), .ZN(new_n1165));
  OAI211_X1 g0965(.A(KEYINPUT116), .B(new_n1131), .C1(new_n1137), .C2(new_n1139), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1142), .A2(new_n1165), .A3(new_n1166), .ZN(G378));
  INV_X1    g0967(.A(KEYINPUT40), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n725), .A2(new_n816), .A3(new_n916), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1168), .B1(new_n921), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n877), .A2(new_n886), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(new_n902), .B2(new_n895), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1170), .B(G330), .C1(new_n1172), .C2(new_n946), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n297), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n308), .A2(new_n1174), .A3(new_n863), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n304), .B(new_n307), .C1(new_n297), .C2(new_n862), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1175), .A2(new_n1176), .A3(new_n1178), .ZN(new_n1181));
  AND3_X1   g0981(.A1(new_n1180), .A2(KEYINPUT118), .A3(new_n1181), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1173), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1180), .A2(KEYINPUT118), .A3(new_n1181), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n948), .B2(G330), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n923), .A2(new_n938), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1173), .A2(new_n1182), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n948), .A2(G330), .A3(new_n1184), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(KEYINPUT119), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n911), .B1(new_n910), .B2(new_n922), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n930), .A2(KEYINPUT105), .A3(new_n937), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1191), .A2(new_n1192), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1186), .A2(new_n1190), .A3(new_n1193), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1189), .B(KEYINPUT119), .C1(new_n938), .C2(new_n923), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1180), .A2(new_n794), .A3(new_n1181), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n824), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n733), .B1(G50), .B2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n260), .A2(G41), .ZN(new_n1200));
  AOI211_X1 g1000(.A(G50), .B(new_n1200), .C1(new_n257), .C2(new_n270), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n750), .A2(new_n202), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n413), .B2(new_n748), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n1099), .B2(new_n758), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(G107), .B2(new_n766), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1056), .A2(new_n1200), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1016), .B(new_n1206), .C1(G97), .C2(new_n756), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1205), .B(new_n1207), .C1(new_n576), .C2(new_n772), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT58), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1201), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1153), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n833), .A2(new_n1211), .B1(new_n748), .B2(G137), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1212), .B1(new_n1146), .B2(new_n755), .C1(new_n286), .C2(new_n739), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n772), .A2(new_n1151), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1213), .B(new_n1214), .C1(G128), .C2(new_n766), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT59), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n257), .B(new_n270), .C1(new_n750), .C2(new_n759), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(G124), .B2(new_n774), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1219), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1210), .B1(new_n1209), .B2(new_n1208), .C1(new_n1217), .C2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1199), .B1(new_n1221), .B2(new_n736), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1196), .A2(new_n732), .B1(new_n1197), .B2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1129), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1224));
  AOI21_X1  g1024(.A(KEYINPUT57), .B1(new_n1224), .B2(new_n1196), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1119), .A2(new_n1136), .A3(new_n1120), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(KEYINPUT115), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1128), .B1(new_n1227), .B2(new_n1138), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1186), .A2(KEYINPUT57), .A3(new_n1193), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n681), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1223), .B1(new_n1225), .B2(new_n1230), .ZN(G375));
  NOR2_X1   g1031(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1232));
  NOR3_X1   g1032(.A1(new_n1232), .A2(new_n992), .A3(new_n1136), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1126), .A2(new_n732), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n786), .B1(G68), .B2(new_n825), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n260), .B(new_n1053), .C1(G77), .C2(new_n751), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n743), .A2(new_n443), .B1(new_n758), .B2(new_n587), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(G107), .B2(new_n748), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1236), .B(new_n1238), .C1(new_n1099), .C2(new_n1026), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n827), .A2(new_n576), .B1(new_n772), .B2(new_n543), .ZN(new_n1240));
  INV_X1    g1040(.A(G128), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n747), .A2(new_n286), .B1(new_n758), .B2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(G159), .B2(new_n833), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n394), .B(new_n1202), .C1(G50), .C2(new_n781), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1243), .B(new_n1244), .C1(new_n1026), .C2(new_n839), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n827), .A2(new_n1153), .B1(new_n772), .B2(new_n1146), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n1239), .A2(new_n1240), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1235), .B1(new_n1247), .B2(new_n736), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(new_n916), .B2(new_n795), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1234), .A2(new_n1249), .ZN(new_n1250));
  OR2_X1    g1050(.A1(new_n1233), .A2(new_n1250), .ZN(G381));
  OR3_X1    g1051(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1252));
  NOR3_X1   g1052(.A1(G390), .A2(G381), .A3(new_n1252), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1253), .B(KEYINPUT120), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT57), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1255), .B1(new_n1256), .B2(new_n1228), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1229), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n682), .B1(new_n1224), .B2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1257), .A2(new_n1259), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1140), .A2(new_n1143), .A3(new_n1163), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1260), .A2(new_n1223), .A3(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  AND2_X1   g1063(.A1(new_n1254), .A2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1253), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT120), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1264), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT121), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1264), .A2(KEYINPUT121), .A3(new_n1267), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(G407));
  INV_X1    g1072(.A(G213), .ZN(new_n1273));
  OR2_X1    g1073(.A1(new_n1273), .A2(G343), .ZN(new_n1274));
  XOR2_X1   g1074(.A(new_n1274), .B(KEYINPUT122), .Z(new_n1275));
  AOI21_X1  g1075(.A(new_n1273), .B1(new_n1263), .B2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(KEYINPUT121), .B1(new_n1264), .B2(new_n1267), .ZN(new_n1277));
  AND4_X1   g1077(.A1(KEYINPUT121), .A2(new_n1267), .A3(new_n1263), .A4(new_n1254), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1276), .B1(new_n1277), .B2(new_n1278), .ZN(G409));
  XNOR2_X1  g1079(.A(G393), .B(new_n805), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1080), .B(new_n1107), .C1(KEYINPUT108), .C2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(G390), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1281), .B1(new_n1282), .B2(new_n1280), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1009), .A2(new_n1035), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1283), .B(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1275), .A2(G2897), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1130), .A2(KEYINPUT60), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1232), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1124), .A2(new_n1128), .A3(new_n1125), .A4(KEYINPUT60), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n681), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1250), .B1(new_n1290), .B2(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(KEYINPUT124), .B1(new_n1294), .B2(G384), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1250), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1232), .B1(KEYINPUT60), .B2(new_n1130), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1296), .B1(new_n1297), .B2(new_n1292), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT124), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1298), .A2(new_n1299), .A3(new_n823), .A4(new_n847), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1294), .A2(KEYINPUT123), .A3(G384), .ZN(new_n1301));
  OAI211_X1 g1101(.A(G384), .B(new_n1296), .C1(new_n1297), .C2(new_n1292), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT123), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  AOI22_X1  g1104(.A1(new_n1295), .A2(new_n1300), .B1(new_n1301), .B2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1275), .ZN(new_n1306));
  OR2_X1    g1106(.A1(new_n1306), .A2(KEYINPUT125), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1287), .B1(new_n1305), .B2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1301), .A2(new_n1304), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1295), .A2(new_n1300), .ZN(new_n1310));
  AND4_X1   g1110(.A1(new_n1309), .A2(new_n1310), .A3(new_n1287), .A4(new_n1307), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1308), .A2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1260), .A2(G378), .A3(new_n1223), .ZN(new_n1313));
  NOR3_X1   g1113(.A1(new_n1256), .A2(new_n1228), .A3(new_n992), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1186), .A2(new_n732), .A3(new_n1193), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1197), .A2(new_n1222), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1261), .B1(new_n1314), .B2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1313), .A2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(new_n1306), .ZN(new_n1320));
  AOI21_X1  g1120(.A(KEYINPUT61), .B1(new_n1312), .B2(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1319), .A2(new_n1306), .A3(new_n1305), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(KEYINPUT62), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1321), .A2(new_n1323), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1322), .A2(KEYINPUT62), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1286), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT63), .ZN(new_n1327));
  OR2_X1    g1127(.A1(new_n1322), .A2(new_n1327), .ZN(new_n1328));
  XNOR2_X1  g1128(.A(new_n1283), .B(new_n1284), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1322), .A2(new_n1327), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1328), .A2(new_n1329), .A3(new_n1321), .A4(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1326), .A2(new_n1331), .ZN(G405));
  INV_X1    g1132(.A(KEYINPUT126), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(G375), .A2(new_n1261), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1310), .A2(new_n1309), .ZN(new_n1335));
  AND3_X1   g1135(.A1(new_n1334), .A2(new_n1313), .A3(new_n1335), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1335), .B1(new_n1334), .B2(new_n1313), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1333), .B1(new_n1336), .B2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1286), .A2(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT127), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1340), .B1(new_n1341), .B2(KEYINPUT126), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1334), .A2(new_n1313), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1343), .A2(new_n1305), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1334), .A2(new_n1313), .A3(new_n1335), .ZN(new_n1345));
  NAND4_X1  g1145(.A1(new_n1344), .A2(KEYINPUT126), .A3(new_n1340), .A4(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1346), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1339), .B1(new_n1342), .B2(new_n1347), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1344), .A2(KEYINPUT126), .A3(new_n1345), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1349), .A2(KEYINPUT127), .ZN(new_n1350));
  NAND4_X1  g1150(.A1(new_n1350), .A2(new_n1286), .A3(new_n1346), .A4(new_n1338), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1348), .A2(new_n1351), .ZN(G402));
endmodule


