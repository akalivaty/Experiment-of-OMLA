

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586;

  XNOR2_X1 U322 ( .A(n467), .B(KEYINPUT37), .ZN(n468) );
  NOR2_X1 U323 ( .A1(n480), .A2(n583), .ZN(n290) );
  AND2_X1 U324 ( .A1(G227GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U325 ( .A(n438), .B(n291), .ZN(n439) );
  XNOR2_X1 U326 ( .A(n319), .B(KEYINPUT65), .ZN(n320) );
  INV_X1 U327 ( .A(KEYINPUT102), .ZN(n467) );
  XNOR2_X1 U328 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U329 ( .A(n321), .B(n320), .ZN(n327) );
  XNOR2_X1 U330 ( .A(n469), .B(n468), .ZN(n512) );
  XNOR2_X1 U331 ( .A(n554), .B(KEYINPUT78), .ZN(n561) );
  XNOR2_X1 U332 ( .A(n446), .B(n445), .ZN(n526) );
  XNOR2_X1 U333 ( .A(n449), .B(G176GAT), .ZN(n450) );
  XNOR2_X1 U334 ( .A(n471), .B(G43GAT), .ZN(n472) );
  XNOR2_X1 U335 ( .A(n451), .B(n450), .ZN(G1349GAT) );
  XNOR2_X1 U336 ( .A(n473), .B(n472), .ZN(G1330GAT) );
  XOR2_X1 U337 ( .A(KEYINPUT15), .B(KEYINPUT82), .Z(n293) );
  XNOR2_X1 U338 ( .A(G64GAT), .B(KEYINPUT80), .ZN(n292) );
  XNOR2_X1 U339 ( .A(n293), .B(n292), .ZN(n308) );
  XOR2_X1 U340 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n295) );
  NAND2_X1 U341 ( .A1(G231GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U342 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U343 ( .A(n296), .B(KEYINPUT81), .Z(n300) );
  XNOR2_X1 U344 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n297) );
  XNOR2_X1 U345 ( .A(n297), .B(KEYINPUT70), .ZN(n344) );
  XNOR2_X1 U346 ( .A(G8GAT), .B(G211GAT), .ZN(n298) );
  XNOR2_X1 U347 ( .A(n298), .B(KEYINPUT79), .ZN(n379) );
  XNOR2_X1 U348 ( .A(n344), .B(n379), .ZN(n299) );
  XNOR2_X1 U349 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U350 ( .A(G15GAT), .B(G127GAT), .Z(n432) );
  XOR2_X1 U351 ( .A(G22GAT), .B(G155GAT), .Z(n416) );
  XOR2_X1 U352 ( .A(n432), .B(n416), .Z(n302) );
  XNOR2_X1 U353 ( .A(G183GAT), .B(G71GAT), .ZN(n301) );
  XNOR2_X1 U354 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U355 ( .A(n304), .B(n303), .Z(n306) );
  XNOR2_X1 U356 ( .A(G1GAT), .B(G78GAT), .ZN(n305) );
  XNOR2_X1 U357 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U358 ( .A(n308), .B(n307), .Z(n580) );
  XOR2_X1 U359 ( .A(KEYINPUT9), .B(KEYINPUT77), .Z(n310) );
  XNOR2_X1 U360 ( .A(KEYINPUT11), .B(KEYINPUT10), .ZN(n309) );
  XNOR2_X1 U361 ( .A(n310), .B(n309), .ZN(n314) );
  XOR2_X1 U362 ( .A(G99GAT), .B(G85GAT), .Z(n329) );
  XOR2_X1 U363 ( .A(KEYINPUT76), .B(KEYINPUT66), .Z(n311) );
  XNOR2_X1 U364 ( .A(n329), .B(n311), .ZN(n312) );
  XOR2_X1 U365 ( .A(G162GAT), .B(G106GAT), .Z(n417) );
  XNOR2_X1 U366 ( .A(n312), .B(n417), .ZN(n313) );
  XOR2_X1 U367 ( .A(n314), .B(n313), .Z(n316) );
  NAND2_X1 U368 ( .A1(G232GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U369 ( .A(n316), .B(n315), .ZN(n321) );
  XOR2_X1 U370 ( .A(G92GAT), .B(G218GAT), .Z(n318) );
  XNOR2_X1 U371 ( .A(G36GAT), .B(G190GAT), .ZN(n317) );
  XNOR2_X1 U372 ( .A(n318), .B(n317), .ZN(n373) );
  XOR2_X1 U373 ( .A(G134GAT), .B(n373), .Z(n319) );
  XNOR2_X1 U374 ( .A(G43GAT), .B(KEYINPUT68), .ZN(n322) );
  XNOR2_X1 U375 ( .A(n322), .B(G29GAT), .ZN(n323) );
  XOR2_X1 U376 ( .A(n323), .B(KEYINPUT7), .Z(n325) );
  XNOR2_X1 U377 ( .A(G50GAT), .B(KEYINPUT8), .ZN(n324) );
  XNOR2_X1 U378 ( .A(n325), .B(n324), .ZN(n350) );
  INV_X1 U379 ( .A(n350), .ZN(n326) );
  XNOR2_X1 U380 ( .A(n327), .B(n326), .ZN(n554) );
  XNOR2_X1 U381 ( .A(KEYINPUT36), .B(n561), .ZN(n583) );
  NOR2_X1 U382 ( .A1(n580), .A2(n583), .ZN(n328) );
  XNOR2_X1 U383 ( .A(n328), .B(KEYINPUT45), .ZN(n363) );
  XOR2_X1 U384 ( .A(G176GAT), .B(G64GAT), .Z(n376) );
  XOR2_X1 U385 ( .A(n376), .B(n329), .Z(n331) );
  XNOR2_X1 U386 ( .A(G106GAT), .B(G92GAT), .ZN(n330) );
  XNOR2_X1 U387 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U388 ( .A(KEYINPUT32), .B(KEYINPUT75), .Z(n333) );
  NAND2_X1 U389 ( .A1(G230GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U390 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U391 ( .A(n335), .B(n334), .Z(n337) );
  XOR2_X1 U392 ( .A(G120GAT), .B(G71GAT), .Z(n433) );
  XNOR2_X1 U393 ( .A(n433), .B(KEYINPUT33), .ZN(n336) );
  XNOR2_X1 U394 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U395 ( .A(KEYINPUT31), .B(KEYINPUT74), .Z(n339) );
  XNOR2_X1 U396 ( .A(G204GAT), .B(KEYINPUT73), .ZN(n338) );
  XNOR2_X1 U397 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U398 ( .A(n341), .B(n340), .Z(n346) );
  XOR2_X1 U399 ( .A(G78GAT), .B(G148GAT), .Z(n343) );
  XNOR2_X1 U400 ( .A(KEYINPUT71), .B(KEYINPUT72), .ZN(n342) );
  XNOR2_X1 U401 ( .A(n343), .B(n342), .ZN(n413) );
  XNOR2_X1 U402 ( .A(n413), .B(n344), .ZN(n345) );
  XNOR2_X1 U403 ( .A(n346), .B(n345), .ZN(n575) );
  XOR2_X1 U404 ( .A(G141GAT), .B(G197GAT), .Z(n348) );
  XNOR2_X1 U405 ( .A(G169GAT), .B(G15GAT), .ZN(n347) );
  XNOR2_X1 U406 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U407 ( .A(n350), .B(n349), .ZN(n360) );
  XOR2_X1 U408 ( .A(G1GAT), .B(KEYINPUT29), .Z(n352) );
  XNOR2_X1 U409 ( .A(G22GAT), .B(G8GAT), .ZN(n351) );
  XNOR2_X1 U410 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U411 ( .A(G113GAT), .B(G36GAT), .Z(n354) );
  XNOR2_X1 U412 ( .A(KEYINPUT67), .B(KEYINPUT30), .ZN(n353) );
  XNOR2_X1 U413 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U414 ( .A(n356), .B(n355), .Z(n358) );
  NAND2_X1 U415 ( .A1(G229GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U416 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U417 ( .A(n360), .B(n359), .ZN(n572) );
  XOR2_X1 U418 ( .A(n572), .B(KEYINPUT69), .Z(n558) );
  INV_X1 U419 ( .A(n558), .ZN(n361) );
  NOR2_X1 U420 ( .A1(n575), .A2(n361), .ZN(n362) );
  AND2_X1 U421 ( .A1(n363), .A2(n362), .ZN(n365) );
  INV_X1 U422 ( .A(KEYINPUT113), .ZN(n364) );
  XNOR2_X1 U423 ( .A(n365), .B(n364), .ZN(n371) );
  XNOR2_X1 U424 ( .A(KEYINPUT112), .B(n580), .ZN(n535) );
  NAND2_X1 U425 ( .A1(n554), .A2(n535), .ZN(n368) );
  XNOR2_X1 U426 ( .A(KEYINPUT41), .B(n575), .ZN(n547) );
  NOR2_X1 U427 ( .A1(n572), .A2(n547), .ZN(n366) );
  XNOR2_X1 U428 ( .A(n366), .B(KEYINPUT46), .ZN(n367) );
  NOR2_X1 U429 ( .A1(n368), .A2(n367), .ZN(n369) );
  XOR2_X1 U430 ( .A(KEYINPUT47), .B(n369), .Z(n370) );
  NOR2_X1 U431 ( .A1(n371), .A2(n370), .ZN(n372) );
  XNOR2_X1 U432 ( .A(n372), .B(KEYINPUT48), .ZN(n527) );
  XNOR2_X1 U433 ( .A(n373), .B(KEYINPUT97), .ZN(n374) );
  XNOR2_X1 U434 ( .A(n374), .B(KEYINPUT96), .ZN(n375) );
  XOR2_X1 U435 ( .A(n376), .B(n375), .Z(n378) );
  NAND2_X1 U436 ( .A1(G226GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U437 ( .A(n378), .B(n377), .ZN(n380) );
  XNOR2_X1 U438 ( .A(n380), .B(n379), .ZN(n388) );
  XNOR2_X1 U439 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n381) );
  XNOR2_X1 U440 ( .A(n381), .B(KEYINPUT17), .ZN(n382) );
  XOR2_X1 U441 ( .A(n382), .B(KEYINPUT87), .Z(n384) );
  XNOR2_X1 U442 ( .A(G169GAT), .B(G183GAT), .ZN(n383) );
  XNOR2_X1 U443 ( .A(n384), .B(n383), .ZN(n446) );
  XOR2_X1 U444 ( .A(G204GAT), .B(KEYINPUT21), .Z(n386) );
  XNOR2_X1 U445 ( .A(G197GAT), .B(KEYINPUT92), .ZN(n385) );
  XNOR2_X1 U446 ( .A(n386), .B(n385), .ZN(n425) );
  XOR2_X1 U447 ( .A(n446), .B(n425), .Z(n387) );
  XNOR2_X1 U448 ( .A(n388), .B(n387), .ZN(n515) );
  XNOR2_X1 U449 ( .A(n515), .B(KEYINPUT120), .ZN(n389) );
  NOR2_X1 U450 ( .A1(n527), .A2(n389), .ZN(n390) );
  XNOR2_X1 U451 ( .A(KEYINPUT54), .B(n390), .ZN(n568) );
  XOR2_X1 U452 ( .A(G85GAT), .B(G162GAT), .Z(n392) );
  XNOR2_X1 U453 ( .A(G29GAT), .B(G120GAT), .ZN(n391) );
  XNOR2_X1 U454 ( .A(n392), .B(n391), .ZN(n396) );
  XOR2_X1 U455 ( .A(G155GAT), .B(G148GAT), .Z(n394) );
  XNOR2_X1 U456 ( .A(G1GAT), .B(G127GAT), .ZN(n393) );
  XNOR2_X1 U457 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U458 ( .A(n396), .B(n395), .Z(n401) );
  XOR2_X1 U459 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n398) );
  NAND2_X1 U460 ( .A1(G225GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U461 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U462 ( .A(KEYINPUT94), .B(n399), .ZN(n400) );
  XNOR2_X1 U463 ( .A(n401), .B(n400), .ZN(n405) );
  XOR2_X1 U464 ( .A(KEYINPUT5), .B(KEYINPUT95), .Z(n403) );
  XNOR2_X1 U465 ( .A(G57GAT), .B(KEYINPUT4), .ZN(n402) );
  XNOR2_X1 U466 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U467 ( .A(n405), .B(n404), .Z(n411) );
  XOR2_X1 U468 ( .A(KEYINPUT85), .B(KEYINPUT0), .Z(n407) );
  XNOR2_X1 U469 ( .A(G113GAT), .B(G134GAT), .ZN(n406) );
  XNOR2_X1 U470 ( .A(n407), .B(n406), .ZN(n442) );
  XOR2_X1 U471 ( .A(KEYINPUT2), .B(KEYINPUT93), .Z(n409) );
  XNOR2_X1 U472 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n408) );
  XNOR2_X1 U473 ( .A(n409), .B(n408), .ZN(n412) );
  XNOR2_X1 U474 ( .A(n442), .B(n412), .ZN(n410) );
  XNOR2_X1 U475 ( .A(n411), .B(n410), .ZN(n567) );
  INV_X1 U476 ( .A(n567), .ZN(n459) );
  XNOR2_X1 U477 ( .A(n413), .B(n412), .ZN(n429) );
  XOR2_X1 U478 ( .A(KEYINPUT91), .B(KEYINPUT22), .Z(n415) );
  XNOR2_X1 U479 ( .A(KEYINPUT23), .B(G211GAT), .ZN(n414) );
  XNOR2_X1 U480 ( .A(n415), .B(n414), .ZN(n421) );
  XOR2_X1 U481 ( .A(G218GAT), .B(n416), .Z(n419) );
  XNOR2_X1 U482 ( .A(G50GAT), .B(n417), .ZN(n418) );
  XNOR2_X1 U483 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U484 ( .A(n421), .B(n420), .Z(n423) );
  NAND2_X1 U485 ( .A1(G228GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U486 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U487 ( .A(n424), .B(KEYINPUT24), .Z(n427) );
  XNOR2_X1 U488 ( .A(n425), .B(KEYINPUT90), .ZN(n426) );
  XNOR2_X1 U489 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U490 ( .A(n429), .B(n428), .ZN(n462) );
  NOR2_X1 U491 ( .A1(n459), .A2(n462), .ZN(n430) );
  AND2_X1 U492 ( .A1(n568), .A2(n430), .ZN(n431) );
  XNOR2_X1 U493 ( .A(n431), .B(KEYINPUT55), .ZN(n447) );
  XOR2_X1 U494 ( .A(G99GAT), .B(G190GAT), .Z(n435) );
  XNOR2_X1 U495 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U496 ( .A(n435), .B(n434), .ZN(n440) );
  XOR2_X1 U497 ( .A(KEYINPUT64), .B(KEYINPUT86), .Z(n437) );
  XNOR2_X1 U498 ( .A(G43GAT), .B(KEYINPUT88), .ZN(n436) );
  XNOR2_X1 U499 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U500 ( .A(n441), .B(G176GAT), .ZN(n444) );
  XOR2_X1 U501 ( .A(n442), .B(KEYINPUT20), .Z(n443) );
  XNOR2_X1 U502 ( .A(n444), .B(n443), .ZN(n445) );
  NOR2_X1 U503 ( .A1(n447), .A2(n526), .ZN(n448) );
  XNOR2_X1 U504 ( .A(KEYINPUT121), .B(n448), .ZN(n560) );
  NOR2_X1 U505 ( .A1(n560), .A2(n547), .ZN(n451) );
  XNOR2_X1 U506 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n449) );
  XNOR2_X1 U507 ( .A(n515), .B(KEYINPUT98), .ZN(n452) );
  XNOR2_X1 U508 ( .A(n452), .B(KEYINPUT27), .ZN(n461) );
  NAND2_X1 U509 ( .A1(n526), .A2(n462), .ZN(n453) );
  XNOR2_X1 U510 ( .A(n453), .B(KEYINPUT26), .ZN(n570) );
  NOR2_X1 U511 ( .A1(n461), .A2(n570), .ZN(n457) );
  NOR2_X1 U512 ( .A1(n515), .A2(n526), .ZN(n454) );
  OR2_X1 U513 ( .A1(n462), .A2(n454), .ZN(n455) );
  XNOR2_X1 U514 ( .A(KEYINPUT25), .B(n455), .ZN(n456) );
  NOR2_X1 U515 ( .A1(n457), .A2(n456), .ZN(n458) );
  NOR2_X1 U516 ( .A1(n459), .A2(n458), .ZN(n460) );
  XNOR2_X1 U517 ( .A(KEYINPUT99), .B(n460), .ZN(n465) );
  NOR2_X1 U518 ( .A1(n567), .A2(n461), .ZN(n544) );
  XOR2_X1 U519 ( .A(n462), .B(KEYINPUT28), .Z(n523) );
  NAND2_X1 U520 ( .A1(n544), .A2(n523), .ZN(n528) );
  XNOR2_X1 U521 ( .A(KEYINPUT89), .B(n526), .ZN(n463) );
  OR2_X1 U522 ( .A1(n528), .A2(n463), .ZN(n464) );
  AND2_X1 U523 ( .A1(n465), .A2(n464), .ZN(n466) );
  XOR2_X1 U524 ( .A(KEYINPUT100), .B(n466), .Z(n485) );
  INV_X1 U525 ( .A(n580), .ZN(n480) );
  AND2_X1 U526 ( .A1(n485), .A2(n290), .ZN(n469) );
  NOR2_X1 U527 ( .A1(n558), .A2(n575), .ZN(n486) );
  NAND2_X1 U528 ( .A1(n512), .A2(n486), .ZN(n470) );
  XNOR2_X1 U529 ( .A(n470), .B(KEYINPUT38), .ZN(n497) );
  NOR2_X1 U530 ( .A1(n497), .A2(n526), .ZN(n473) );
  INV_X1 U531 ( .A(KEYINPUT40), .ZN(n471) );
  INV_X1 U532 ( .A(G50GAT), .ZN(n476) );
  NOR2_X1 U533 ( .A1(n523), .A2(n497), .ZN(n474) );
  XNOR2_X1 U534 ( .A(KEYINPUT104), .B(n474), .ZN(n475) );
  XNOR2_X1 U535 ( .A(n476), .B(n475), .ZN(G1331GAT) );
  NOR2_X1 U536 ( .A1(n560), .A2(n535), .ZN(n477) );
  XNOR2_X1 U537 ( .A(KEYINPUT122), .B(n477), .ZN(n479) );
  INV_X1 U538 ( .A(G183GAT), .ZN(n478) );
  XNOR2_X1 U539 ( .A(n479), .B(n478), .ZN(G1350GAT) );
  XOR2_X1 U540 ( .A(KEYINPUT16), .B(KEYINPUT84), .Z(n482) );
  NAND2_X1 U541 ( .A1(n561), .A2(n480), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U543 ( .A(n483), .B(KEYINPUT83), .Z(n484) );
  AND2_X1 U544 ( .A1(n485), .A2(n484), .ZN(n501) );
  NAND2_X1 U545 ( .A1(n486), .A2(n501), .ZN(n492) );
  NOR2_X1 U546 ( .A1(n567), .A2(n492), .ZN(n487) );
  XOR2_X1 U547 ( .A(G1GAT), .B(n487), .Z(n488) );
  XNOR2_X1 U548 ( .A(KEYINPUT34), .B(n488), .ZN(G1324GAT) );
  NOR2_X1 U549 ( .A1(n515), .A2(n492), .ZN(n489) );
  XOR2_X1 U550 ( .A(G8GAT), .B(n489), .Z(G1325GAT) );
  NOR2_X1 U551 ( .A1(n526), .A2(n492), .ZN(n491) );
  XNOR2_X1 U552 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n491), .B(n490), .ZN(G1326GAT) );
  NOR2_X1 U554 ( .A1(n523), .A2(n492), .ZN(n494) );
  XNOR2_X1 U555 ( .A(G22GAT), .B(KEYINPUT101), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n494), .B(n493), .ZN(G1327GAT) );
  XNOR2_X1 U557 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n496) );
  NOR2_X1 U558 ( .A1(n567), .A2(n497), .ZN(n495) );
  XNOR2_X1 U559 ( .A(n496), .B(n495), .ZN(G1328GAT) );
  XNOR2_X1 U560 ( .A(G36GAT), .B(KEYINPUT103), .ZN(n499) );
  NOR2_X1 U561 ( .A1(n497), .A2(n515), .ZN(n498) );
  XNOR2_X1 U562 ( .A(n499), .B(n498), .ZN(G1329GAT) );
  INV_X1 U563 ( .A(n572), .ZN(n500) );
  NOR2_X1 U564 ( .A1(n500), .A2(n547), .ZN(n513) );
  NAND2_X1 U565 ( .A1(n513), .A2(n501), .ZN(n508) );
  NOR2_X1 U566 ( .A1(n567), .A2(n508), .ZN(n503) );
  XNOR2_X1 U567 ( .A(KEYINPUT105), .B(KEYINPUT42), .ZN(n502) );
  XNOR2_X1 U568 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(n504), .ZN(G1332GAT) );
  NOR2_X1 U570 ( .A1(n515), .A2(n508), .ZN(n505) );
  XOR2_X1 U571 ( .A(KEYINPUT106), .B(n505), .Z(n506) );
  XNOR2_X1 U572 ( .A(G64GAT), .B(n506), .ZN(G1333GAT) );
  NOR2_X1 U573 ( .A1(n526), .A2(n508), .ZN(n507) );
  XOR2_X1 U574 ( .A(G71GAT), .B(n507), .Z(G1334GAT) );
  NOR2_X1 U575 ( .A1(n523), .A2(n508), .ZN(n510) );
  XNOR2_X1 U576 ( .A(KEYINPUT107), .B(KEYINPUT43), .ZN(n509) );
  XNOR2_X1 U577 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U578 ( .A(G78GAT), .B(n511), .Z(G1335GAT) );
  NAND2_X1 U579 ( .A1(n513), .A2(n512), .ZN(n522) );
  NOR2_X1 U580 ( .A1(n567), .A2(n522), .ZN(n514) );
  XOR2_X1 U581 ( .A(G85GAT), .B(n514), .Z(G1336GAT) );
  NOR2_X1 U582 ( .A1(n515), .A2(n522), .ZN(n516) );
  XOR2_X1 U583 ( .A(KEYINPUT108), .B(n516), .Z(n517) );
  XNOR2_X1 U584 ( .A(G92GAT), .B(n517), .ZN(G1337GAT) );
  NOR2_X1 U585 ( .A1(n526), .A2(n522), .ZN(n519) );
  XNOR2_X1 U586 ( .A(G99GAT), .B(KEYINPUT109), .ZN(n518) );
  XNOR2_X1 U587 ( .A(n519), .B(n518), .ZN(G1338GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT110), .B(KEYINPUT44), .Z(n521) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(KEYINPUT111), .ZN(n520) );
  XNOR2_X1 U590 ( .A(n521), .B(n520), .ZN(n525) );
  NOR2_X1 U591 ( .A1(n523), .A2(n522), .ZN(n524) );
  XOR2_X1 U592 ( .A(n525), .B(n524), .Z(G1339GAT) );
  INV_X1 U593 ( .A(n526), .ZN(n530) );
  BUF_X1 U594 ( .A(n527), .Z(n542) );
  NOR2_X1 U595 ( .A1(n542), .A2(n528), .ZN(n529) );
  NAND2_X1 U596 ( .A1(n530), .A2(n529), .ZN(n539) );
  NOR2_X1 U597 ( .A1(n558), .A2(n539), .ZN(n531) );
  XOR2_X1 U598 ( .A(G113GAT), .B(n531), .Z(G1340GAT) );
  NOR2_X1 U599 ( .A1(n547), .A2(n539), .ZN(n533) );
  XNOR2_X1 U600 ( .A(KEYINPUT114), .B(KEYINPUT49), .ZN(n532) );
  XNOR2_X1 U601 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U602 ( .A(G120GAT), .B(n534), .ZN(G1341GAT) );
  NOR2_X1 U603 ( .A1(n535), .A2(n539), .ZN(n537) );
  XNOR2_X1 U604 ( .A(KEYINPUT50), .B(KEYINPUT115), .ZN(n536) );
  XNOR2_X1 U605 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  NOR2_X1 U607 ( .A1(n561), .A2(n539), .ZN(n541) );
  XNOR2_X1 U608 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n540) );
  XNOR2_X1 U609 ( .A(n541), .B(n540), .ZN(G1343GAT) );
  NOR2_X1 U610 ( .A1(n542), .A2(n570), .ZN(n543) );
  NAND2_X1 U611 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U612 ( .A(KEYINPUT116), .B(n545), .ZN(n553) );
  NOR2_X1 U613 ( .A1(n572), .A2(n553), .ZN(n546) );
  XOR2_X1 U614 ( .A(G141GAT), .B(n546), .Z(G1344GAT) );
  NOR2_X1 U615 ( .A1(n547), .A2(n553), .ZN(n551) );
  XOR2_X1 U616 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n549) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(KEYINPUT117), .ZN(n548) );
  XNOR2_X1 U618 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(G1345GAT) );
  NOR2_X1 U620 ( .A1(n580), .A2(n553), .ZN(n552) );
  XOR2_X1 U621 ( .A(G155GAT), .B(n552), .Z(G1346GAT) );
  XNOR2_X1 U622 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n556) );
  NOR2_X1 U623 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U625 ( .A(G162GAT), .B(n557), .ZN(G1347GAT) );
  OR2_X1 U626 ( .A1(n560), .A2(n558), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n559), .B(G169GAT), .ZN(G1348GAT) );
  NOR2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n563) );
  INV_X1 U629 ( .A(KEYINPUT58), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(G190GAT), .ZN(G1351GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n566) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n565) );
  XNOR2_X1 U634 ( .A(n566), .B(n565), .ZN(n574) );
  NAND2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(KEYINPUT123), .B(n571), .ZN(n582) );
  NOR2_X1 U638 ( .A1(n572), .A2(n582), .ZN(n573) );
  XOR2_X1 U639 ( .A(n574), .B(n573), .Z(G1352GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n578) );
  INV_X1 U641 ( .A(n582), .ZN(n576) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n579) );
  XOR2_X1 U644 ( .A(G204GAT), .B(n579), .Z(G1353GAT) );
  NOR2_X1 U645 ( .A1(n580), .A2(n582), .ZN(n581) );
  XOR2_X1 U646 ( .A(G211GAT), .B(n581), .Z(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n585) );
  XNOR2_X1 U648 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XOR2_X1 U650 ( .A(G218GAT), .B(n586), .Z(G1355GAT) );
endmodule

