

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735;

  XNOR2_X1 U367 ( .A(n427), .B(KEYINPUT19), .ZN(n562) );
  AND2_X1 U368 ( .A1(n635), .A2(n722), .ZN(n346) );
  NOR2_X2 U369 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X2 U370 ( .A1(G902), .A2(n705), .ZN(n379) );
  XNOR2_X1 U371 ( .A(n457), .B(n370), .ZN(n386) );
  NAND2_X2 U372 ( .A1(n362), .A2(n361), .ZN(n704) );
  NOR2_X1 U373 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X2 U374 ( .A1(n591), .A2(n590), .ZN(n722) );
  AND2_X1 U375 ( .A1(n526), .A2(n525), .ZN(n534) );
  XNOR2_X1 U376 ( .A(n472), .B(n471), .ZN(n528) );
  NOR2_X1 U377 ( .A1(n510), .A2(n519), .ZN(n500) );
  OR2_X1 U378 ( .A1(n575), .A2(n426), .ZN(n427) );
  XNOR2_X1 U379 ( .A(n386), .B(KEYINPUT91), .ZN(n716) );
  XNOR2_X1 U380 ( .A(n412), .B(G134), .ZN(n457) );
  XNOR2_X1 U381 ( .A(n368), .B(n367), .ZN(n412) );
  NOR2_X1 U382 ( .A1(n568), .A2(n575), .ZN(n569) );
  AND2_X1 U383 ( .A1(n530), .A2(n359), .ZN(n358) );
  OR2_X1 U384 ( .A1(n732), .A2(n357), .ZN(n356) );
  AND2_X1 U385 ( .A1(n528), .A2(KEYINPUT44), .ZN(n359) );
  XNOR2_X1 U386 ( .A(G146), .B(G101), .ZN(n374) );
  XNOR2_X1 U387 ( .A(G146), .B(G125), .ZN(n410) );
  XNOR2_X1 U388 ( .A(n371), .B(G104), .ZN(n406) );
  XNOR2_X1 U389 ( .A(G110), .B(G107), .ZN(n371) );
  XNOR2_X1 U390 ( .A(KEYINPUT12), .B(KEYINPUT11), .ZN(n440) );
  XOR2_X1 U391 ( .A(G122), .B(G113), .Z(n444) );
  XNOR2_X1 U392 ( .A(G104), .B(G143), .ZN(n443) );
  XNOR2_X1 U393 ( .A(G143), .B(KEYINPUT66), .ZN(n368) );
  NOR2_X1 U394 ( .A1(n481), .A2(n480), .ZN(n482) );
  OR2_X1 U395 ( .A1(n615), .A2(n418), .ZN(n423) );
  XNOR2_X1 U396 ( .A(n462), .B(n461), .ZN(n516) );
  XNOR2_X1 U397 ( .A(n451), .B(KEYINPUT13), .ZN(n515) );
  XNOR2_X1 U398 ( .A(G475), .B(n450), .ZN(n451) );
  BUF_X1 U399 ( .A(n499), .Z(n658) );
  INV_X1 U400 ( .A(KEYINPUT84), .ZN(n357) );
  XNOR2_X1 U401 ( .A(G113), .B(G101), .ZN(n354) );
  XNOR2_X1 U402 ( .A(KEYINPUT70), .B(KEYINPUT71), .ZN(n355) );
  XNOR2_X1 U403 ( .A(n387), .B(G472), .ZN(n665) );
  XNOR2_X1 U404 ( .A(n403), .B(n402), .ZN(n550) );
  XNOR2_X1 U405 ( .A(n587), .B(n586), .ZN(n591) );
  XNOR2_X1 U406 ( .A(n353), .B(n351), .ZN(n407) );
  XNOR2_X1 U407 ( .A(n352), .B(KEYINPUT3), .ZN(n351) );
  XNOR2_X1 U408 ( .A(n355), .B(n354), .ZN(n353) );
  XNOR2_X1 U409 ( .A(G119), .B(G116), .ZN(n352) );
  XNOR2_X1 U410 ( .A(G128), .B(G119), .ZN(n388) );
  XNOR2_X1 U411 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U412 ( .A(n406), .B(n373), .ZN(n376) );
  XNOR2_X1 U413 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n409) );
  XNOR2_X1 U414 ( .A(n460), .B(n459), .ZN(n711) );
  XNOR2_X1 U415 ( .A(G107), .B(G116), .ZN(n455) );
  XNOR2_X1 U416 ( .A(n446), .B(n445), .ZN(n449) );
  NAND2_X1 U417 ( .A1(n346), .A2(n350), .ZN(n362) );
  NAND2_X1 U418 ( .A1(n632), .A2(n349), .ZN(n361) );
  NAND2_X1 U419 ( .A1(n704), .A2(G210), .ZN(n617) );
  AND2_X1 U420 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U421 ( .A(n569), .B(KEYINPUT36), .ZN(n572) );
  XNOR2_X1 U422 ( .A(n360), .B(n494), .ZN(n530) );
  NOR2_X1 U423 ( .A1(n491), .A2(n492), .ZN(n360) );
  INV_X1 U424 ( .A(KEYINPUT102), .ZN(n473) );
  XOR2_X1 U425 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n347) );
  OR2_X1 U426 ( .A1(n498), .A2(n497), .ZN(n348) );
  AND2_X1 U427 ( .A1(n418), .A2(n593), .ZN(n349) );
  AND2_X1 U428 ( .A1(n418), .A2(n348), .ZN(n350) );
  NAND2_X1 U429 ( .A1(n358), .A2(n356), .ZN(n509) );
  XNOR2_X2 U430 ( .A(n507), .B(n506), .ZN(n732) );
  OR2_X1 U431 ( .A1(n592), .A2(n633), .ZN(n632) );
  XOR2_X1 U432 ( .A(n454), .B(n453), .Z(n363) );
  XOR2_X1 U433 ( .A(KEYINPUT78), .B(KEYINPUT24), .Z(n364) );
  AND2_X1 U434 ( .A1(G214), .A2(n441), .ZN(n365) );
  AND2_X1 U435 ( .A1(n697), .A2(n482), .ZN(n366) );
  XNOR2_X1 U436 ( .A(n536), .B(n535), .ZN(n592) );
  INV_X1 U437 ( .A(KEYINPUT47), .ZN(n566) );
  XNOR2_X1 U438 ( .A(n567), .B(n566), .ZN(n583) );
  INV_X1 U439 ( .A(n550), .ZN(n480) );
  NOR2_X1 U440 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U441 ( .A(KEYINPUT48), .B(KEYINPUT82), .ZN(n586) );
  XNOR2_X1 U442 ( .A(n442), .B(n365), .ZN(n446) );
  INV_X1 U443 ( .A(G469), .ZN(n378) );
  INV_X1 U444 ( .A(n539), .ZN(n540) );
  XNOR2_X1 U445 ( .A(n458), .B(n457), .ZN(n459) );
  AND2_X1 U446 ( .A1(n541), .A2(n540), .ZN(n542) );
  INV_X1 U447 ( .A(n570), .ZN(n571) );
  AND2_X1 U448 ( .A1(n543), .A2(n542), .ZN(n578) );
  OR2_X1 U449 ( .A1(n723), .A2(G952), .ZN(n611) );
  INV_X1 U450 ( .A(G128), .ZN(n367) );
  INV_X1 U451 ( .A(KEYINPUT69), .ZN(n369) );
  XNOR2_X1 U452 ( .A(n369), .B(KEYINPUT4), .ZN(n413) );
  XNOR2_X1 U453 ( .A(G137), .B(n413), .ZN(n370) );
  INV_X1 U454 ( .A(KEYINPUT64), .ZN(n372) );
  XNOR2_X2 U455 ( .A(n372), .B(G953), .ZN(n723) );
  NAND2_X1 U456 ( .A1(n723), .A2(G227), .ZN(n373) );
  XOR2_X1 U457 ( .A(G140), .B(G131), .Z(n447) );
  XNOR2_X1 U458 ( .A(n374), .B(n447), .ZN(n375) );
  XNOR2_X1 U459 ( .A(n716), .B(n377), .ZN(n705) );
  XNOR2_X2 U460 ( .A(n379), .B(n378), .ZN(n554) );
  XNOR2_X1 U461 ( .A(n554), .B(KEYINPUT1), .ZN(n499) );
  XOR2_X1 U462 ( .A(KEYINPUT5), .B(KEYINPUT94), .Z(n381) );
  XNOR2_X1 U463 ( .A(G146), .B(G131), .ZN(n380) );
  XNOR2_X1 U464 ( .A(n381), .B(n380), .ZN(n383) );
  NOR2_X1 U465 ( .A1(G953), .A2(G237), .ZN(n441) );
  NAND2_X1 U466 ( .A1(n441), .A2(G210), .ZN(n382) );
  XNOR2_X1 U467 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U468 ( .A(n384), .B(n407), .ZN(n385) );
  XNOR2_X1 U469 ( .A(n386), .B(n385), .ZN(n595) );
  INV_X1 U470 ( .A(G902), .ZN(n398) );
  NAND2_X1 U471 ( .A1(n595), .A2(n398), .ZN(n387) );
  XOR2_X1 U472 ( .A(G137), .B(G110), .Z(n389) );
  XNOR2_X1 U473 ( .A(n389), .B(n388), .ZN(n392) );
  XNOR2_X1 U474 ( .A(G140), .B(KEYINPUT23), .ZN(n390) );
  XNOR2_X1 U475 ( .A(n364), .B(n390), .ZN(n391) );
  XNOR2_X1 U476 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U477 ( .A(n410), .B(KEYINPUT10), .ZN(n448) );
  XNOR2_X1 U478 ( .A(n393), .B(n448), .ZN(n397) );
  NAND2_X1 U479 ( .A1(n723), .A2(G234), .ZN(n395) );
  XNOR2_X1 U480 ( .A(KEYINPUT79), .B(KEYINPUT8), .ZN(n394) );
  XNOR2_X1 U481 ( .A(n395), .B(n394), .ZN(n456) );
  AND2_X1 U482 ( .A1(n456), .A2(G221), .ZN(n396) );
  XNOR2_X1 U483 ( .A(n397), .B(n396), .ZN(n609) );
  NAND2_X1 U484 ( .A1(n609), .A2(n398), .ZN(n403) );
  XNOR2_X1 U485 ( .A(KEYINPUT15), .B(G902), .ZN(n594) );
  NAND2_X1 U486 ( .A1(n594), .A2(G234), .ZN(n400) );
  XNOR2_X1 U487 ( .A(KEYINPUT20), .B(KEYINPUT92), .ZN(n399) );
  XNOR2_X1 U488 ( .A(n400), .B(n399), .ZN(n464) );
  NAND2_X1 U489 ( .A1(G217), .A2(n464), .ZN(n401) );
  XNOR2_X1 U490 ( .A(KEYINPUT25), .B(n401), .ZN(n402) );
  OR2_X1 U491 ( .A1(n665), .A2(n480), .ZN(n404) );
  NOR2_X1 U492 ( .A1(n658), .A2(n404), .ZN(n470) );
  XNOR2_X1 U493 ( .A(KEYINPUT16), .B(G122), .ZN(n405) );
  XNOR2_X1 U494 ( .A(n406), .B(n405), .ZN(n408) );
  XNOR2_X1 U495 ( .A(n408), .B(n407), .ZN(n628) );
  XNOR2_X1 U496 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U497 ( .A(n412), .B(n411), .ZN(n416) );
  NAND2_X1 U498 ( .A1(n723), .A2(G224), .ZN(n414) );
  XNOR2_X1 U499 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U500 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U501 ( .A(n628), .B(n417), .ZN(n615) );
  INV_X1 U502 ( .A(n594), .ZN(n418) );
  NOR2_X1 U503 ( .A1(G237), .A2(G902), .ZN(n420) );
  INV_X1 U504 ( .A(KEYINPUT73), .ZN(n419) );
  XNOR2_X1 U505 ( .A(n420), .B(n419), .ZN(n425) );
  INV_X1 U506 ( .A(G210), .ZN(n421) );
  OR2_X1 U507 ( .A1(n425), .A2(n421), .ZN(n422) );
  XNOR2_X2 U508 ( .A(n423), .B(n422), .ZN(n575) );
  INV_X1 U509 ( .A(G214), .ZN(n424) );
  OR2_X1 U510 ( .A1(n425), .A2(n424), .ZN(n643) );
  INV_X1 U511 ( .A(n643), .ZN(n426) );
  INV_X1 U512 ( .A(G953), .ZN(n428) );
  NOR2_X1 U513 ( .A1(G898), .A2(n428), .ZN(n626) );
  NAND2_X1 U514 ( .A1(G237), .A2(G234), .ZN(n429) );
  XNOR2_X1 U515 ( .A(n429), .B(KEYINPUT14), .ZN(n432) );
  NAND2_X1 U516 ( .A1(n432), .A2(G902), .ZN(n430) );
  XOR2_X1 U517 ( .A(KEYINPUT88), .B(n430), .Z(n474) );
  NAND2_X1 U518 ( .A1(n626), .A2(n474), .ZN(n431) );
  XNOR2_X1 U519 ( .A(KEYINPUT89), .B(n431), .ZN(n434) );
  NAND2_X1 U520 ( .A1(n432), .A2(G952), .ZN(n433) );
  XOR2_X1 U521 ( .A(KEYINPUT87), .B(n433), .Z(n675) );
  NOR2_X1 U522 ( .A1(G953), .A2(n675), .ZN(n479) );
  NOR2_X1 U523 ( .A1(n434), .A2(n479), .ZN(n436) );
  INV_X1 U524 ( .A(KEYINPUT90), .ZN(n435) );
  XNOR2_X1 U525 ( .A(n436), .B(n435), .ZN(n437) );
  NAND2_X1 U526 ( .A1(n562), .A2(n437), .ZN(n439) );
  XNOR2_X1 U527 ( .A(KEYINPUT68), .B(KEYINPUT0), .ZN(n438) );
  XNOR2_X1 U528 ( .A(n439), .B(n438), .ZN(n501) );
  XNOR2_X1 U529 ( .A(n347), .B(n440), .ZN(n442) );
  XNOR2_X1 U530 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U531 ( .A(n448), .B(n447), .ZN(n717) );
  XNOR2_X1 U532 ( .A(n449), .B(n717), .ZN(n604) );
  NOR2_X1 U533 ( .A1(n604), .A2(G902), .ZN(n450) );
  INV_X1 U534 ( .A(n515), .ZN(n463) );
  XNOR2_X1 U535 ( .A(G122), .B(KEYINPUT98), .ZN(n452) );
  XNOR2_X1 U536 ( .A(n452), .B(KEYINPUT9), .ZN(n454) );
  XOR2_X1 U537 ( .A(KEYINPUT7), .B(KEYINPUT97), .Z(n453) );
  XNOR2_X1 U538 ( .A(n363), .B(n455), .ZN(n460) );
  NAND2_X1 U539 ( .A1(n456), .A2(G217), .ZN(n458) );
  NOR2_X1 U540 ( .A1(G902), .A2(n711), .ZN(n462) );
  XOR2_X1 U541 ( .A(KEYINPUT99), .B(G478), .Z(n461) );
  NAND2_X1 U542 ( .A1(n463), .A2(n516), .ZN(n646) );
  AND2_X1 U543 ( .A1(n464), .A2(G221), .ZN(n466) );
  INV_X1 U544 ( .A(KEYINPUT21), .ZN(n465) );
  XNOR2_X1 U545 ( .A(n466), .B(n465), .ZN(n654) );
  OR2_X1 U546 ( .A1(n646), .A2(n654), .ZN(n467) );
  OR2_X2 U547 ( .A1(n501), .A2(n467), .ZN(n469) );
  XNOR2_X1 U548 ( .A(KEYINPUT67), .B(KEYINPUT22), .ZN(n468) );
  XNOR2_X2 U549 ( .A(n469), .B(n468), .ZN(n521) );
  NAND2_X1 U550 ( .A1(n470), .A2(n521), .ZN(n472) );
  INV_X1 U551 ( .A(KEYINPUT101), .ZN(n471) );
  XNOR2_X1 U552 ( .A(n528), .B(G110), .ZN(G12) );
  NAND2_X1 U553 ( .A1(n516), .A2(n515), .ZN(n546) );
  XNOR2_X2 U554 ( .A(n546), .B(n473), .ZN(n697) );
  INV_X1 U555 ( .A(n723), .ZN(n475) );
  NAND2_X1 U556 ( .A1(n475), .A2(n474), .ZN(n476) );
  NOR2_X1 U557 ( .A1(G900), .A2(n476), .ZN(n477) );
  XOR2_X1 U558 ( .A(KEYINPUT103), .B(n477), .Z(n478) );
  NOR2_X1 U559 ( .A1(n479), .A2(n478), .ZN(n539) );
  NOR2_X1 U560 ( .A1(n539), .A2(n654), .ZN(n549) );
  NAND2_X1 U561 ( .A1(n549), .A2(n643), .ZN(n481) );
  XNOR2_X1 U562 ( .A(n665), .B(KEYINPUT6), .ZN(n519) );
  INV_X1 U563 ( .A(n519), .ZN(n483) );
  NAND2_X1 U564 ( .A1(n366), .A2(n483), .ZN(n568) );
  OR2_X1 U565 ( .A1(n658), .A2(n568), .ZN(n484) );
  XNOR2_X1 U566 ( .A(n484), .B(KEYINPUT43), .ZN(n485) );
  AND2_X1 U567 ( .A1(n485), .A2(n575), .ZN(n589) );
  XOR2_X1 U568 ( .A(G140), .B(KEYINPUT111), .Z(n486) );
  XOR2_X1 U569 ( .A(n589), .B(n486), .Z(G42) );
  INV_X1 U570 ( .A(KEYINPUT86), .ZN(n487) );
  XNOR2_X1 U571 ( .A(n658), .B(n487), .ZN(n570) );
  INV_X1 U572 ( .A(KEYINPUT100), .ZN(n488) );
  XNOR2_X1 U573 ( .A(n550), .B(n488), .ZN(n656) );
  INV_X1 U574 ( .A(n656), .ZN(n489) );
  NAND2_X1 U575 ( .A1(n519), .A2(n489), .ZN(n490) );
  OR2_X1 U576 ( .A1(n570), .A2(n490), .ZN(n492) );
  INV_X1 U577 ( .A(n521), .ZN(n491) );
  INV_X1 U578 ( .A(KEYINPUT76), .ZN(n493) );
  XNOR2_X1 U579 ( .A(n493), .B(KEYINPUT32), .ZN(n494) );
  XNOR2_X1 U580 ( .A(n530), .B(G119), .ZN(G21) );
  INV_X1 U581 ( .A(KEYINPUT2), .ZN(n495) );
  INV_X1 U582 ( .A(KEYINPUT74), .ZN(n496) );
  NOR2_X1 U583 ( .A1(KEYINPUT2), .A2(n496), .ZN(n498) );
  NOR2_X1 U584 ( .A1(n495), .A2(KEYINPUT74), .ZN(n497) );
  NOR2_X1 U585 ( .A1(n550), .A2(n654), .ZN(n659) );
  NAND2_X1 U586 ( .A1(n659), .A2(n499), .ZN(n510) );
  XNOR2_X1 U587 ( .A(n500), .B(KEYINPUT33), .ZN(n652) );
  NOR2_X1 U588 ( .A1(n652), .A2(n501), .ZN(n503) );
  XOR2_X1 U589 ( .A(KEYINPUT34), .B(KEYINPUT75), .Z(n502) );
  XNOR2_X1 U590 ( .A(n503), .B(n502), .ZN(n505) );
  INV_X1 U591 ( .A(n516), .ZN(n504) );
  AND2_X1 U592 ( .A1(n504), .A2(n515), .ZN(n574) );
  NAND2_X1 U593 ( .A1(n505), .A2(n574), .ZN(n507) );
  INV_X1 U594 ( .A(KEYINPUT35), .ZN(n506) );
  INV_X1 U595 ( .A(KEYINPUT44), .ZN(n527) );
  NAND2_X1 U596 ( .A1(n527), .A2(KEYINPUT84), .ZN(n508) );
  NAND2_X1 U597 ( .A1(n509), .A2(n508), .ZN(n526) );
  INV_X1 U598 ( .A(n665), .ZN(n551) );
  NOR2_X1 U599 ( .A1(n510), .A2(n551), .ZN(n667) );
  INV_X1 U600 ( .A(n501), .ZN(n513) );
  NAND2_X1 U601 ( .A1(n667), .A2(n513), .ZN(n511) );
  XNOR2_X1 U602 ( .A(n511), .B(KEYINPUT31), .ZN(n700) );
  NAND2_X1 U603 ( .A1(n659), .A2(n554), .ZN(n512) );
  XNOR2_X1 U604 ( .A(n512), .B(KEYINPUT93), .ZN(n543) );
  AND2_X1 U605 ( .A1(n543), .A2(n551), .ZN(n514) );
  AND2_X1 U606 ( .A1(n514), .A2(n513), .ZN(n687) );
  OR2_X1 U607 ( .A1(n700), .A2(n687), .ZN(n518) );
  NOR2_X1 U608 ( .A1(n516), .A2(n515), .ZN(n699) );
  INV_X1 U609 ( .A(n699), .ZN(n692) );
  AND2_X1 U610 ( .A1(n546), .A2(n692), .ZN(n648) );
  INV_X1 U611 ( .A(n648), .ZN(n517) );
  NAND2_X1 U612 ( .A1(n518), .A2(n517), .ZN(n524) );
  NAND2_X1 U613 ( .A1(n519), .A2(n656), .ZN(n520) );
  NOR2_X1 U614 ( .A1(n658), .A2(n520), .ZN(n522) );
  AND2_X1 U615 ( .A1(n522), .A2(n521), .ZN(n685) );
  INV_X1 U616 ( .A(n685), .ZN(n523) );
  AND2_X1 U617 ( .A1(n524), .A2(n523), .ZN(n525) );
  AND2_X1 U618 ( .A1(n528), .A2(n527), .ZN(n529) );
  NAND2_X1 U619 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U620 ( .A1(n531), .A2(KEYINPUT84), .ZN(n532) );
  NAND2_X1 U621 ( .A1(n732), .A2(n532), .ZN(n533) );
  NAND2_X1 U622 ( .A1(n534), .A2(n533), .ZN(n536) );
  XNOR2_X1 U623 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n535) );
  INV_X1 U624 ( .A(n592), .ZN(n635) );
  XOR2_X1 U625 ( .A(KEYINPUT72), .B(KEYINPUT39), .Z(n545) );
  XOR2_X1 U626 ( .A(KEYINPUT30), .B(KEYINPUT104), .Z(n538) );
  NAND2_X1 U627 ( .A1(n665), .A2(n643), .ZN(n537) );
  XNOR2_X1 U628 ( .A(n538), .B(n537), .ZN(n541) );
  XNOR2_X1 U629 ( .A(n575), .B(KEYINPUT38), .ZN(n644) );
  NAND2_X1 U630 ( .A1(n578), .A2(n644), .ZN(n544) );
  XNOR2_X1 U631 ( .A(n545), .B(n544), .ZN(n588) );
  NOR2_X1 U632 ( .A1(n588), .A2(n546), .ZN(n548) );
  INV_X1 U633 ( .A(KEYINPUT40), .ZN(n547) );
  XNOR2_X1 U634 ( .A(n548), .B(n547), .ZN(n729) );
  NAND2_X1 U635 ( .A1(n550), .A2(n549), .ZN(n552) );
  XNOR2_X1 U636 ( .A(n553), .B(KEYINPUT28), .ZN(n555) );
  NAND2_X1 U637 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U638 ( .A(n556), .B(KEYINPUT106), .ZN(n564) );
  NAND2_X1 U639 ( .A1(n644), .A2(n643), .ZN(n647) );
  NOR2_X1 U640 ( .A1(n647), .A2(n646), .ZN(n558) );
  XOR2_X1 U641 ( .A(KEYINPUT41), .B(KEYINPUT107), .Z(n557) );
  XNOR2_X1 U642 ( .A(n558), .B(n557), .ZN(n677) );
  NOR2_X1 U643 ( .A1(n564), .A2(n677), .ZN(n559) );
  XOR2_X1 U644 ( .A(KEYINPUT42), .B(n559), .Z(n730) );
  NAND2_X1 U645 ( .A1(n729), .A2(n730), .ZN(n561) );
  XNOR2_X1 U646 ( .A(KEYINPUT46), .B(KEYINPUT83), .ZN(n560) );
  XNOR2_X1 U647 ( .A(n561), .B(n560), .ZN(n585) );
  INV_X1 U648 ( .A(n562), .ZN(n563) );
  NOR2_X1 U649 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U650 ( .A(n565), .B(KEYINPUT77), .ZN(n691) );
  NOR2_X1 U651 ( .A1(n691), .A2(n648), .ZN(n567) );
  XNOR2_X1 U652 ( .A(KEYINPUT108), .B(n573), .ZN(n734) );
  INV_X1 U653 ( .A(n734), .ZN(n581) );
  INV_X1 U654 ( .A(n574), .ZN(n576) );
  NOR2_X1 U655 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U656 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U657 ( .A(KEYINPUT105), .B(n579), .ZN(n728) );
  INV_X1 U658 ( .A(n728), .ZN(n580) );
  NAND2_X1 U659 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U660 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U661 ( .A1(n585), .A2(n584), .ZN(n587) );
  NOR2_X1 U662 ( .A1(n588), .A2(n692), .ZN(n702) );
  OR2_X1 U663 ( .A1(n702), .A2(n589), .ZN(n590) );
  NAND2_X1 U664 ( .A1(n722), .A2(KEYINPUT2), .ZN(n633) );
  AND2_X1 U665 ( .A1(KEYINPUT74), .A2(KEYINPUT2), .ZN(n593) );
  NAND2_X1 U666 ( .A1(n704), .A2(G472), .ZN(n597) );
  XNOR2_X1 U667 ( .A(n595), .B(KEYINPUT62), .ZN(n596) );
  XNOR2_X1 U668 ( .A(n597), .B(n596), .ZN(n598) );
  NAND2_X1 U669 ( .A1(n598), .A2(n611), .ZN(n601) );
  XNOR2_X1 U670 ( .A(KEYINPUT109), .B(KEYINPUT63), .ZN(n599) );
  XNOR2_X1 U671 ( .A(n599), .B(KEYINPUT85), .ZN(n600) );
  XNOR2_X1 U672 ( .A(n601), .B(n600), .ZN(G57) );
  NAND2_X1 U673 ( .A1(n704), .A2(G475), .ZN(n606) );
  XNOR2_X1 U674 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n602) );
  XNOR2_X1 U675 ( .A(n602), .B(KEYINPUT59), .ZN(n603) );
  XNOR2_X1 U676 ( .A(n604), .B(n603), .ZN(n605) );
  XNOR2_X1 U677 ( .A(n606), .B(n605), .ZN(n607) );
  INV_X1 U678 ( .A(n611), .ZN(n715) );
  NOR2_X1 U679 ( .A1(n607), .A2(n715), .ZN(n608) );
  XNOR2_X1 U680 ( .A(n608), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U681 ( .A1(n704), .A2(G217), .ZN(n610) );
  XNOR2_X1 U682 ( .A(n610), .B(n609), .ZN(n612) );
  NAND2_X1 U683 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U684 ( .A(n613), .B(KEYINPUT121), .ZN(G66) );
  XOR2_X1 U685 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n614) );
  XNOR2_X1 U686 ( .A(n615), .B(n614), .ZN(n616) );
  XNOR2_X1 U687 ( .A(n617), .B(n616), .ZN(n618) );
  NOR2_X1 U688 ( .A1(n618), .A2(n715), .ZN(n619) );
  XNOR2_X1 U689 ( .A(n619), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X1 U690 ( .A1(n592), .A2(G953), .ZN(n625) );
  NAND2_X1 U691 ( .A1(G224), .A2(G953), .ZN(n620) );
  XNOR2_X1 U692 ( .A(n620), .B(KEYINPUT122), .ZN(n621) );
  XNOR2_X1 U693 ( .A(KEYINPUT61), .B(n621), .ZN(n622) );
  NAND2_X1 U694 ( .A1(n622), .A2(G898), .ZN(n623) );
  XNOR2_X1 U695 ( .A(n623), .B(KEYINPUT123), .ZN(n624) );
  NOR2_X1 U696 ( .A1(n625), .A2(n624), .ZN(n630) );
  INV_X1 U697 ( .A(n626), .ZN(n627) );
  NAND2_X1 U698 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U699 ( .A(n630), .B(n629), .ZN(G69) );
  NOR2_X1 U700 ( .A1(n635), .A2(KEYINPUT2), .ZN(n631) );
  XNOR2_X1 U701 ( .A(n631), .B(KEYINPUT80), .ZN(n641) );
  NAND2_X1 U702 ( .A1(n632), .A2(KEYINPUT74), .ZN(n637) );
  NOR2_X1 U703 ( .A1(n633), .A2(KEYINPUT74), .ZN(n634) );
  NAND2_X1 U704 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U705 ( .A1(n637), .A2(n636), .ZN(n639) );
  OR2_X1 U706 ( .A1(n722), .A2(KEYINPUT2), .ZN(n638) );
  NAND2_X1 U707 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U708 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U709 ( .A(n642), .B(KEYINPUT81), .ZN(n682) );
  NOR2_X1 U710 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U711 ( .A1(n646), .A2(n645), .ZN(n651) );
  NOR2_X1 U712 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U713 ( .A(n649), .B(KEYINPUT114), .ZN(n650) );
  NOR2_X1 U714 ( .A1(n651), .A2(n650), .ZN(n653) );
  NOR2_X1 U715 ( .A1(n653), .A2(n652), .ZN(n672) );
  INV_X1 U716 ( .A(n654), .ZN(n655) );
  NOR2_X1 U717 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U718 ( .A(KEYINPUT49), .B(n657), .ZN(n663) );
  NOR2_X1 U719 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U720 ( .A(KEYINPUT112), .B(n660), .Z(n661) );
  XNOR2_X1 U721 ( .A(KEYINPUT50), .B(n661), .ZN(n662) );
  NAND2_X1 U722 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U723 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U724 ( .A1(n667), .A2(n666), .ZN(n668) );
  XOR2_X1 U725 ( .A(KEYINPUT51), .B(n668), .Z(n669) );
  NOR2_X1 U726 ( .A1(n677), .A2(n669), .ZN(n670) );
  XOR2_X1 U727 ( .A(KEYINPUT113), .B(n670), .Z(n671) );
  XOR2_X1 U728 ( .A(KEYINPUT115), .B(n673), .Z(n674) );
  XNOR2_X1 U729 ( .A(n674), .B(KEYINPUT52), .ZN(n676) );
  NOR2_X1 U730 ( .A1(n676), .A2(n675), .ZN(n680) );
  NOR2_X1 U731 ( .A1(n652), .A2(n677), .ZN(n678) );
  OR2_X1 U732 ( .A1(n678), .A2(G953), .ZN(n679) );
  NAND2_X1 U733 ( .A1(n682), .A2(n681), .ZN(n684) );
  XOR2_X1 U734 ( .A(KEYINPUT116), .B(KEYINPUT53), .Z(n683) );
  XNOR2_X1 U735 ( .A(n684), .B(n683), .ZN(G75) );
  XOR2_X1 U736 ( .A(G101), .B(n685), .Z(G3) );
  NAND2_X1 U737 ( .A1(n697), .A2(n687), .ZN(n686) );
  XNOR2_X1 U738 ( .A(n686), .B(G104), .ZN(G6) );
  XOR2_X1 U739 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n689) );
  NAND2_X1 U740 ( .A1(n687), .A2(n699), .ZN(n688) );
  XNOR2_X1 U741 ( .A(n689), .B(n688), .ZN(n690) );
  XNOR2_X1 U742 ( .A(G107), .B(n690), .ZN(G9) );
  NOR2_X1 U743 ( .A1(n692), .A2(n691), .ZN(n694) );
  XNOR2_X1 U744 ( .A(G128), .B(KEYINPUT29), .ZN(n693) );
  XNOR2_X1 U745 ( .A(n694), .B(n693), .ZN(G30) );
  INV_X1 U746 ( .A(n697), .ZN(n695) );
  NOR2_X1 U747 ( .A1(n695), .A2(n691), .ZN(n696) );
  XOR2_X1 U748 ( .A(G146), .B(n696), .Z(G48) );
  NAND2_X1 U749 ( .A1(n697), .A2(n700), .ZN(n698) );
  XNOR2_X1 U750 ( .A(n698), .B(G113), .ZN(G15) );
  NAND2_X1 U751 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U752 ( .A(n701), .B(G116), .ZN(G18) );
  XOR2_X1 U753 ( .A(G134), .B(n702), .Z(n703) );
  XNOR2_X1 U754 ( .A(KEYINPUT110), .B(n703), .ZN(G36) );
  NAND2_X1 U755 ( .A1(n704), .A2(G469), .ZN(n709) );
  XNOR2_X1 U756 ( .A(KEYINPUT58), .B(KEYINPUT117), .ZN(n707) );
  XNOR2_X1 U757 ( .A(n705), .B(KEYINPUT57), .ZN(n706) );
  XNOR2_X1 U758 ( .A(n707), .B(n706), .ZN(n708) );
  XNOR2_X1 U759 ( .A(n709), .B(n708), .ZN(n710) );
  NOR2_X1 U760 ( .A1(n715), .A2(n710), .ZN(G54) );
  NAND2_X1 U761 ( .A1(n704), .A2(G478), .ZN(n713) );
  XNOR2_X1 U762 ( .A(n711), .B(KEYINPUT120), .ZN(n712) );
  XNOR2_X1 U763 ( .A(n713), .B(n712), .ZN(n714) );
  NOR2_X1 U764 ( .A1(n715), .A2(n714), .ZN(G63) );
  XOR2_X1 U765 ( .A(n716), .B(n717), .Z(n721) );
  XOR2_X1 U766 ( .A(G227), .B(n721), .Z(n718) );
  NAND2_X1 U767 ( .A1(n718), .A2(G900), .ZN(n719) );
  XNOR2_X1 U768 ( .A(n719), .B(KEYINPUT124), .ZN(n720) );
  NAND2_X1 U769 ( .A1(n720), .A2(G953), .ZN(n726) );
  XNOR2_X1 U770 ( .A(n722), .B(n721), .ZN(n724) );
  NAND2_X1 U771 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U772 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U773 ( .A(KEYINPUT125), .B(n727), .Z(G72) );
  XOR2_X1 U774 ( .A(G143), .B(n728), .Z(G45) );
  XNOR2_X1 U775 ( .A(G131), .B(n729), .ZN(G33) );
  XOR2_X1 U776 ( .A(G137), .B(n730), .Z(n731) );
  XNOR2_X1 U777 ( .A(KEYINPUT127), .B(n731), .ZN(G39) );
  XNOR2_X1 U778 ( .A(G122), .B(KEYINPUT126), .ZN(n733) );
  XNOR2_X1 U779 ( .A(n733), .B(n732), .ZN(G24) );
  XNOR2_X1 U780 ( .A(G125), .B(KEYINPUT37), .ZN(n735) );
  XNOR2_X1 U781 ( .A(n735), .B(n734), .ZN(G27) );
endmodule

