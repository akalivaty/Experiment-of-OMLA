//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 0 1 1 0 0 0 1 1 0 0 1 0 1 0 0 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 0 0 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 1 1 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n639, new_n640, new_n641, new_n642, new_n645, new_n646,
    new_n648, new_n649, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT65), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n462), .B1(new_n467), .B2(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n464), .A2(new_n466), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  NOR3_X1   g045(.A1(new_n469), .A2(KEYINPUT65), .A3(new_n470), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n461), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(G101), .A2(G2104), .ZN(new_n474));
  OAI21_X1  g049(.A(KEYINPUT66), .B1(new_n465), .B2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT66), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n476), .A2(new_n463), .A3(KEYINPUT3), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n475), .A2(new_n477), .A3(new_n466), .ZN(new_n478));
  INV_X1    g053(.A(G137), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n474), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AND2_X1   g057(.A1(new_n473), .A2(new_n482), .ZN(G160));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n481), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT69), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n478), .A2(KEYINPUT67), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n475), .A2(new_n477), .A3(new_n488), .A4(new_n466), .ZN(new_n489));
  AOI21_X1  g064(.A(G2105), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n490), .A2(G136), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n481), .B1(new_n487), .B2(new_n489), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT68), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n492), .B(new_n493), .ZN(new_n494));
  AOI211_X1 g069(.A(new_n486), .B(new_n491), .C1(new_n494), .C2(G124), .ZN(G162));
  INV_X1    g070(.A(KEYINPUT70), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n481), .A2(G114), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OR3_X1    g074(.A1(new_n497), .A2(new_n498), .A3(new_n496), .ZN(new_n500));
  AND3_X1   g075(.A1(new_n475), .A2(new_n477), .A3(new_n466), .ZN(new_n501));
  AND2_X1   g076(.A1(G126), .A2(G2105), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n499), .A2(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G138), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n504), .A2(G2105), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n475), .A2(new_n477), .A3(new_n466), .A4(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n507));
  NOR3_X1   g082(.A1(new_n504), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n467), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n503), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(G164));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n513), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G50), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n516), .A2(new_n517), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(KEYINPUT71), .A2(KEYINPUT5), .ZN(new_n522));
  NOR2_X1   g097(.A1(KEYINPUT71), .A2(KEYINPUT5), .ZN(new_n523));
  OAI21_X1  g098(.A(G543), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT5), .ZN(new_n525));
  OAI21_X1  g100(.A(KEYINPUT72), .B1(new_n525), .B2(G543), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT72), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n529), .B(G543), .C1(new_n522), .C2(new_n523), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n521), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G88), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n519), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT71), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(new_n525), .ZN(new_n536));
  NAND2_X1  g111(.A1(KEYINPUT71), .A2(KEYINPUT5), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n513), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n530), .B1(new_n538), .B2(new_n526), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n539), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n515), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n534), .A2(new_n541), .ZN(G166));
  NAND2_X1  g117(.A1(G63), .A2(G651), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n539), .A2(KEYINPUT73), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT73), .ZN(new_n545));
  OAI211_X1 g120(.A(new_n530), .B(new_n545), .C1(new_n538), .C2(new_n526), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n543), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n539), .A2(G89), .A3(new_n520), .ZN(new_n548));
  NAND3_X1  g123(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n549));
  OR2_X1    g124(.A1(KEYINPUT74), .A2(KEYINPUT7), .ZN(new_n550));
  NAND2_X1  g125(.A1(KEYINPUT74), .A2(KEYINPUT7), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n550), .A2(new_n549), .A3(new_n551), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n553), .A2(new_n554), .B1(new_n518), .B2(G51), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n548), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n547), .A2(new_n556), .ZN(G168));
  XOR2_X1   g132(.A(KEYINPUT75), .B(G90), .Z(new_n558));
  NAND3_X1  g133(.A1(new_n539), .A2(new_n520), .A3(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT76), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n518), .A2(G52), .ZN(new_n561));
  AND3_X1   g136(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n560), .B1(new_n559), .B2(new_n561), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n546), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n545), .B1(new_n528), .B2(new_n530), .ZN(new_n566));
  OAI21_X1  g141(.A(G64), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(G77), .A2(G543), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n515), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n564), .A2(new_n569), .ZN(G171));
  OAI21_X1  g145(.A(G56), .B1(new_n565), .B2(new_n566), .ZN(new_n571));
  INV_X1    g146(.A(G68), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(new_n513), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n515), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n531), .A2(G81), .B1(G43), .B2(new_n518), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G860), .ZN(G153));
  NAND4_X1  g154(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g155(.A1(G1), .A2(G3), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT77), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT8), .ZN(new_n583));
  NAND4_X1  g158(.A1(G319), .A2(G483), .A3(G661), .A4(new_n583), .ZN(G188));
  AOI22_X1  g159(.A1(new_n539), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n585), .A2(new_n515), .ZN(new_n586));
  INV_X1    g161(.A(new_n518), .ZN(new_n587));
  INV_X1    g162(.A(G53), .ZN(new_n588));
  OR3_X1    g163(.A1(new_n587), .A2(KEYINPUT9), .A3(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(KEYINPUT9), .B1(new_n587), .B2(new_n588), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n589), .A2(new_n590), .B1(new_n531), .B2(G91), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n586), .A2(new_n591), .ZN(G299));
  INV_X1    g167(.A(G171), .ZN(G301));
  INV_X1    g168(.A(KEYINPUT78), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n594), .B1(new_n547), .B2(new_n556), .ZN(new_n595));
  INV_X1    g170(.A(new_n543), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n596), .B1(new_n565), .B2(new_n566), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n520), .A2(G51), .A3(G543), .ZN(new_n598));
  INV_X1    g173(.A(new_n554), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(new_n552), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n600), .B1(new_n531), .B2(G89), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n597), .A2(new_n601), .A3(KEYINPUT78), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n595), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G286));
  INV_X1    g179(.A(G166), .ZN(G303));
  NAND2_X1  g180(.A1(new_n544), .A2(new_n546), .ZN(new_n606));
  OAI21_X1  g181(.A(G651), .B1(new_n606), .B2(G74), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n531), .A2(G87), .B1(G49), .B2(new_n518), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(G288));
  AOI22_X1  g184(.A1(new_n539), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n610), .A2(new_n515), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT79), .ZN(new_n612));
  INV_X1    g187(.A(G48), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n587), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n518), .A2(KEYINPUT79), .A3(G48), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n531), .A2(G86), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n611), .A2(new_n616), .ZN(G305));
  AOI22_X1  g192(.A1(new_n606), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n618), .A2(new_n515), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n518), .A2(G47), .ZN(new_n620));
  INV_X1    g195(.A(G85), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n532), .B2(new_n621), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(G290));
  NAND2_X1  g199(.A1(new_n539), .A2(G66), .ZN(new_n625));
  INV_X1    g200(.A(G79), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(new_n513), .ZN(new_n627));
  AOI22_X1  g202(.A1(new_n627), .A2(G651), .B1(G54), .B2(new_n518), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n531), .A2(G92), .ZN(new_n629));
  INV_X1    g204(.A(KEYINPUT10), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n531), .A2(KEYINPUT10), .A3(G92), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n628), .A2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(G868), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(new_n635), .B2(G171), .ZN(G284));
  OAI21_X1  g212(.A(new_n636), .B1(new_n635), .B2(G171), .ZN(G321));
  NAND2_X1  g213(.A1(G286), .A2(G868), .ZN(new_n639));
  INV_X1    g214(.A(KEYINPUT80), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g216(.A(KEYINPUT80), .B1(G299), .B2(new_n635), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n641), .B1(new_n639), .B2(new_n642), .ZN(G297));
  AOI21_X1  g218(.A(new_n641), .B1(new_n639), .B2(new_n642), .ZN(G280));
  INV_X1    g219(.A(new_n634), .ZN(new_n645));
  INV_X1    g220(.A(G559), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n645), .B1(new_n646), .B2(G860), .ZN(G148));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(G868), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n649), .B1(G868), .B2(new_n578), .ZN(G323));
  XNOR2_X1  g225(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g226(.A1(new_n481), .A2(G2104), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n469), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT12), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT13), .ZN(new_n655));
  INV_X1    g230(.A(G2100), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT81), .Z(new_n658));
  NAND2_X1  g233(.A1(new_n494), .A2(G123), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n490), .A2(G135), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n481), .A2(G111), .ZN(new_n661));
  OAI21_X1  g236(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n662));
  OAI211_X1 g237(.A(new_n659), .B(new_n660), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(KEYINPUT83), .B(G2096), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n655), .A2(new_n656), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT82), .Z(new_n667));
  NAND3_X1  g242(.A1(new_n658), .A2(new_n665), .A3(new_n667), .ZN(G156));
  XNOR2_X1  g243(.A(G1341), .B(G1348), .ZN(new_n669));
  XOR2_X1   g244(.A(G2443), .B(G2446), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT85), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2451), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2427), .B(G2438), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(G2430), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT15), .B(G2435), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n676), .A2(KEYINPUT14), .A3(new_n677), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n678), .A2(KEYINPUT86), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(KEYINPUT86), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n681), .B1(new_n679), .B2(new_n680), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n672), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n684), .ZN(new_n686));
  INV_X1    g261(.A(new_n672), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n686), .A2(new_n682), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT87), .B(G2454), .ZN(new_n689));
  AND3_X1   g264(.A1(new_n685), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n689), .B1(new_n685), .B2(new_n688), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n669), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(KEYINPUT88), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT88), .ZN(new_n694));
  OAI211_X1 g269(.A(new_n694), .B(new_n669), .C1(new_n690), .C2(new_n691), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NOR3_X1   g271(.A1(new_n690), .A2(new_n691), .A3(new_n669), .ZN(new_n697));
  INV_X1    g272(.A(G14), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n696), .A2(new_n699), .ZN(G401));
  INV_X1    g275(.A(KEYINPUT18), .ZN(new_n701));
  XOR2_X1   g276(.A(G2084), .B(G2090), .Z(new_n702));
  XNOR2_X1  g277(.A(G2067), .B(G2678), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(KEYINPUT17), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n702), .A2(new_n703), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n701), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(new_n656), .ZN(new_n708));
  XOR2_X1   g283(.A(G2072), .B(G2078), .Z(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(new_n704), .B2(KEYINPUT18), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(G2096), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n708), .B(new_n711), .ZN(G227));
  XOR2_X1   g287(.A(KEYINPUT89), .B(KEYINPUT19), .Z(new_n713));
  XNOR2_X1  g288(.A(G1971), .B(G1976), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(G1956), .B(G2474), .ZN(new_n716));
  XNOR2_X1  g291(.A(G1961), .B(G1966), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT20), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n716), .B(new_n717), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n716), .A2(new_n717), .ZN(new_n722));
  MUX2_X1   g297(.A(new_n721), .B(new_n722), .S(new_n715), .Z(new_n723));
  NAND2_X1  g298(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  XOR2_X1   g301(.A(G1991), .B(G1996), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(G1981), .B(G1986), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n728), .A2(new_n729), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n730), .A2(new_n731), .ZN(G229));
  INV_X1    g307(.A(G16), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G6), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n611), .A2(new_n616), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(new_n733), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT92), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT32), .B(G1981), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n736), .A2(KEYINPUT92), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n736), .A2(KEYINPUT92), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n741), .A2(new_n738), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n733), .A2(G23), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G288), .B2(G16), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT33), .B(G1976), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n746), .A2(new_n747), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n733), .A2(KEYINPUT90), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n733), .A2(KEYINPUT90), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(G166), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G22), .B2(new_n752), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n754), .A2(G1971), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n754), .A2(G1971), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n748), .B(new_n749), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n744), .A2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT34), .ZN(new_n759));
  OAI21_X1  g334(.A(KEYINPUT93), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT93), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n761), .B(KEYINPUT34), .C1(new_n744), .C2(new_n757), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(G29), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n764), .A2(G25), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n494), .A2(G119), .ZN(new_n766));
  OAI21_X1  g341(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n767));
  INV_X1    g342(.A(G107), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n767), .B1(new_n768), .B2(G2105), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n490), .B2(G131), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n765), .B1(new_n771), .B2(G29), .ZN(new_n772));
  XOR2_X1   g347(.A(KEYINPUT35), .B(G1991), .Z(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT95), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(KEYINPUT36), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n623), .A2(new_n752), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n752), .A2(G24), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(KEYINPUT91), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT91), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n777), .A2(new_n781), .A3(new_n778), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(G1986), .ZN(new_n784));
  INV_X1    g359(.A(G1986), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n780), .A2(new_n785), .A3(new_n782), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n776), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(new_n759), .B2(new_n758), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT94), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n775), .B1(new_n789), .B2(KEYINPUT36), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n763), .A2(new_n788), .A3(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n791), .B1(new_n763), .B2(new_n788), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT31), .B(G11), .ZN(new_n795));
  INV_X1    g370(.A(G28), .ZN(new_n796));
  AOI21_X1  g371(.A(G29), .B1(new_n796), .B2(KEYINPUT30), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n797), .A2(KEYINPUT103), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(KEYINPUT30), .B2(new_n796), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n797), .A2(KEYINPUT103), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n795), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n733), .A2(G21), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G168), .B2(new_n733), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT102), .B(G1966), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(G2078), .ZN(new_n807));
  NAND2_X1  g382(.A1(G164), .A2(G29), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G27), .B2(G29), .ZN(new_n809));
  AOI211_X1 g384(.A(new_n801), .B(new_n806), .C1(new_n807), .C2(new_n809), .ZN(new_n810));
  OAI221_X1 g385(.A(new_n810), .B1(new_n764), .B2(new_n663), .C1(new_n803), .C2(new_n805), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n645), .A2(G16), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G4), .B2(G16), .ZN(new_n813));
  INV_X1    g388(.A(G1348), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n813), .A2(new_n814), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT24), .ZN(new_n817));
  INV_X1    g392(.A(G34), .ZN(new_n818));
  AOI21_X1  g393(.A(G29), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(new_n817), .B2(new_n818), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G160), .B2(new_n764), .ZN(new_n821));
  OAI22_X1  g396(.A1(new_n821), .A2(G2084), .B1(new_n809), .B2(new_n807), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(G2084), .B2(new_n821), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n815), .A2(new_n816), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n764), .A2(G33), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n490), .A2(G139), .ZN(new_n826));
  NAND2_X1  g401(.A1(G115), .A2(G2104), .ZN(new_n827));
  INV_X1    g402(.A(G127), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n827), .B1(new_n469), .B2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT25), .ZN(new_n830));
  NAND2_X1  g405(.A1(G103), .A2(G2104), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n831), .B2(G2105), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n481), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n833));
  AOI22_X1  g408(.A1(new_n829), .A2(G2105), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n826), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n825), .B1(new_n836), .B2(new_n764), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(G2072), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n750), .A2(G20), .A3(new_n751), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT23), .Z(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(G299), .B2(G16), .ZN(new_n841));
  XOR2_X1   g416(.A(KEYINPUT105), .B(G1956), .Z(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  NOR4_X1   g418(.A1(new_n811), .A2(new_n824), .A3(new_n838), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n764), .A2(G32), .ZN(new_n845));
  NAND3_X1  g420(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT26), .Z(new_n847));
  INV_X1    g422(.A(G105), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n847), .B1(new_n848), .B2(new_n652), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n849), .B1(new_n490), .B2(G141), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n487), .A2(new_n489), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n493), .B1(new_n852), .B2(G2105), .ZN(new_n853));
  AOI211_X1 g428(.A(KEYINPUT68), .B(new_n481), .C1(new_n487), .C2(new_n489), .ZN(new_n854));
  OAI21_X1  g429(.A(G129), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT100), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI211_X1 g432(.A(KEYINPUT100), .B(G129), .C1(new_n853), .C2(new_n854), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n851), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n845), .B1(new_n859), .B2(new_n764), .ZN(new_n860));
  XOR2_X1   g435(.A(KEYINPUT27), .B(G1996), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT101), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n860), .B(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(KEYINPUT98), .B(KEYINPUT28), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n764), .A2(G26), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n494), .A2(G128), .ZN(new_n867));
  OR2_X1    g442(.A1(G104), .A2(G2105), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n868), .B(G2104), .C1(G116), .C2(new_n481), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT97), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n870), .B1(new_n490), .B2(G140), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n867), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n866), .B1(new_n872), .B2(G29), .ZN(new_n873));
  XNOR2_X1  g448(.A(KEYINPUT99), .B(G2067), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n873), .B(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n733), .A2(G5), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(G171), .B2(new_n733), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(G1961), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(G29), .A2(G35), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n880), .B1(G162), .B2(G29), .ZN(new_n881));
  XNOR2_X1  g456(.A(KEYINPUT104), .B(KEYINPUT29), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(G2090), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n881), .B(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n752), .A2(G19), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n885), .B1(new_n578), .B2(new_n752), .ZN(new_n886));
  XNOR2_X1  g461(.A(KEYINPUT96), .B(G1341), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n886), .B(new_n887), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n844), .A2(new_n863), .A3(new_n879), .A4(new_n889), .ZN(new_n890));
  NOR3_X1   g465(.A1(new_n793), .A2(new_n794), .A3(new_n890), .ZN(G311));
  NOR2_X1   g466(.A1(new_n794), .A2(new_n890), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(new_n792), .ZN(G150));
  NAND2_X1  g468(.A1(new_n645), .A2(G559), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT38), .ZN(new_n895));
  OAI21_X1  g470(.A(G67), .B1(new_n565), .B2(new_n566), .ZN(new_n896));
  INV_X1    g471(.A(G80), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n897), .A2(new_n513), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n515), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  AOI22_X1  g475(.A1(new_n531), .A2(G93), .B1(G55), .B2(new_n518), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  OAI22_X1  g477(.A1(new_n575), .A2(new_n577), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(G56), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n904), .B1(new_n544), .B2(new_n546), .ZN(new_n905));
  OAI21_X1  g480(.A(G651), .B1(new_n905), .B2(new_n573), .ZN(new_n906));
  INV_X1    g481(.A(G67), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n907), .B1(new_n544), .B2(new_n546), .ZN(new_n908));
  OAI21_X1  g483(.A(G651), .B1(new_n908), .B2(new_n898), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n906), .A2(new_n909), .A3(new_n576), .A4(new_n901), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n903), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n895), .B(new_n911), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n912), .A2(KEYINPUT39), .ZN(new_n913));
  INV_X1    g488(.A(G860), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(KEYINPUT39), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n900), .A2(new_n902), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n917), .A2(new_n914), .ZN(new_n918));
  XNOR2_X1  g493(.A(KEYINPUT106), .B(KEYINPUT37), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n918), .B(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n916), .A2(new_n920), .ZN(G145));
  INV_X1    g496(.A(KEYINPUT40), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n494), .A2(G130), .ZN(new_n923));
  OAI21_X1  g498(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n924), .A2(KEYINPUT109), .ZN(new_n925));
  INV_X1    g500(.A(G118), .ZN(new_n926));
  AOI22_X1  g501(.A1(new_n924), .A2(KEYINPUT109), .B1(new_n926), .B2(G2105), .ZN(new_n927));
  AOI22_X1  g502(.A1(new_n490), .A2(G142), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n923), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n929), .B(new_n654), .ZN(new_n930));
  INV_X1    g505(.A(new_n771), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n930), .B(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n857), .A2(new_n858), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n850), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n511), .A2(KEYINPUT107), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n503), .A2(new_n510), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n936), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n872), .ZN(new_n942));
  INV_X1    g517(.A(new_n940), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n859), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n941), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n859), .A2(new_n943), .ZN(new_n946));
  AOI211_X1 g521(.A(new_n851), .B(new_n940), .C1(new_n857), .C2(new_n858), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n872), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AOI211_X1 g523(.A(new_n934), .B(new_n835), .C1(new_n945), .C2(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n835), .A2(new_n934), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n835), .A2(new_n934), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n945), .A2(new_n948), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n933), .B1(new_n949), .B2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(G162), .B(G160), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n956), .B(new_n663), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n945), .A2(new_n948), .A3(new_n952), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n950), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n959), .A2(new_n932), .A3(new_n953), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n955), .A2(new_n957), .A3(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(G37), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n957), .B1(new_n955), .B2(new_n960), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n922), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n955), .A2(new_n960), .ZN(new_n966));
  INV_X1    g541(.A(new_n957), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n968), .A2(KEYINPUT40), .A3(new_n962), .A4(new_n961), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n965), .A2(new_n969), .ZN(G395));
  OAI21_X1  g545(.A(KEYINPUT112), .B1(new_n917), .B2(G868), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n903), .A2(new_n910), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n972), .B(new_n648), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n634), .A2(G299), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT41), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n628), .A2(new_n633), .A3(new_n586), .A4(new_n591), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n974), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  XOR2_X1   g552(.A(KEYINPUT111), .B(KEYINPUT41), .Z(new_n978));
  AOI21_X1  g553(.A(new_n978), .B1(new_n974), .B2(new_n976), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  OR2_X1    g555(.A1(new_n973), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n974), .A2(new_n976), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n982), .B(KEYINPUT110), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n973), .ZN(new_n984));
  NAND2_X1  g559(.A1(G290), .A2(new_n735), .ZN(new_n985));
  INV_X1    g560(.A(G288), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n986), .A2(G303), .ZN(new_n987));
  NOR2_X1   g562(.A1(G288), .A2(G166), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NOR3_X1   g564(.A1(new_n735), .A2(new_n619), .A3(new_n622), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n985), .A2(new_n989), .A3(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n623), .A2(G305), .ZN(new_n993));
  OAI22_X1  g568(.A1(new_n993), .A2(new_n990), .B1(new_n987), .B2(new_n988), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n992), .A2(new_n994), .A3(KEYINPUT42), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT42), .B1(new_n992), .B2(new_n994), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n981), .B(new_n984), .C1(new_n995), .C2(new_n996), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n997), .A2(G868), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n981), .A2(new_n984), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n995), .A2(new_n996), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n971), .B1(new_n998), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT112), .ZN(new_n1003));
  AND4_X1   g578(.A1(new_n1003), .A2(new_n1001), .A3(G868), .A4(new_n997), .ZN(new_n1004));
  OAI21_X1  g579(.A(KEYINPUT113), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n998), .A2(new_n1003), .A3(new_n1001), .ZN(new_n1006));
  INV_X1    g581(.A(new_n971), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1001), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n997), .A2(G868), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1007), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1006), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1005), .A2(new_n1012), .ZN(G295));
  NOR2_X1   g588(.A1(new_n1002), .A2(new_n1004), .ZN(G331));
  NAND2_X1  g589(.A1(new_n992), .A2(new_n994), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n1017));
  OAI21_X1  g592(.A(G168), .B1(new_n564), .B2(new_n569), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n559), .A2(new_n561), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT76), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G64), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1023), .B1(new_n544), .B2(new_n546), .ZN(new_n1024));
  INV_X1    g599(.A(new_n568), .ZN(new_n1025));
  OAI21_X1  g600(.A(G651), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1022), .A2(new_n595), .A3(new_n1026), .A4(new_n602), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT115), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1018), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(G286), .A2(G171), .A3(KEYINPUT115), .ZN(new_n1030));
  AOI221_X4 g605(.A(new_n1017), .B1(new_n903), .B2(new_n910), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT116), .B1(new_n1032), .B2(new_n972), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n911), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1035));
  INV_X1    g610(.A(new_n982), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n978), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n982), .A2(KEYINPUT41), .ZN(new_n1038));
  AOI22_X1  g613(.A1(new_n1034), .A2(new_n1035), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1032), .A2(new_n972), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n983), .A2(new_n1040), .A3(new_n1035), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1016), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n980), .B1(new_n1040), .B2(new_n1035), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1044), .B1(new_n1034), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(G37), .B1(new_n1046), .B2(new_n1015), .ZN(new_n1047));
  XNOR2_X1  g622(.A(KEYINPUT114), .B(KEYINPUT43), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1043), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1048), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1040), .A2(new_n1017), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1032), .A2(KEYINPUT116), .A3(new_n972), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1045), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1040), .A2(new_n1035), .ZN(new_n1054));
  INV_X1    g629(.A(new_n980), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1053), .A2(new_n1015), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(new_n962), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1015), .B1(new_n1053), .B2(new_n1056), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1050), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT44), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1049), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1051), .A2(new_n1035), .A3(new_n1052), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1015), .B1(new_n1065), .B2(new_n1041), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT43), .B1(new_n1066), .B2(new_n1058), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1059), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1047), .A2(new_n1068), .A3(new_n1048), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1061), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1062), .A2(new_n1070), .ZN(G397));
  INV_X1    g646(.A(G8), .ZN(new_n1072));
  NOR2_X1   g647(.A1(G166), .A2(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n1073), .B(KEYINPUT55), .ZN(new_n1074));
  INV_X1    g649(.A(G1384), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n500), .A2(new_n499), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n501), .A2(new_n502), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  AOI22_X1  g653(.A1(new_n506), .A2(KEYINPUT4), .B1(new_n467), .B2(new_n508), .ZN(new_n1079));
  OAI211_X1 g654(.A(KEYINPUT45), .B(new_n1075), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT45), .B1(new_n511), .B2(new_n1075), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n467), .A2(new_n462), .A3(G125), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT65), .B1(new_n469), .B2(new_n470), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1084), .A2(new_n1085), .B1(G113), .B2(G2104), .ZN(new_n1086));
  OAI211_X1 g661(.A(G40), .B(new_n482), .C1(new_n1086), .C2(new_n481), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT117), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n473), .A2(KEYINPUT117), .A3(G40), .A4(new_n482), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1083), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT50), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1094), .B(new_n1075), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n511), .A2(KEYINPUT120), .A3(new_n1094), .A4(new_n1075), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n511), .A2(new_n1075), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(KEYINPUT50), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1091), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  OAI22_X1  g677(.A1(new_n1093), .A2(G1971), .B1(new_n1102), .B2(G2090), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1074), .B1(new_n1103), .B2(G8), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1092), .A2(new_n804), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1089), .A2(new_n1090), .B1(KEYINPUT50), .B2(new_n1100), .ZN(new_n1106));
  INV_X1    g681(.A(G2084), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1106), .A2(new_n1107), .A3(new_n1095), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT63), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1109), .A2(new_n1110), .A3(G8), .A4(new_n603), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1074), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1091), .A2(new_n1095), .A3(new_n1101), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1113), .A2(G2090), .ZN(new_n1114));
  AOI21_X1  g689(.A(G1971), .B1(new_n1083), .B2(new_n1091), .ZN(new_n1115));
  OAI21_X1  g690(.A(G8), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  OAI22_X1  g691(.A1(new_n1104), .A2(new_n1111), .B1(new_n1112), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT119), .B1(G305), .B2(G1981), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT119), .ZN(new_n1119));
  INV_X1    g694(.A(G1981), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n611), .A2(new_n616), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(G305), .A2(G1981), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT49), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AOI22_X1  g701(.A1(new_n1118), .A2(new_n1121), .B1(G1981), .B2(G305), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT49), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1100), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1072), .B1(new_n1091), .B2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1126), .A2(new_n1128), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT52), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n986), .A2(G1976), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1132), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1134));
  AND2_X1   g709(.A1(new_n1130), .A2(new_n1133), .ZN(new_n1135));
  INV_X1    g710(.A(G1976), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT52), .B1(G288), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1134), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1117), .A2(new_n1131), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1116), .A2(new_n1112), .ZN(new_n1140));
  AOI211_X1 g715(.A(new_n1072), .B(G286), .C1(new_n1105), .C2(new_n1108), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1140), .A2(new_n1131), .A3(new_n1138), .A4(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(KEYINPUT63), .ZN(new_n1143));
  NOR2_X1   g718(.A1(G288), .A2(G1976), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1128), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1130), .B1(new_n1127), .B2(KEYINPUT49), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1144), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(new_n1122), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(new_n1130), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1139), .A2(new_n1143), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(G168), .ZN(new_n1151));
  OAI21_X1  g726(.A(G8), .B1(new_n1109), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT123), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1152), .A2(new_n1153), .A3(KEYINPUT51), .ZN(new_n1154));
  XNOR2_X1  g729(.A(KEYINPUT123), .B(KEYINPUT51), .ZN(new_n1155));
  OAI211_X1 g730(.A(G8), .B(new_n1155), .C1(new_n1109), .C2(new_n1151), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1109), .A2(G8), .A3(new_n1151), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1154), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(KEYINPUT62), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT62), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1154), .A2(new_n1160), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1131), .A2(new_n1138), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1116), .A2(new_n1112), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n1162), .A2(new_n1104), .A3(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT53), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1165), .B1(new_n1092), .B2(G2078), .ZN(new_n1166));
  INV_X1    g741(.A(G1961), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1113), .A2(new_n1167), .ZN(new_n1168));
  AND2_X1   g743(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1093), .A2(KEYINPUT53), .A3(new_n807), .ZN(new_n1170));
  AOI21_X1  g745(.A(G301), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1159), .A2(new_n1161), .A3(new_n1164), .A4(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g747(.A(G299), .B(KEYINPUT57), .ZN(new_n1173));
  AOI21_X1  g748(.A(G1956), .B1(new_n1106), .B2(new_n1099), .ZN(new_n1174));
  XNOR2_X1  g749(.A(KEYINPUT56), .B(G2072), .ZN(new_n1175));
  AND3_X1   g750(.A1(new_n1083), .A2(new_n1091), .A3(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1173), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT121), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(G1348), .B1(new_n1106), .B2(new_n1095), .ZN(new_n1180));
  INV_X1    g755(.A(G2067), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1091), .A2(new_n1181), .A3(new_n1129), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1182), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n645), .B1(new_n1180), .B2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g759(.A(KEYINPUT121), .B(new_n1173), .C1(new_n1174), .C2(new_n1176), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1179), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(G1956), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1102), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT57), .ZN(new_n1189));
  XNOR2_X1  g764(.A(G299), .B(new_n1189), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1083), .A2(new_n1091), .A3(new_n1175), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1188), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  AND2_X1   g767(.A1(new_n1186), .A2(new_n1192), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1179), .A2(KEYINPUT61), .A3(new_n1185), .A4(new_n1192), .ZN(new_n1194));
  INV_X1    g769(.A(G1996), .ZN(new_n1195));
  AND3_X1   g770(.A1(new_n1083), .A2(new_n1091), .A3(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g771(.A(KEYINPUT58), .B(G1341), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1197), .B1(new_n1091), .B2(new_n1129), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n578), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1199), .A2(KEYINPUT59), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT59), .ZN(new_n1201));
  OAI211_X1 g776(.A(new_n1201), .B(new_n578), .C1(new_n1196), .C2(new_n1198), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1180), .A2(new_n1183), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n634), .A2(KEYINPUT60), .ZN(new_n1204));
  AOI22_X1  g779(.A1(new_n1200), .A2(new_n1202), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g780(.A(new_n1180), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n634), .B1(new_n1206), .B2(new_n1182), .ZN(new_n1207));
  NOR3_X1   g782(.A1(new_n1180), .A2(new_n1183), .A3(new_n645), .ZN(new_n1208));
  OAI21_X1  g783(.A(KEYINPUT60), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  AND3_X1   g784(.A1(new_n1194), .A2(new_n1205), .A3(new_n1209), .ZN(new_n1210));
  AOI21_X1  g785(.A(KEYINPUT61), .B1(new_n1177), .B2(new_n1192), .ZN(new_n1211));
  XNOR2_X1  g786(.A(new_n1211), .B(KEYINPUT122), .ZN(new_n1212));
  AOI21_X1  g787(.A(new_n1193), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n1169), .A2(G301), .A3(new_n1170), .ZN(new_n1214));
  OR2_X1    g789(.A1(new_n1086), .A2(KEYINPUT125), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1086), .A2(KEYINPUT125), .ZN(new_n1216));
  NAND3_X1  g791(.A1(new_n1215), .A2(new_n1216), .A3(G2105), .ZN(new_n1217));
  AND4_X1   g792(.A1(KEYINPUT53), .A2(new_n482), .A3(G40), .A4(new_n807), .ZN(new_n1218));
  NAND3_X1  g793(.A1(new_n1083), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  AND2_X1   g794(.A1(new_n1169), .A2(new_n1219), .ZN(new_n1220));
  OAI211_X1 g795(.A(KEYINPUT54), .B(new_n1214), .C1(new_n1220), .C2(G301), .ZN(new_n1221));
  XNOR2_X1  g796(.A(KEYINPUT124), .B(KEYINPUT54), .ZN(new_n1222));
  AND4_X1   g797(.A1(G301), .A2(new_n1166), .A3(new_n1168), .A4(new_n1219), .ZN(new_n1223));
  OAI21_X1  g798(.A(new_n1222), .B1(new_n1171), .B2(new_n1223), .ZN(new_n1224));
  NAND4_X1  g799(.A1(new_n1164), .A2(new_n1221), .A3(new_n1158), .A4(new_n1224), .ZN(new_n1225));
  OAI211_X1 g800(.A(new_n1150), .B(new_n1172), .C1(new_n1213), .C2(new_n1225), .ZN(new_n1226));
  AND2_X1   g801(.A1(new_n1091), .A2(new_n1082), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n623), .A2(new_n785), .ZN(new_n1228));
  XOR2_X1   g803(.A(new_n1228), .B(KEYINPUT118), .Z(new_n1229));
  INV_X1    g804(.A(new_n1229), .ZN(new_n1230));
  OAI21_X1  g805(.A(new_n1230), .B1(new_n785), .B2(new_n623), .ZN(new_n1231));
  XNOR2_X1  g806(.A(new_n859), .B(G1996), .ZN(new_n1232));
  XNOR2_X1  g807(.A(new_n872), .B(new_n1181), .ZN(new_n1233));
  OR2_X1    g808(.A1(new_n931), .A2(new_n773), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n931), .A2(new_n773), .ZN(new_n1235));
  NAND4_X1  g810(.A1(new_n1232), .A2(new_n1233), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  OAI21_X1  g811(.A(new_n1227), .B1(new_n1231), .B2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g812(.A1(new_n1226), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g813(.A1(new_n1227), .A2(new_n1195), .ZN(new_n1239));
  XNOR2_X1  g814(.A(new_n1239), .B(KEYINPUT46), .ZN(new_n1240));
  INV_X1    g815(.A(new_n1227), .ZN(new_n1241));
  AND2_X1   g816(.A1(new_n1233), .A2(new_n859), .ZN(new_n1242));
  OAI21_X1  g817(.A(new_n1240), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  XNOR2_X1  g818(.A(new_n1243), .B(KEYINPUT47), .ZN(new_n1244));
  NAND2_X1  g819(.A1(new_n1229), .A2(new_n1227), .ZN(new_n1245));
  INV_X1    g820(.A(KEYINPUT48), .ZN(new_n1246));
  XNOR2_X1  g821(.A(new_n1245), .B(new_n1246), .ZN(new_n1247));
  AND2_X1   g822(.A1(new_n1236), .A2(new_n1227), .ZN(new_n1248));
  OAI21_X1  g823(.A(new_n1244), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g824(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1250));
  NAND2_X1  g825(.A1(new_n1250), .A2(new_n1227), .ZN(new_n1251));
  XNOR2_X1  g826(.A(new_n1235), .B(KEYINPUT126), .ZN(new_n1252));
  AOI22_X1  g827(.A1(new_n1251), .A2(new_n1252), .B1(new_n1181), .B2(new_n942), .ZN(new_n1253));
  OR2_X1    g828(.A1(new_n1253), .A2(KEYINPUT127), .ZN(new_n1254));
  AOI21_X1  g829(.A(new_n1241), .B1(new_n1253), .B2(KEYINPUT127), .ZN(new_n1255));
  AOI21_X1  g830(.A(new_n1249), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g831(.A1(new_n1238), .A2(new_n1256), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g832(.A1(new_n1066), .A2(new_n1058), .A3(new_n1050), .ZN(new_n1259));
  AOI21_X1  g833(.A(new_n1048), .B1(new_n1047), .B2(new_n1068), .ZN(new_n1260));
  NOR2_X1   g834(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NOR2_X1   g835(.A1(G227), .A2(new_n459), .ZN(new_n1262));
  OAI21_X1  g836(.A(new_n1262), .B1(new_n730), .B2(new_n731), .ZN(new_n1263));
  AOI21_X1  g837(.A(new_n1263), .B1(new_n696), .B2(new_n699), .ZN(new_n1264));
  OAI21_X1  g838(.A(new_n1264), .B1(new_n963), .B2(new_n964), .ZN(new_n1265));
  NOR2_X1   g839(.A1(new_n1261), .A2(new_n1265), .ZN(G308));
  OAI221_X1 g840(.A(new_n1264), .B1(new_n963), .B2(new_n964), .C1(new_n1259), .C2(new_n1260), .ZN(G225));
endmodule


