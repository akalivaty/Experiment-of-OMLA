//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 0 0 0 0 1 0 1 1 0 0 1 1 0 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 0 0 0 0 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n559, new_n561, new_n562, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n581,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n620, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1193, new_n1195, new_n1196, new_n1197;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT66), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n465), .A2(G137), .ZN(new_n469));
  NAND2_X1  g044(.A1(G101), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n468), .A2(new_n471), .ZN(G160));
  INV_X1    g047(.A(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(KEYINPUT3), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(new_n464), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n477), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  NAND4_X1  g060(.A1(new_n474), .A2(new_n476), .A3(G126), .A4(G2105), .ZN(new_n486));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n487), .A2(new_n489), .A3(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT67), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n474), .A2(new_n476), .A3(G138), .A4(new_n464), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n465), .A2(KEYINPUT4), .A3(G138), .A4(new_n464), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT67), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n486), .A2(new_n497), .A3(new_n490), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n492), .A2(new_n495), .A3(new_n496), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT68), .ZN(new_n500));
  AND2_X1   g075(.A1(new_n495), .A2(new_n496), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT68), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n501), .A2(new_n502), .A3(new_n492), .A4(new_n498), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n506), .A2(KEYINPUT6), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT69), .B(G651), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(KEYINPUT6), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G50), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n508), .A2(KEYINPUT6), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT70), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g090(.A1(KEYINPUT70), .A2(KEYINPUT5), .A3(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n507), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n512), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n510), .A2(new_n511), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n522), .A2(new_n508), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n521), .A2(new_n523), .ZN(G166));
  AND2_X1   g099(.A1(new_n509), .A2(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G51), .ZN(new_n526));
  INV_X1    g101(.A(new_n519), .ZN(new_n527));
  XOR2_X1   g102(.A(KEYINPUT72), .B(G89), .Z(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT7), .ZN(new_n530));
  NAND2_X1  g105(.A1(G76), .A2(G543), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n531), .B2(new_n506), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n526), .A2(new_n529), .A3(new_n532), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n517), .B(KEYINPUT71), .ZN(new_n534));
  INV_X1    g109(.A(G63), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n534), .A2(new_n535), .B1(new_n530), .B2(new_n531), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n533), .B1(G651), .B2(new_n536), .ZN(G168));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G64), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n534), .B2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n508), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(G52), .ZN(new_n543));
  INV_X1    g118(.A(G90), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n510), .A2(new_n543), .B1(new_n519), .B2(new_n544), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n545), .A2(KEYINPUT73), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n545), .A2(KEYINPUT73), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n542), .B1(new_n546), .B2(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n534), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(new_n541), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n525), .A2(G43), .B1(new_n527), .B2(G81), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT74), .ZN(G153));
  AND3_X1   g133(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G36), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n562), .ZN(G188));
  NAND4_X1  g138(.A1(new_n512), .A2(G91), .A3(new_n517), .A4(new_n518), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT76), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n509), .A2(KEYINPUT76), .A3(G91), .A4(new_n517), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n569), .A2(KEYINPUT75), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n525), .A2(G53), .A3(new_n570), .ZN(new_n571));
  XNOR2_X1  g146(.A(KEYINPUT75), .B(KEYINPUT9), .ZN(new_n572));
  INV_X1    g147(.A(G53), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n510), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(G78), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(new_n517), .ZN(new_n576));
  XOR2_X1   g151(.A(KEYINPUT77), .B(G65), .Z(new_n577));
  OAI21_X1  g152(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G651), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n568), .A2(new_n571), .A3(new_n574), .A4(new_n579), .ZN(G299));
  NAND2_X1  g155(.A1(new_n536), .A2(G651), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n581), .A2(new_n526), .A3(new_n532), .A4(new_n529), .ZN(G286));
  INV_X1    g157(.A(G166), .ZN(G303));
  AOI22_X1  g158(.A1(new_n525), .A2(G49), .B1(new_n527), .B2(G87), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT71), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n517), .B(new_n585), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n586), .B2(G74), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n584), .A2(new_n587), .ZN(G288));
  NAND4_X1  g163(.A1(new_n512), .A2(G86), .A3(new_n517), .A4(new_n518), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT78), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n517), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n525), .A2(G48), .B1(new_n592), .B2(new_n541), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(KEYINPUT79), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT79), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n590), .A2(new_n596), .A3(new_n593), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(G305));
  NAND2_X1  g174(.A1(G72), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G60), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n534), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(new_n541), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n525), .A2(G47), .B1(new_n527), .B2(G85), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n576), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n525), .A2(G54), .B1(new_n609), .B2(G651), .ZN(new_n610));
  INV_X1    g185(.A(G92), .ZN(new_n611));
  OAI21_X1  g186(.A(KEYINPUT10), .B1(new_n519), .B2(new_n611), .ZN(new_n612));
  OR3_X1    g187(.A1(new_n519), .A2(KEYINPUT10), .A3(new_n611), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n610), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n606), .B1(G868), .B2(new_n615), .ZN(G284));
  OAI21_X1  g191(.A(new_n606), .B1(G868), .B2(new_n615), .ZN(G321));
  MUX2_X1   g192(.A(G299), .B(G286), .S(G868), .Z(G280));
  XOR2_X1   g193(.A(G280), .B(KEYINPUT80), .Z(G297));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n615), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n615), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g200(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT12), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  INV_X1    g203(.A(G2100), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n478), .A2(G123), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n480), .A2(G135), .ZN(new_n632));
  NOR2_X1   g207(.A1(G99), .A2(G2105), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(new_n464), .B2(G111), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n631), .B(new_n632), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(G2096), .Z(new_n636));
  NAND2_X1  g211(.A1(new_n630), .A2(new_n636), .ZN(G156));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT81), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2427), .B(G2430), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(KEYINPUT14), .ZN(new_n643));
  XOR2_X1   g218(.A(G2451), .B(G2454), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G1341), .B(G1348), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2443), .B(G2446), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(G14), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT82), .Z(G401));
  XNOR2_X1  g227(.A(G2084), .B(G2090), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT83), .Z(new_n654));
  XOR2_X1   g229(.A(G2067), .B(G2678), .Z(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2072), .B(G2078), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT18), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n657), .B(KEYINPUT17), .Z(new_n660));
  AOI21_X1  g235(.A(new_n660), .B1(new_n654), .B2(new_n655), .ZN(new_n661));
  INV_X1    g236(.A(new_n655), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n662), .A2(new_n657), .ZN(new_n663));
  AOI211_X1 g238(.A(new_n656), .B(new_n661), .C1(new_n654), .C2(new_n663), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n659), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2096), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(new_n629), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(G227));
  XNOR2_X1  g243(.A(G1971), .B(G1976), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  XOR2_X1   g245(.A(G1956), .B(G2474), .Z(new_n671));
  XOR2_X1   g246(.A(G1961), .B(G1966), .Z(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT20), .Z(new_n675));
  NOR2_X1   g250(.A1(new_n671), .A2(new_n672), .ZN(new_n676));
  INV_X1    g251(.A(new_n673), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n676), .B1(new_n670), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n670), .A2(KEYINPUT84), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n675), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(G1986), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G1991), .B(G1996), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT22), .B(G1981), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n687), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(G229));
  OAI21_X1  g265(.A(G2104), .B1(new_n464), .B2(G107), .ZN(new_n691));
  INV_X1    g266(.A(G95), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n691), .B1(new_n692), .B2(new_n464), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT85), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n693), .A2(new_n694), .ZN(new_n696));
  AOI22_X1  g271(.A1(new_n695), .A2(new_n696), .B1(G131), .B2(new_n480), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n478), .A2(G119), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  MUX2_X1   g274(.A(G25), .B(new_n699), .S(G29), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT86), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT35), .B(G1991), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n701), .B(new_n702), .Z(new_n703));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G24), .ZN(new_n705));
  INV_X1    g280(.A(G290), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(new_n704), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G1986), .ZN(new_n708));
  AND2_X1   g283(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n709));
  NOR3_X1   g284(.A1(new_n703), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n704), .A2(G22), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G166), .B2(new_n704), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n712), .A2(G1971), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n712), .A2(G1971), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n704), .A2(G23), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G288), .B2(G16), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT87), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n717), .A2(new_n718), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT33), .B(G1976), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  NOR3_X1   g298(.A1(new_n720), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n721), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n722), .B1(new_n725), .B2(new_n719), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n714), .B(new_n715), .C1(new_n724), .C2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n598), .A2(G16), .ZN(new_n728));
  OR2_X1    g303(.A1(G6), .A2(G16), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(KEYINPUT32), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT32), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n728), .A2(new_n732), .A3(new_n729), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G1981), .ZN(new_n735));
  INV_X1    g310(.A(G1981), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n731), .A2(new_n736), .A3(new_n733), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n727), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n738), .A2(KEYINPUT34), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT34), .ZN(new_n740));
  AOI211_X1 g315(.A(new_n740), .B(new_n727), .C1(new_n735), .C2(new_n737), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n710), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI221_X1 g319(.A(new_n710), .B1(KEYINPUT88), .B2(KEYINPUT36), .C1(new_n739), .C2(new_n741), .ZN(new_n745));
  AOI22_X1  g320(.A1(G129), .A2(new_n478), .B1(new_n480), .B2(G141), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n464), .A2(G105), .A3(G2104), .ZN(new_n747));
  NAND3_X1  g322(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT26), .Z(new_n749));
  NAND3_X1  g324(.A1(new_n746), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  MUX2_X1   g325(.A(G32), .B(new_n750), .S(G29), .Z(new_n751));
  XOR2_X1   g326(.A(KEYINPUT27), .B(G1996), .Z(new_n752));
  NOR2_X1   g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  OR2_X1    g328(.A1(KEYINPUT24), .A2(G34), .ZN(new_n754));
  INV_X1    g329(.A(G29), .ZN(new_n755));
  NAND2_X1  g330(.A1(KEYINPUT24), .A2(G34), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G160), .B2(new_n755), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G2084), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n753), .A2(new_n759), .ZN(new_n760));
  OR2_X1    g335(.A1(G29), .A2(G33), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT89), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT25), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(G115), .A2(G2104), .ZN(new_n766));
  INV_X1    g341(.A(G127), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n766), .B1(new_n477), .B2(new_n767), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n768), .A2(G2105), .B1(new_n480), .B2(G139), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n763), .A2(new_n764), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n765), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n761), .B1(new_n771), .B2(new_n755), .ZN(new_n772));
  INV_X1    g347(.A(G2072), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT30), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n775), .A2(G28), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(G28), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n774), .B1(new_n755), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n751), .A2(new_n752), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n635), .A2(new_n755), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n760), .A2(new_n779), .A3(new_n780), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n772), .A2(new_n773), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT90), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT31), .B(G11), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n755), .A2(G27), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G164), .B2(new_n755), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n786), .B1(new_n788), .B2(G2078), .ZN(new_n789));
  NOR3_X1   g364(.A1(new_n783), .A2(new_n785), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n704), .A2(G21), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G168), .B2(new_n704), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT91), .B(G1966), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G5), .A2(G16), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G171), .B2(G16), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n796), .A2(G1961), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n788), .A2(G2078), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n790), .A2(new_n794), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n796), .A2(G1961), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT92), .ZN(new_n801));
  OR3_X1    g376(.A1(new_n799), .A2(KEYINPUT93), .A3(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(KEYINPUT93), .B1(new_n799), .B2(new_n801), .ZN(new_n803));
  NAND2_X1  g378(.A1(G299), .A2(G16), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n704), .A2(KEYINPUT23), .A3(G20), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT23), .ZN(new_n806));
  INV_X1    g381(.A(G20), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n806), .B1(new_n807), .B2(G16), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n804), .A2(new_n805), .A3(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(G1956), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n704), .A2(G19), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(new_n556), .B2(new_n704), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(G1341), .Z(new_n814));
  AND4_X1   g389(.A1(new_n802), .A2(new_n803), .A3(new_n811), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n755), .A2(G35), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G162), .B2(new_n755), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT29), .ZN(new_n818));
  INV_X1    g393(.A(G2090), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n744), .A2(new_n745), .A3(new_n815), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n755), .A2(G26), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n478), .A2(G128), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n480), .A2(G140), .ZN(new_n824));
  OR2_X1    g399(.A1(G104), .A2(G2105), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n825), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n823), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n822), .B1(new_n828), .B2(new_n755), .ZN(new_n829));
  MUX2_X1   g404(.A(new_n822), .B(new_n829), .S(KEYINPUT28), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(G2067), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n704), .A2(G4), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n615), .B2(new_n704), .ZN(new_n833));
  INV_X1    g408(.A(G1348), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  NOR3_X1   g411(.A1(new_n821), .A2(new_n831), .A3(new_n836), .ZN(G311));
  AND3_X1   g412(.A1(new_n744), .A2(new_n745), .A3(new_n815), .ZN(new_n838));
  INV_X1    g413(.A(new_n831), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n838), .A2(new_n839), .A3(new_n835), .A4(new_n820), .ZN(G150));
  NAND2_X1  g415(.A1(G80), .A2(G543), .ZN(new_n841));
  INV_X1    g416(.A(G67), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n841), .B1(new_n534), .B2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT94), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI211_X1 g420(.A(KEYINPUT94), .B(new_n841), .C1(new_n534), .C2(new_n842), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n845), .A2(new_n541), .A3(new_n846), .ZN(new_n847));
  AOI22_X1  g422(.A1(new_n525), .A2(G55), .B1(new_n527), .B2(G93), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XOR2_X1   g424(.A(KEYINPUT96), .B(G860), .Z(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT37), .Z(new_n852));
  NAND2_X1  g427(.A1(new_n615), .A2(G559), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT38), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT39), .Z(new_n855));
  INV_X1    g430(.A(KEYINPUT95), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n553), .A2(new_n856), .A3(new_n554), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n555), .A2(KEYINPUT95), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n849), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n556), .A2(new_n847), .A3(new_n856), .A4(new_n848), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n855), .B(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n852), .B1(new_n862), .B2(new_n850), .ZN(G145));
  XOR2_X1   g438(.A(new_n635), .B(G160), .Z(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n484), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n478), .A2(G130), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n480), .A2(G142), .ZN(new_n867));
  NOR2_X1   g442(.A1(G106), .A2(G2105), .ZN(new_n868));
  OAI21_X1  g443(.A(G2104), .B1(new_n464), .B2(G118), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n866), .B(new_n867), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n699), .B(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT98), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n872), .A2(new_n627), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n627), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n495), .A2(new_n496), .A3(new_n486), .A4(new_n490), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n827), .B(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n750), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT97), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n771), .A2(new_n879), .ZN(new_n880));
  AND2_X1   g455(.A1(new_n771), .A2(new_n879), .ZN(new_n881));
  OR3_X1    g456(.A1(new_n878), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT99), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n878), .A2(new_n880), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n865), .B1(new_n875), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n882), .A2(new_n884), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n883), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n886), .B1(new_n875), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(G37), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n873), .A2(KEYINPUT100), .A3(new_n874), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n891), .A2(new_n887), .ZN(new_n892));
  INV_X1    g467(.A(new_n865), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n893), .B1(new_n891), .B2(new_n887), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n890), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n889), .A2(new_n895), .ZN(new_n896));
  XOR2_X1   g471(.A(new_n896), .B(KEYINPUT40), .Z(G395));
  NOR2_X1   g472(.A1(new_n849), .A2(G868), .ZN(new_n898));
  INV_X1    g473(.A(G288), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n899), .A2(G290), .ZN(new_n900));
  AOI21_X1  g475(.A(G288), .B1(new_n603), .B2(new_n604), .ZN(new_n901));
  OAI21_X1  g476(.A(KEYINPUT102), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n706), .A2(G288), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT102), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n899), .A2(G290), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(G166), .B1(new_n595), .B2(new_n597), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n595), .A2(G166), .A3(new_n597), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n902), .A2(new_n906), .A3(new_n908), .A4(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n900), .A2(new_n901), .ZN(new_n911));
  INV_X1    g486(.A(new_n909), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n911), .B(new_n904), .C1(new_n912), .C2(new_n907), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT42), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n914), .B(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT103), .ZN(new_n917));
  XNOR2_X1  g492(.A(G299), .B(new_n614), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n918), .A2(KEYINPUT41), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(KEYINPUT41), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n919), .A2(KEYINPUT101), .A3(new_n920), .ZN(new_n921));
  OR2_X1    g496(.A1(new_n920), .A2(KEYINPUT101), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n861), .B(new_n622), .ZN(new_n924));
  OAI22_X1  g499(.A1(new_n916), .A2(new_n917), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n918), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n925), .B1(new_n926), .B2(new_n924), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n916), .A2(new_n917), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n927), .B(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n898), .B1(new_n929), .B2(G868), .ZN(G295));
  AOI21_X1  g505(.A(new_n898), .B1(new_n929), .B2(G868), .ZN(G331));
  NAND2_X1  g506(.A1(G301), .A2(G168), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n545), .B(KEYINPUT73), .ZN(new_n933));
  NAND3_X1  g508(.A1(G286), .A2(new_n933), .A3(new_n542), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n861), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n932), .A2(new_n934), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n936), .A2(new_n859), .A3(new_n860), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n938), .A2(new_n922), .A3(new_n921), .ZN(new_n939));
  INV_X1    g514(.A(new_n914), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n935), .A2(new_n926), .A3(new_n937), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n942), .A2(new_n890), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n919), .A2(new_n920), .ZN(new_n944));
  INV_X1    g519(.A(new_n937), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n936), .B1(new_n859), .B2(new_n860), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n947), .A2(new_n941), .A3(KEYINPUT105), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT105), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n938), .A2(new_n949), .A3(new_n944), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n948), .A2(new_n914), .A3(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n943), .A2(KEYINPUT43), .A3(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT43), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n942), .A2(new_n890), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n940), .B1(new_n939), .B2(new_n941), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n952), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT44), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT43), .B1(new_n954), .B2(new_n955), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT104), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT104), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n961), .B(KEYINPUT43), .C1(new_n954), .C2(new_n955), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n951), .A2(new_n953), .A3(new_n890), .A4(new_n942), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT106), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT106), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n943), .A2(new_n965), .A3(new_n953), .A4(new_n951), .ZN(new_n966));
  AOI22_X1  g541(.A1(new_n960), .A2(new_n962), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n958), .B1(new_n967), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g543(.A(G1384), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n876), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT45), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n468), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n469), .A2(new_n470), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(new_n464), .ZN(new_n975));
  XNOR2_X1  g550(.A(KEYINPUT107), .B(G40), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n973), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n972), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n827), .B(G2067), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OR2_X1    g556(.A1(new_n981), .A2(KEYINPUT108), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(KEYINPUT108), .ZN(new_n983));
  INV_X1    g558(.A(new_n979), .ZN(new_n984));
  XOR2_X1   g559(.A(new_n750), .B(G1996), .Z(new_n985));
  OAI211_X1 g560(.A(new_n982), .B(new_n983), .C1(new_n984), .C2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n699), .A2(new_n702), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n699), .A2(new_n702), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n979), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  OR2_X1    g566(.A1(G290), .A2(G1986), .ZN(new_n992));
  NAND2_X1  g567(.A1(G290), .A2(G1986), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n984), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT121), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n996), .A2(KEYINPUT61), .ZN(new_n997));
  XNOR2_X1  g572(.A(G299), .B(KEYINPUT57), .ZN(new_n998));
  XNOR2_X1  g573(.A(KEYINPUT56), .B(G2072), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n468), .A2(new_n471), .A3(new_n976), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n876), .A2(KEYINPUT45), .A3(new_n969), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n500), .A2(new_n969), .A3(new_n503), .ZN(new_n1004));
  AOI211_X1 g579(.A(new_n1000), .B(new_n1003), .C1(new_n1004), .C2(new_n971), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n500), .A2(new_n1006), .A3(new_n969), .A4(new_n503), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n978), .B1(new_n970), .B2(KEYINPUT50), .ZN(new_n1008));
  AOI21_X1  g583(.A(G1956), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n998), .B1(new_n1005), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1003), .B1(new_n1004), .B2(new_n971), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n999), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n810), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT57), .ZN(new_n1015));
  XNOR2_X1  g590(.A(G299), .B(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1012), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1010), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n996), .A2(KEYINPUT61), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n997), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1004), .A2(new_n971), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1003), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n978), .A2(new_n970), .ZN(new_n1024));
  XNOR2_X1  g599(.A(KEYINPUT58), .B(G1341), .ZN(new_n1025));
  OAI22_X1  g600(.A1(new_n1023), .A2(G1996), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  AND4_X1   g601(.A1(KEYINPUT120), .A2(new_n1026), .A3(KEYINPUT59), .A4(new_n556), .ZN(new_n1027));
  INV_X1    g602(.A(new_n997), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1028), .B1(new_n1010), .B2(new_n1017), .ZN(new_n1029));
  XNOR2_X1  g604(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1030), .B1(new_n1026), .B2(new_n556), .ZN(new_n1031));
  NOR4_X1   g606(.A1(new_n1020), .A2(new_n1027), .A3(new_n1029), .A4(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1004), .A2(KEYINPUT50), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT109), .B1(new_n970), .B2(KEYINPUT50), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT109), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n876), .A2(new_n1035), .A3(new_n1006), .A4(new_n969), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n978), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1033), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n834), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT119), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1001), .A2(new_n969), .A3(new_n876), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1041), .A2(G2067), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1039), .A2(new_n1040), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT60), .ZN(new_n1045));
  AOI21_X1  g620(.A(G1348), .B1(new_n1033), .B2(new_n1037), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT119), .B1(new_n1046), .B2(new_n1042), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1044), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n1048), .A2(new_n615), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1040), .B1(new_n1039), .B2(new_n1043), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n1046), .A2(KEYINPUT119), .A3(new_n1042), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT60), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT122), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1044), .A2(new_n1047), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1055), .A2(KEYINPUT122), .A3(KEYINPUT60), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1049), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1048), .A2(new_n615), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT122), .B1(new_n1055), .B2(KEYINPUT60), .ZN(new_n1059));
  AOI211_X1 g634(.A(new_n1053), .B(new_n1045), .C1(new_n1044), .C2(new_n1047), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1058), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1032), .A2(new_n1057), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT123), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1010), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1055), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n1017), .A2(new_n615), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1064), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n1062), .A2(new_n1063), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1063), .B1(new_n1062), .B2(new_n1067), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT51), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n972), .B(new_n1001), .C1(new_n1004), .C2(new_n971), .ZN(new_n1071));
  INV_X1    g646(.A(G1966), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1073), .B(G168), .C1(G2084), .C2(new_n1038), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1070), .B1(new_n1074), .B2(G8), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1038), .ZN(new_n1076));
  INV_X1    g651(.A(G2084), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n1076), .A2(new_n1077), .B1(new_n1072), .B2(new_n1071), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT51), .B1(new_n1078), .B2(G168), .ZN(new_n1079));
  INV_X1    g654(.A(G8), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1080), .B1(new_n1078), .B2(G168), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1075), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(G1961), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1038), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n1085));
  OR2_X1    g660(.A1(new_n1085), .A2(G2078), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1084), .B(KEYINPUT124), .C1(new_n1071), .C2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT124), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1071), .A2(new_n1086), .ZN(new_n1089));
  AOI21_X1  g664(.A(G1961), .B1(new_n1033), .B2(new_n1037), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1088), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1085), .B1(new_n1023), .B2(G2078), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1087), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(G171), .ZN(new_n1094));
  NAND2_X1  g669(.A1(G160), .A2(G40), .ZN(new_n1095));
  XOR2_X1   g670(.A(new_n1095), .B(KEYINPUT125), .Z(new_n1096));
  NAND2_X1  g671(.A1(new_n972), .A2(new_n1002), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1096), .A2(new_n1086), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT126), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1090), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1100), .B(new_n1092), .C1(new_n1099), .C2(new_n1098), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1094), .B1(new_n1101), .B2(G171), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1082), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(G303), .A2(G8), .ZN(new_n1105));
  XOR2_X1   g680(.A(new_n1105), .B(KEYINPUT55), .Z(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  OR2_X1    g682(.A1(new_n1011), .A2(G1971), .ZN(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT115), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT115), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n819), .B1(new_n1013), .B2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1108), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1112), .A2(KEYINPUT116), .ZN(new_n1113));
  OAI21_X1  g688(.A(G8), .B1(new_n1112), .B2(KEYINPUT116), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1107), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1108), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1038), .A2(G2090), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1106), .B(G8), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT110), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1076), .A2(new_n819), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1080), .B1(new_n1120), .B2(new_n1108), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT110), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1121), .A2(new_n1122), .A3(new_n1106), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1119), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(G1976), .ZN(new_n1125));
  OAI211_X1 g700(.A(G8), .B(new_n1041), .C1(G288), .C2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(KEYINPUT111), .A2(KEYINPUT52), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1024), .A2(new_n1080), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1127), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1129), .B(new_n1130), .C1(new_n1125), .C2(G288), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT52), .ZN(new_n1132));
  NAND3_X1  g707(.A1(G288), .A2(new_n1132), .A3(new_n1125), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1128), .A2(new_n1131), .A3(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g709(.A(KEYINPUT112), .B(G1981), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n590), .A2(new_n593), .A3(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n509), .A2(G48), .A3(G543), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1137), .B(new_n589), .C1(new_n591), .C2(new_n508), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT113), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1138), .A2(new_n1139), .A3(G1981), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1139), .B1(new_n1138), .B2(G1981), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1136), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT49), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1136), .B(KEYINPUT49), .C1(new_n1140), .C2(new_n1141), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1144), .A2(new_n1129), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1134), .A2(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1147), .B(KEYINPUT117), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1115), .A2(new_n1124), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1103), .B1(new_n1101), .B2(G171), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1150), .B1(G171), .B2(new_n1093), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1104), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n1068), .A2(new_n1069), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT63), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1115), .A2(new_n1124), .A3(new_n1148), .ZN(new_n1155));
  NOR3_X1   g730(.A1(new_n1078), .A2(new_n1080), .A3(G286), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1154), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1147), .A2(KEYINPUT114), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT114), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1134), .A2(new_n1146), .A3(new_n1160), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n1159), .B(new_n1161), .C1(new_n1106), .C2(new_n1121), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT118), .ZN(new_n1163));
  OR2_X1    g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1154), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1164), .A2(new_n1165), .A3(new_n1124), .A4(new_n1156), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1158), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1124), .ZN(new_n1168));
  AND2_X1   g743(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1146), .A2(new_n1125), .A3(new_n899), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(new_n1136), .ZN(new_n1171));
  AOI22_X1  g746(.A1(new_n1168), .A2(new_n1169), .B1(new_n1129), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT62), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1094), .B1(new_n1082), .B2(new_n1173), .ZN(new_n1174));
  OAI211_X1 g749(.A(new_n1149), .B(new_n1174), .C1(new_n1173), .C2(new_n1082), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1167), .A2(new_n1172), .A3(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n995), .B1(new_n1153), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT46), .ZN(new_n1178));
  OR3_X1    g753(.A1(new_n984), .A2(new_n1178), .A3(G1996), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n979), .B1(new_n980), .B2(new_n750), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1178), .B1(new_n984), .B2(G1996), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  XOR2_X1   g757(.A(new_n1182), .B(KEYINPUT47), .Z(new_n1183));
  NOR2_X1   g758(.A1(new_n992), .A2(new_n984), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n1184), .B(KEYINPUT127), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n1185), .B(KEYINPUT48), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1186), .A2(new_n991), .ZN(new_n1187));
  INV_X1    g762(.A(new_n989), .ZN(new_n1188));
  OAI22_X1  g763(.A1(new_n986), .A2(new_n1188), .B1(G2067), .B2(new_n827), .ZN(new_n1189));
  AOI211_X1 g764(.A(new_n1183), .B(new_n1187), .C1(new_n979), .C2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1177), .A2(new_n1190), .ZN(G329));
  assign    G231 = 1'b0;
  NAND4_X1  g766(.A1(new_n651), .A2(new_n688), .A3(new_n667), .A4(new_n689), .ZN(new_n1193));
  NOR4_X1   g767(.A1(new_n967), .A2(new_n462), .A3(new_n896), .A4(new_n1193), .ZN(G308));
  INV_X1    g768(.A(new_n967), .ZN(new_n1195));
  INV_X1    g769(.A(new_n896), .ZN(new_n1196));
  INV_X1    g770(.A(new_n1193), .ZN(new_n1197));
  NAND4_X1  g771(.A1(new_n1195), .A2(G319), .A3(new_n1196), .A4(new_n1197), .ZN(G225));
endmodule


