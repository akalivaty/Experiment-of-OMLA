//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 0 1 0 1 0 1 0 0 1 1 1 0 0 0 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  OR2_X1    g0004(.A1(KEYINPUT64), .A2(G20), .ZN(new_n205));
  NAND2_X1  g0005(.A1(KEYINPUT64), .A2(G20), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND3_X1  g0011(.A1(new_n207), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT0), .ZN(new_n216));
  XOR2_X1   g0016(.A(KEYINPUT65), .B(G77), .Z(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G97), .B2(G257), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G50), .A2(G226), .ZN(new_n224));
  NAND4_X1  g0024(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n213), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n212), .B(new_n216), .C1(new_n226), .C2(KEYINPUT1), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(G226), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G250), .B(G257), .Z(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G58), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  NOR2_X1   g0044(.A1(G20), .A2(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(G150), .ZN(new_n246));
  INV_X1    g0046(.A(G20), .ZN(new_n247));
  AND2_X1   g0047(.A1(KEYINPUT64), .A2(G20), .ZN(new_n248));
  NOR2_X1   g0048(.A1(KEYINPUT64), .A2(G20), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G33), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT8), .B(G58), .ZN(new_n252));
  OAI221_X1 g0052(.A(new_n246), .B1(new_n247), .B2(new_n201), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n208), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT67), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT67), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n254), .A2(new_n257), .A3(new_n208), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n253), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G1), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(G13), .A3(G20), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT68), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n262), .A2(KEYINPUT68), .A3(G13), .A4(G20), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G50), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n256), .A2(new_n258), .B1(new_n265), .B2(new_n266), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n262), .A2(G20), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n261), .B(new_n270), .C1(new_n269), .C2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT3), .ZN(new_n275));
  INV_X1    g0075(.A(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  AOI21_X1  g0078(.A(G1698), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AND2_X1   g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI22_X1  g0082(.A1(G222), .A2(new_n279), .B1(new_n217), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G223), .ZN(new_n284));
  INV_X1    g0084(.A(G1698), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n285), .B1(new_n277), .B2(new_n278), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n283), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(G33), .A2(G41), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n289), .A2(G1), .A3(G13), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G41), .ZN(new_n293));
  INV_X1    g0093(.A(G45), .ZN(new_n294));
  AOI21_X1  g0094(.A(G1), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G274), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n262), .B1(G41), .B2(G45), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n290), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n297), .B1(new_n300), .B2(G226), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n292), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n274), .B1(new_n302), .B2(G169), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT69), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI211_X1 g0105(.A(KEYINPUT69), .B(new_n274), .C1(new_n302), .C2(G169), .ZN(new_n306));
  INV_X1    g0106(.A(G179), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n305), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT70), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n305), .A2(KEYINPUT70), .A3(new_n306), .A4(new_n308), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n250), .A2(G33), .A3(G77), .ZN(new_n314));
  INV_X1    g0114(.A(G68), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n245), .A2(G50), .B1(G20), .B2(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n259), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  XOR2_X1   g0117(.A(new_n317), .B(KEYINPUT11), .Z(new_n318));
  INV_X1    g0118(.A(new_n273), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G68), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n268), .A2(new_n315), .ZN(new_n321));
  XNOR2_X1  g0121(.A(new_n321), .B(KEYINPUT12), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n318), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT13), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n279), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n325));
  INV_X1    g0125(.A(G232), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n325), .B1(new_n326), .B2(new_n287), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n291), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n297), .B1(new_n300), .B2(G238), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n324), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n328), .A2(new_n324), .A3(new_n329), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G200), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G190), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n331), .A2(new_n336), .A3(new_n332), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n323), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n332), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n339), .A2(new_n330), .ZN(new_n340));
  INV_X1    g0140(.A(G169), .ZN(new_n341));
  OAI21_X1  g0141(.A(KEYINPUT14), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT14), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n333), .A2(new_n343), .A3(G169), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n340), .A2(G179), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n342), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n338), .B1(new_n346), .B2(new_n323), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT9), .ZN(new_n348));
  OR2_X1    g0148(.A1(new_n274), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n274), .A2(new_n348), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n302), .A2(G190), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n292), .A2(new_n301), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(G200), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n349), .A2(new_n350), .A3(new_n351), .A4(new_n353), .ZN(new_n354));
  XNOR2_X1  g0154(.A(new_n354), .B(KEYINPUT10), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n217), .A2(new_n207), .ZN(new_n356));
  INV_X1    g0156(.A(new_n245), .ZN(new_n357));
  XNOR2_X1  g0157(.A(KEYINPUT15), .B(G87), .ZN(new_n358));
  OAI221_X1 g0158(.A(new_n356), .B1(new_n357), .B2(new_n252), .C1(new_n251), .C2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n260), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n271), .A2(G77), .A3(new_n272), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n268), .A2(new_n218), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT71), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n279), .A2(G232), .B1(new_n282), .B2(G107), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n286), .A2(G238), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n290), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n296), .B1(new_n299), .B2(new_n219), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n341), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n363), .A2(new_n364), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n365), .A2(new_n366), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n368), .B1(new_n371), .B2(new_n291), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n307), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n364), .B1(new_n363), .B2(new_n369), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n372), .A2(G200), .ZN(new_n377));
  NOR3_X1   g0177(.A1(new_n367), .A2(G190), .A3(new_n368), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n379), .A2(new_n363), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n313), .A2(new_n347), .A3(new_n355), .A4(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT17), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n290), .A2(G232), .A3(new_n298), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n384), .A2(KEYINPUT74), .A3(new_n296), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT74), .B1(new_n384), .B2(new_n296), .ZN(new_n387));
  NOR3_X1   g0187(.A1(new_n386), .A2(new_n387), .A3(G190), .ZN(new_n388));
  OAI211_X1 g0188(.A(G223), .B(new_n285), .C1(new_n280), .C2(new_n281), .ZN(new_n389));
  OAI211_X1 g0189(.A(G226), .B(G1698), .C1(new_n280), .C2(new_n281), .ZN(new_n390));
  INV_X1    g0190(.A(G87), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n389), .B(new_n390), .C1(new_n276), .C2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n291), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(KEYINPUT73), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT73), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n392), .A2(new_n395), .A3(new_n291), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n388), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n387), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n393), .A2(new_n398), .A3(new_n385), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n334), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT75), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n397), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT7), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n277), .A2(new_n278), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n403), .B1(new_n207), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n282), .A2(KEYINPUT7), .A3(new_n247), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G68), .ZN(new_n408));
  INV_X1    g0208(.A(G58), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n409), .A2(new_n315), .ZN(new_n410));
  NOR2_X1   g0210(.A1(G58), .A2(G68), .ZN(new_n411));
  OAI21_X1  g0211(.A(G20), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n245), .A2(G159), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n408), .A2(KEYINPUT16), .A3(new_n415), .ZN(new_n416));
  XNOR2_X1  g0216(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n403), .B1(new_n404), .B2(G20), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n250), .A2(new_n282), .A3(KEYINPUT7), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n315), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n417), .B1(new_n420), .B2(new_n414), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n416), .A2(new_n421), .A3(new_n260), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n267), .A2(new_n252), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(new_n319), .B2(new_n252), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n402), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n401), .B1(new_n397), .B2(new_n400), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n383), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n422), .A2(new_n424), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  NOR3_X1   g0229(.A1(new_n386), .A2(new_n387), .A3(G179), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n430), .A2(new_n394), .A3(new_n396), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n399), .A2(new_n341), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT18), .B1(new_n429), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n397), .A2(new_n400), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT75), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n429), .A2(new_n436), .A3(KEYINPUT17), .A4(new_n402), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n431), .A2(new_n432), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT18), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(new_n428), .A3(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n427), .A2(new_n434), .A3(new_n437), .A4(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n382), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(G274), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n294), .A2(G1), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n443), .A2(new_n444), .B1(new_n209), .B2(new_n289), .ZN(new_n445));
  OR2_X1    g0245(.A1(new_n444), .A2(G250), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI211_X1 g0247(.A(G238), .B(new_n285), .C1(new_n280), .C2(new_n281), .ZN(new_n448));
  NAND2_X1  g0248(.A1(G33), .A2(G116), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT80), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT79), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n452), .B1(new_n286), .B2(G244), .ZN(new_n453));
  OAI211_X1 g0253(.A(G244), .B(G1698), .C1(new_n280), .C2(new_n281), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(KEYINPUT79), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n450), .B(new_n451), .C1(new_n453), .C2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n291), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n448), .A2(new_n449), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n286), .A2(new_n452), .A3(G244), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n454), .A2(KEYINPUT79), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(new_n451), .ZN(new_n462));
  OAI211_X1 g0262(.A(G190), .B(new_n447), .C1(new_n457), .C2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(G97), .ZN(new_n464));
  INV_X1    g0264(.A(G107), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n391), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT19), .ZN(new_n467));
  NOR3_X1   g0267(.A1(new_n467), .A2(new_n276), .A3(new_n464), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n466), .B1(new_n468), .B2(new_n207), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n205), .A2(G33), .A3(G97), .A4(new_n206), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n467), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n404), .A2(new_n250), .A3(G68), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n469), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n473), .A2(new_n260), .B1(new_n268), .B2(new_n358), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n262), .A2(G33), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n271), .A2(G87), .A3(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT81), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n271), .A2(KEYINPUT81), .A3(G87), .A4(new_n475), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n474), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n290), .B1(new_n461), .B2(new_n451), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n450), .B1(new_n453), .B2(new_n455), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT80), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n481), .A2(new_n483), .B1(new_n445), .B2(new_n446), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n463), .B(new_n480), .C1(new_n484), .C2(new_n334), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n307), .B(new_n447), .C1(new_n457), .C2(new_n462), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n271), .A2(new_n475), .ZN(new_n487));
  INV_X1    g0287(.A(new_n358), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n474), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n486), .B(new_n490), .C1(new_n484), .C2(G169), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n485), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT6), .ZN(new_n493));
  NOR3_X1   g0293(.A1(new_n493), .A2(new_n464), .A3(G107), .ZN(new_n494));
  XNOR2_X1  g0294(.A(G97), .B(G107), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n494), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  OAI22_X1  g0296(.A1(new_n496), .A2(new_n250), .B1(new_n202), .B2(new_n357), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n465), .B1(new_n418), .B2(new_n419), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n260), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n487), .A2(G97), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n268), .A2(new_n464), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AND2_X1   g0302(.A1(KEYINPUT4), .A2(G244), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n285), .B(new_n503), .C1(new_n280), .C2(new_n281), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G283), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n219), .B1(new_n277), .B2(new_n278), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n504), .B(new_n505), .C1(new_n506), .C2(KEYINPUT4), .ZN(new_n507));
  OAI21_X1  g0307(.A(G250), .B1(new_n280), .B2(new_n281), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n285), .B1(new_n508), .B2(KEYINPUT4), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n291), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT77), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT5), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n511), .B1(new_n512), .B2(G41), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  AND2_X1   g0314(.A1(KEYINPUT76), .A2(KEYINPUT5), .ZN(new_n515));
  NOR2_X1   g0315(.A1(KEYINPUT76), .A2(KEYINPUT5), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n293), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(KEYINPUT77), .B(new_n293), .C1(new_n515), .C2(new_n516), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n518), .A2(new_n445), .A3(new_n519), .A4(new_n444), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n444), .ZN(new_n521));
  XNOR2_X1  g0321(.A(KEYINPUT76), .B(KEYINPUT5), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n513), .B1(new_n522), .B2(new_n293), .ZN(new_n523));
  OAI211_X1 g0323(.A(G257), .B(new_n290), .C1(new_n521), .C2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n510), .A2(new_n520), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n341), .ZN(new_n526));
  AND2_X1   g0326(.A1(new_n502), .A2(new_n526), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n524), .A2(new_n520), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT78), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n528), .A2(new_n529), .A3(new_n307), .A4(new_n510), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n510), .A2(new_n307), .A3(new_n524), .A4(new_n520), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(KEYINPUT78), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n525), .A2(new_n334), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(G190), .B2(new_n525), .ZN(new_n535));
  AND3_X1   g0335(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n527), .A2(new_n533), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n492), .A2(KEYINPUT82), .A3(new_n537), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n531), .A2(KEYINPUT78), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n531), .A2(KEYINPUT78), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n526), .B(new_n502), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(G200), .B1(new_n528), .B2(new_n510), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n525), .A2(G190), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n536), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n541), .A2(new_n485), .A3(new_n491), .A4(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT82), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI211_X1 g0347(.A(G270), .B(new_n290), .C1(new_n521), .C2(new_n523), .ZN(new_n548));
  OAI211_X1 g0348(.A(G264), .B(G1698), .C1(new_n280), .C2(new_n281), .ZN(new_n549));
  OAI211_X1 g0349(.A(G257), .B(new_n285), .C1(new_n280), .C2(new_n281), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n277), .A2(G303), .A3(new_n278), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT83), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n552), .A2(new_n553), .A3(new_n291), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n553), .B1(new_n552), .B2(new_n291), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n520), .B(new_n548), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n276), .A2(G97), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n205), .A2(new_n558), .A3(new_n206), .A4(new_n505), .ZN(new_n559));
  INV_X1    g0359(.A(G116), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n254), .A2(new_n208), .B1(G20), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT20), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n559), .A2(KEYINPUT20), .A3(new_n561), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n564), .A2(new_n565), .B1(new_n560), .B2(new_n268), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n271), .A2(G116), .A3(new_n475), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n341), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n557), .A2(new_n568), .A3(KEYINPUT21), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n566), .A2(new_n567), .ZN(new_n570));
  AND2_X1   g0370(.A1(new_n548), .A2(new_n520), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n552), .A2(new_n291), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(KEYINPUT83), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n554), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n570), .A2(new_n571), .A3(new_n574), .A4(G179), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n569), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT21), .B1(new_n557), .B2(new_n568), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n271), .A2(G107), .A3(new_n475), .ZN(new_n579));
  OR3_X1    g0379(.A1(new_n267), .A2(KEYINPUT25), .A3(G107), .ZN(new_n580));
  OAI21_X1  g0380(.A(KEYINPUT25), .B1(new_n267), .B2(G107), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n404), .A2(new_n250), .A3(G87), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(KEYINPUT22), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT22), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n404), .A2(new_n250), .A3(new_n585), .A4(G87), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT85), .ZN(new_n588));
  NOR2_X1   g0388(.A1(KEYINPUT23), .A2(G107), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n207), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n589), .B1(new_n248), .B2(new_n249), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT85), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT23), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n449), .A2(new_n593), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n594), .A2(new_n247), .B1(KEYINPUT23), .B2(G107), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n590), .A2(new_n592), .A3(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n587), .A2(new_n596), .A3(KEYINPUT24), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n260), .ZN(new_n598));
  AOI21_X1  g0398(.A(KEYINPUT24), .B1(new_n587), .B2(new_n596), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n582), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OAI211_X1 g0400(.A(G264), .B(new_n290), .C1(new_n521), .C2(new_n523), .ZN(new_n601));
  OAI211_X1 g0401(.A(G257), .B(G1698), .C1(new_n280), .C2(new_n281), .ZN(new_n602));
  NAND2_X1  g0402(.A1(G33), .A2(G294), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n602), .B(new_n603), .C1(new_n508), .C2(G1698), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n291), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n601), .A2(new_n605), .A3(new_n520), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(G169), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n607), .B1(new_n307), .B2(new_n606), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n600), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n606), .A2(new_n334), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n601), .A2(new_n605), .A3(new_n336), .A4(new_n520), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n587), .A2(new_n596), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT24), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n615), .A2(new_n260), .A3(new_n597), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n612), .A2(new_n616), .A3(new_n582), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n609), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n570), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n557), .A2(G190), .ZN(new_n620));
  AOI21_X1  g0420(.A(G200), .B1(new_n571), .B2(new_n574), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(KEYINPUT84), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT84), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n624), .B(new_n619), .C1(new_n620), .C2(new_n621), .ZN(new_n625));
  AND4_X1   g0425(.A1(new_n578), .A2(new_n618), .A3(new_n623), .A4(new_n625), .ZN(new_n626));
  AND4_X1   g0426(.A1(new_n442), .A2(new_n538), .A3(new_n547), .A4(new_n626), .ZN(G372));
  INV_X1    g0427(.A(new_n617), .ZN(new_n628));
  OAI21_X1  g0428(.A(KEYINPUT86), .B1(new_n545), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT86), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n492), .A2(new_n630), .A3(new_n537), .A4(new_n617), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n557), .A2(new_n568), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT21), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n635), .A2(new_n569), .A3(new_n575), .ZN(new_n636));
  INV_X1    g0436(.A(new_n609), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n632), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT26), .ZN(new_n641));
  INV_X1    g0441(.A(new_n541), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n492), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n485), .A2(new_n491), .ZN(new_n644));
  OAI21_X1  g0444(.A(KEYINPUT26), .B1(new_n644), .B2(new_n541), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n643), .A2(new_n645), .A3(new_n491), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n640), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n442), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n338), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n649), .A2(new_n427), .A3(new_n437), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n376), .B1(new_n346), .B2(new_n323), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n434), .B(new_n440), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n652), .A2(new_n355), .B1(new_n311), .B2(new_n312), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n648), .A2(new_n653), .ZN(G369));
  AND3_X1   g0454(.A1(new_n623), .A2(new_n578), .A3(new_n625), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n250), .A2(new_n262), .A3(G13), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(G213), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(G343), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(new_n619), .ZN(new_n663));
  MUX2_X1   g0463(.A(new_n655), .B(new_n636), .S(new_n663), .Z(new_n664));
  AND2_X1   g0464(.A1(new_n664), .A2(G330), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n600), .A2(new_n661), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n637), .B1(new_n617), .B2(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n609), .A2(new_n661), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n636), .A2(new_n662), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n668), .B1(new_n669), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n670), .A2(new_n673), .ZN(G399));
  INV_X1    g0474(.A(new_n214), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(G41), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(new_n262), .ZN(new_n677));
  NOR4_X1   g0477(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n678));
  AOI22_X1  g0478(.A1(new_n677), .A2(new_n678), .B1(new_n211), .B2(new_n676), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n679), .B(KEYINPUT87), .ZN(new_n680));
  XOR2_X1   g0480(.A(new_n680), .B(KEYINPUT28), .Z(new_n681));
  AND2_X1   g0481(.A1(new_n525), .A2(new_n606), .ZN(new_n682));
  INV_X1    g0482(.A(new_n484), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n682), .A2(new_n683), .A3(new_n307), .A4(new_n557), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT88), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n684), .B(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n557), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n601), .A2(new_n605), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n525), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n687), .A2(new_n484), .A3(G179), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT30), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n662), .B1(new_n686), .B2(new_n691), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n626), .A2(new_n538), .A3(new_n547), .A4(new_n662), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n692), .B1(new_n693), .B2(KEYINPUT31), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT31), .ZN(new_n695));
  AOI211_X1 g0495(.A(new_n695), .B(new_n662), .C1(new_n691), .C2(new_n684), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G330), .ZN(new_n698));
  OAI21_X1  g0498(.A(KEYINPUT89), .B1(new_n636), .B2(new_n637), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT89), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n578), .A2(new_n700), .A3(new_n609), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n545), .A2(new_n628), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n643), .A2(new_n645), .A3(new_n491), .ZN(new_n705));
  OAI211_X1 g0505(.A(KEYINPUT29), .B(new_n662), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n661), .B1(new_n640), .B2(new_n646), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n706), .B1(new_n707), .B2(KEYINPUT29), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n698), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n681), .B1(new_n709), .B2(G1), .ZN(new_n710));
  XOR2_X1   g0510(.A(new_n710), .B(KEYINPUT90), .Z(G364));
  INV_X1    g0511(.A(G13), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n207), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G45), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n677), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n675), .A2(new_n282), .ZN(new_n716));
  XNOR2_X1  g0516(.A(G355), .B(KEYINPUT91), .ZN(new_n717));
  AOI22_X1  g0517(.A1(new_n716), .A2(new_n717), .B1(new_n560), .B2(new_n675), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n211), .A2(G45), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n719), .B1(new_n240), .B2(G45), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n675), .A2(new_n404), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n718), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(G13), .A2(G33), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G20), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n208), .B1(G20), .B2(new_n341), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n715), .B1(new_n723), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n207), .A2(new_n336), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n731), .A2(new_n307), .A3(G200), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n732), .A2(KEYINPUT94), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(KEYINPUT94), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G107), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G179), .A2(G200), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G190), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n207), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  OR2_X1    g0542(.A1(new_n742), .A2(KEYINPUT95), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(KEYINPUT95), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n464), .ZN(new_n746));
  NOR4_X1   g0546(.A1(new_n247), .A2(new_n336), .A3(new_n334), .A4(G179), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n730), .A2(new_n307), .A3(G200), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OAI221_X1 g0550(.A(new_n404), .B1(new_n391), .B2(new_n748), .C1(new_n750), .C2(new_n218), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n738), .A2(new_n746), .A3(new_n751), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n207), .A2(G179), .A3(G190), .A4(new_n334), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(KEYINPUT92), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n753), .A2(KEYINPUT92), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n731), .A2(new_n739), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n760), .A2(KEYINPUT32), .A3(G159), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT32), .ZN(new_n762));
  INV_X1    g0562(.A(G159), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n762), .B1(new_n759), .B2(new_n763), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n758), .A2(G58), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n207), .A2(G179), .A3(G200), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT93), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n766), .A2(new_n767), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n768), .A2(G190), .A3(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n768), .A2(new_n336), .A3(new_n769), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI22_X1  g0573(.A1(G50), .A2(new_n771), .B1(new_n773), .B2(G68), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n752), .A2(new_n765), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT96), .ZN(new_n776));
  INV_X1    g0576(.A(G322), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n757), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n760), .A2(G329), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n404), .B1(new_n747), .B2(G303), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n749), .A2(G311), .B1(new_n780), .B2(KEYINPUT98), .ZN(new_n781));
  OAI211_X1 g0581(.A(new_n779), .B(new_n781), .C1(KEYINPUT98), .C2(new_n780), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n778), .B(new_n782), .C1(G283), .C2(new_n736), .ZN(new_n783));
  INV_X1    g0583(.A(G326), .ZN(new_n784));
  INV_X1    g0584(.A(G294), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n770), .A2(new_n784), .B1(new_n785), .B2(new_n742), .ZN(new_n786));
  INV_X1    g0586(.A(KEYINPUT97), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n786), .A2(new_n787), .ZN(new_n789));
  XNOR2_X1  g0589(.A(KEYINPUT33), .B(G317), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n773), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n783), .A2(new_n788), .A3(new_n789), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n776), .A2(new_n792), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n793), .A2(KEYINPUT99), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n727), .B1(new_n793), .B2(KEYINPUT99), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n729), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT100), .ZN(new_n797));
  INV_X1    g0597(.A(new_n726), .ZN(new_n798));
  OR2_X1    g0598(.A1(new_n664), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n715), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n665), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(G330), .B2(new_n664), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(G396));
  AOI22_X1  g0605(.A1(new_n758), .A2(G143), .B1(G159), .B2(new_n749), .ZN(new_n806));
  INV_X1    g0606(.A(G137), .ZN(new_n807));
  INV_X1    g0607(.A(G150), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n806), .B1(new_n807), .B2(new_n770), .C1(new_n808), .C2(new_n772), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT34), .Z(new_n810));
  OAI21_X1  g0610(.A(new_n404), .B1(new_n748), .B2(new_n269), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(G58), .B2(new_n741), .ZN(new_n812));
  INV_X1    g0612(.A(G132), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n812), .B1(new_n813), .B2(new_n759), .C1(new_n735), .C2(new_n315), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n736), .A2(G87), .ZN(new_n816));
  INV_X1    g0616(.A(G311), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n816), .B1(new_n817), .B2(new_n759), .ZN(new_n818));
  XOR2_X1   g0618(.A(new_n818), .B(KEYINPUT102), .Z(new_n819));
  OAI221_X1 g0619(.A(new_n282), .B1(new_n465), .B2(new_n748), .C1(new_n750), .C2(new_n560), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n746), .B(new_n820), .C1(G294), .C2(new_n758), .ZN(new_n821));
  INV_X1    g0621(.A(G283), .ZN(new_n822));
  INV_X1    g0622(.A(G303), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n821), .B1(new_n822), .B2(new_n772), .C1(new_n823), .C2(new_n770), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n819), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n727), .B1(new_n815), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n727), .A2(new_n724), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n801), .B1(G77), .B2(new_n828), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT101), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT103), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n363), .A2(new_n661), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n379), .B2(new_n363), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n374), .B2(new_n375), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT104), .ZN(new_n836));
  INV_X1    g0636(.A(new_n375), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n837), .A2(new_n370), .A3(new_n373), .A4(new_n833), .ZN(new_n838));
  AND3_X1   g0638(.A1(new_n835), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n836), .B1(new_n835), .B2(new_n838), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n832), .B1(new_n725), .B2(new_n841), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT105), .ZN(new_n843));
  INV_X1    g0643(.A(new_n698), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n707), .A2(new_n841), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n638), .B1(new_n629), .B2(new_n631), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n662), .B(new_n841), .C1(new_n846), .C2(new_n705), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n801), .B1(new_n844), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n848), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n850), .B1(new_n698), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n843), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(G384));
  INV_X1    g0654(.A(new_n496), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n855), .A2(KEYINPUT35), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n855), .A2(KEYINPUT35), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n207), .A2(G116), .A3(new_n209), .ZN(new_n858));
  NOR3_X1   g0658(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  OR2_X1    g0659(.A1(new_n859), .A2(KEYINPUT36), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(KEYINPUT36), .ZN(new_n861));
  NOR3_X1   g0661(.A1(new_n218), .A2(new_n210), .A3(new_n410), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n315), .A2(G50), .ZN(new_n863));
  OAI211_X1 g0663(.A(G1), .B(new_n712), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n860), .A2(new_n861), .A3(new_n864), .ZN(new_n865));
  XOR2_X1   g0665(.A(new_n865), .B(KEYINPUT106), .Z(new_n866));
  INV_X1    g0666(.A(new_n417), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n414), .B1(new_n407), .B2(G68), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n416), .B(new_n260), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n659), .B1(new_n869), .B2(new_n424), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n441), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n425), .A2(new_n426), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n433), .A2(new_n659), .B1(new_n869), .B2(new_n424), .ZN(new_n873));
  OAI21_X1  g0673(.A(KEYINPUT37), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT107), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n659), .B(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n428), .B1(new_n438), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT37), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n877), .B(new_n878), .C1(new_n426), .C2(new_n425), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n874), .A2(new_n879), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n871), .A2(new_n880), .A3(KEYINPUT38), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT38), .B1(new_n871), .B2(new_n880), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT39), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n876), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n429), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n441), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n877), .B1(new_n426), .B2(new_n425), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT37), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n879), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT38), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT39), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n871), .A2(new_n880), .A3(KEYINPUT38), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n883), .A2(new_n895), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n346), .A2(new_n323), .A3(new_n662), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n376), .A2(new_n662), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n847), .A2(new_n899), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n323), .A2(new_n661), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n347), .B(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n900), .B(new_n903), .C1(new_n882), .C2(new_n881), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n434), .A2(new_n440), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n884), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n898), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n442), .B(new_n706), .C1(new_n707), .C2(KEYINPUT29), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n653), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n907), .B(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT40), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n686), .A2(new_n691), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n661), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n913), .A2(new_n695), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n903), .B(new_n841), .C1(new_n694), .C2(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n881), .A2(new_n882), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n911), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n693), .A2(KEYINPUT31), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n913), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n692), .A2(KEYINPUT31), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n911), .B1(new_n892), .B2(new_n894), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n921), .A2(new_n841), .A3(new_n903), .A4(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n917), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n921), .A2(new_n442), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n924), .B(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(G330), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n910), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n262), .B2(new_n713), .ZN(new_n929));
  NOR3_X1   g0729(.A1(new_n926), .A2(new_n910), .A3(new_n927), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n866), .B1(new_n929), .B2(new_n930), .ZN(G367));
  OAI21_X1  g0731(.A(new_n537), .B1(new_n536), .B2(new_n662), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n642), .A2(new_n661), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n669), .A2(new_n934), .A3(new_n672), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n935), .A2(KEYINPUT42), .ZN(new_n936));
  INV_X1    g0736(.A(new_n544), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n541), .B1(new_n937), .B2(new_n609), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n935), .A2(KEYINPUT42), .B1(new_n662), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n480), .A2(new_n662), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n492), .A2(new_n940), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n491), .A2(new_n940), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n936), .A2(new_n939), .B1(KEYINPUT43), .B2(new_n943), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n943), .A2(KEYINPUT43), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n945), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n934), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n670), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n948), .B(new_n950), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n676), .B(KEYINPUT41), .Z(new_n952));
  INV_X1    g0752(.A(KEYINPUT44), .ZN(new_n953));
  INV_X1    g0753(.A(new_n673), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n953), .B1(new_n954), .B2(new_n949), .ZN(new_n955));
  NOR3_X1   g0755(.A1(new_n673), .A2(KEYINPUT44), .A3(new_n934), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT45), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n954), .B2(new_n949), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n673), .A2(KEYINPUT45), .A3(new_n934), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT108), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n665), .A2(new_n962), .A3(new_n669), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n957), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n964), .A2(KEYINPUT108), .A3(new_n670), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n670), .A2(KEYINPUT108), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n966), .A2(new_n957), .A3(new_n961), .A4(new_n963), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n669), .B(new_n672), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n665), .B(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n968), .A2(new_n709), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n952), .B1(new_n971), .B2(new_n709), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n714), .A2(G1), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n951), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n236), .A2(new_n722), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n728), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(new_n675), .B2(new_n488), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n715), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n404), .B1(new_n409), .B2(new_n748), .C1(new_n759), .C2(new_n807), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n745), .A2(new_n315), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n980), .B(new_n981), .C1(G50), .C2(new_n749), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n736), .A2(new_n217), .B1(G150), .B2(new_n758), .ZN(new_n983));
  AOI22_X1  g0783(.A1(G143), .A2(new_n771), .B1(new_n773), .B2(G159), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n736), .A2(G97), .B1(G303), .B2(new_n758), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n748), .A2(new_n560), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(KEYINPUT46), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT109), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n282), .B1(new_n465), .B2(new_n742), .C1(new_n987), .C2(KEYINPUT46), .ZN(new_n990));
  INV_X1    g0790(.A(G317), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n750), .A2(new_n822), .B1(new_n759), .B2(new_n991), .ZN(new_n992));
  NOR3_X1   g0792(.A1(new_n989), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  AOI22_X1  g0793(.A1(G294), .A2(new_n773), .B1(new_n771), .B2(G311), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n986), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n985), .A2(KEYINPUT47), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n727), .ZN(new_n997));
  AOI21_X1  g0797(.A(KEYINPUT47), .B1(new_n985), .B2(new_n995), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n979), .B1(new_n997), .B2(new_n998), .C1(new_n798), .C2(new_n943), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n974), .A2(new_n999), .ZN(G387));
  INV_X1    g0800(.A(new_n716), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n1001), .A2(new_n678), .B1(G107), .B2(new_n214), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n233), .A2(G45), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n678), .B(new_n294), .C1(new_n315), .C2(new_n202), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT110), .Z(new_n1005));
  NOR2_X1   g0805(.A1(new_n252), .A2(G50), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n722), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1002), .B1(new_n1003), .B2(new_n1009), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n801), .B1(new_n977), .B2(new_n1010), .C1(new_n669), .C2(new_n798), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n735), .A2(new_n464), .B1(new_n269), .B2(new_n757), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n748), .A2(new_n218), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n282), .B(new_n1013), .C1(new_n749), .C2(G68), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n808), .B2(new_n759), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n745), .A2(new_n358), .ZN(new_n1016));
  NOR3_X1   g0816(.A1(new_n1012), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1017), .B1(new_n763), .B2(new_n770), .C1(new_n252), .C2(new_n772), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n817), .A2(new_n772), .B1(new_n770), .B2(new_n777), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT112), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n757), .A2(new_n991), .B1(new_n823), .B2(new_n750), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(KEYINPUT48), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1022), .A2(KEYINPUT48), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n742), .A2(new_n822), .B1(new_n748), .B2(new_n785), .ZN(new_n1026));
  NOR3_X1   g0826(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(KEYINPUT49), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n404), .B1(new_n760), .B2(G326), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1028), .B(new_n1029), .C1(new_n560), .C2(new_n735), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1027), .A2(KEYINPUT49), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1018), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1011), .B1(new_n1032), .B2(new_n727), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1033), .A2(KEYINPUT113), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(KEYINPUT113), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n1034), .A2(new_n1035), .B1(new_n970), .B2(new_n973), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n676), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n709), .B2(new_n970), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n709), .B2(new_n970), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1036), .A2(new_n1039), .ZN(G393));
  NAND2_X1  g0840(.A1(new_n709), .A2(new_n970), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1041), .A2(new_n965), .A3(new_n967), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n971), .A2(new_n1042), .A3(new_n676), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n404), .B1(new_n315), .B2(new_n748), .C1(new_n750), .C2(new_n252), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(G143), .B2(new_n760), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n745), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(G77), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n816), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n757), .A2(new_n763), .B1(new_n770), .B2(new_n808), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT51), .Z(new_n1050));
  AOI211_X1 g0850(.A(new_n1048), .B(new_n1050), .C1(G50), .C2(new_n773), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n757), .A2(new_n817), .B1(new_n770), .B2(new_n991), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT52), .Z(new_n1053));
  NOR2_X1   g0853(.A1(new_n772), .A2(new_n823), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n282), .B1(new_n748), .B2(new_n822), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(G116), .B2(new_n741), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1056), .B1(new_n777), .B2(new_n759), .C1(new_n785), .C2(new_n750), .ZN(new_n1057));
  NOR4_X1   g0857(.A1(new_n1053), .A2(new_n738), .A3(new_n1054), .A4(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n727), .B1(new_n1051), .B2(new_n1058), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n728), .B1(new_n464), .B2(new_n214), .C1(new_n243), .C2(new_n722), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1059), .A2(new_n801), .A3(new_n1060), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT114), .Z(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n726), .B2(new_n949), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(new_n968), .B2(new_n973), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1043), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(KEYINPUT115), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT115), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1043), .A2(new_n1067), .A3(new_n1064), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1066), .A2(new_n1068), .ZN(G390));
  NAND4_X1  g0869(.A1(new_n921), .A2(G330), .A3(new_n841), .A4(new_n903), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n902), .B1(new_n847), .B2(new_n899), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n883), .B(new_n895), .C1(new_n1071), .C2(new_n897), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n897), .B1(new_n892), .B2(new_n894), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n899), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n702), .A2(new_n703), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n661), .B1(new_n646), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1074), .B1(new_n1076), .B2(new_n841), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1073), .B1(new_n1077), .B2(new_n902), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1070), .B1(new_n1072), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n897), .B1(new_n900), .B2(new_n903), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1078), .B1(new_n1080), .B2(new_n896), .ZN(new_n1081));
  OAI211_X1 g0881(.A(G330), .B(new_n841), .C1(new_n694), .C2(new_n696), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1082), .A2(new_n902), .ZN(new_n1083));
  OAI21_X1  g0883(.A(KEYINPUT116), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n1082), .A2(new_n902), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT116), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1085), .A2(new_n1086), .A3(new_n1072), .A4(new_n1078), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1079), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n973), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT119), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1088), .A2(KEYINPUT119), .A3(new_n973), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n883), .A2(new_n895), .A3(new_n724), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n827), .A2(new_n252), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n282), .B1(new_n760), .B2(G125), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n747), .A2(G150), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT53), .Z(new_n1097));
  XOR2_X1   g0897(.A(KEYINPUT54), .B(G143), .Z(new_n1098));
  NAND2_X1  g0898(.A1(new_n749), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1095), .A2(new_n1097), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(G159), .B2(new_n1046), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n736), .A2(G50), .B1(G132), .B2(new_n758), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(G128), .A2(new_n771), .B1(new_n773), .B2(G137), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  OR2_X1    g0905(.A1(new_n1105), .A2(KEYINPUT120), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(KEYINPUT120), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n736), .A2(G68), .B1(G116), .B2(new_n758), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n282), .B1(new_n391), .B2(new_n748), .C1(new_n759), .C2(new_n785), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(G97), .B2(new_n749), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(G107), .A2(new_n773), .B1(new_n771), .B2(G283), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1108), .A2(new_n1047), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1106), .A2(new_n1107), .A3(new_n1112), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n715), .B(new_n1094), .C1(new_n1113), .C2(new_n727), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1091), .A2(new_n1092), .B1(new_n1093), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1079), .ZN(new_n1117));
  OAI211_X1 g0917(.A(G330), .B(new_n442), .C1(new_n694), .C2(new_n914), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n908), .A2(new_n1118), .A3(new_n653), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT117), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n908), .A2(new_n1118), .A3(KEYINPUT117), .A4(new_n653), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n1082), .A2(new_n902), .ZN(new_n1124));
  OAI211_X1 g0924(.A(G330), .B(new_n841), .C1(new_n694), .C2(new_n914), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1125), .A2(new_n902), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n900), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1125), .A2(new_n902), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1085), .A2(new_n1077), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1116), .A2(new_n1117), .A3(new_n1123), .A4(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1128), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1077), .B1(new_n1082), .B2(new_n902), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n900), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1082), .A2(new_n902), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1135), .B1(new_n1070), .B2(new_n1136), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1121), .B(new_n1122), .C1(new_n1134), .C2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(KEYINPUT118), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT118), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1130), .A2(new_n1123), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n676), .B(new_n1131), .C1(new_n1142), .C2(new_n1088), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1115), .A2(new_n1143), .ZN(G378));
  INV_X1    g0944(.A(KEYINPUT57), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1131), .A2(new_n1123), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n659), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n274), .A2(new_n1147), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n355), .A2(new_n309), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1148), .B1(new_n355), .B2(new_n309), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT122), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  OR3_X1    g0953(.A1(new_n1149), .A2(new_n1150), .A3(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1153), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n907), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n917), .A2(G330), .A3(new_n923), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1156), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n898), .A2(new_n1159), .A3(new_n904), .A4(new_n906), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n1157), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1158), .B1(new_n1157), .B2(new_n1160), .ZN(new_n1162));
  OR2_X1    g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1145), .B1(new_n1146), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(new_n1088), .B2(new_n1130), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n1166), .A2(new_n1167), .A3(KEYINPUT57), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n676), .B1(new_n1164), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1159), .A2(new_n724), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n801), .B1(G50), .B2(new_n828), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n757), .A2(new_n465), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT121), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1173), .B1(new_n464), .B2(new_n772), .C1(new_n560), .C2(new_n770), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n735), .A2(new_n409), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n282), .A2(new_n293), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n1013), .B(new_n1176), .C1(new_n760), .C2(G283), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n358), .B2(new_n750), .ZN(new_n1178));
  NOR4_X1   g0978(.A1(new_n1174), .A2(new_n981), .A3(new_n1175), .A4(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(G50), .B1(new_n276), .B2(new_n293), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n1179), .A2(KEYINPUT58), .B1(new_n1176), .B2(new_n1180), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n749), .A2(G137), .B1(new_n747), .B2(new_n1098), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n745), .B2(new_n808), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(G128), .B2(new_n758), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n771), .A2(G125), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1184), .B(new_n1185), .C1(new_n813), .C2(new_n772), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1186), .A2(KEYINPUT59), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(KEYINPUT59), .ZN(new_n1188));
  AOI211_X1 g0988(.A(G33), .B(G41), .C1(new_n760), .C2(G124), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1188), .B(new_n1189), .C1(new_n763), .C2(new_n735), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1181), .B1(KEYINPUT58), .B2(new_n1179), .C1(new_n1187), .C2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1171), .B1(new_n1191), .B2(new_n727), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1163), .A2(new_n973), .B1(new_n1170), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1169), .A2(new_n1193), .ZN(G375));
  NOR2_X1   g0994(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n952), .B1(new_n1195), .B2(new_n1165), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1139), .A2(new_n1196), .A3(new_n1141), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n902), .A2(new_n724), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n801), .B1(G68), .B2(new_n828), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n735), .A2(new_n202), .B1(new_n822), .B2(new_n757), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n404), .B1(new_n747), .B2(G97), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1201), .B1(new_n759), .B2(new_n823), .C1(new_n750), .C2(new_n465), .ZN(new_n1202));
  NOR3_X1   g1002(.A1(new_n1200), .A2(new_n1016), .A3(new_n1202), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1203), .B1(new_n560), .B2(new_n772), .C1(new_n785), .C2(new_n770), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n757), .A2(new_n807), .B1(new_n770), .B2(new_n813), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(new_n773), .B2(new_n1098), .ZN(new_n1206));
  XOR2_X1   g1006(.A(new_n1206), .B(KEYINPUT123), .Z(new_n1207));
  OAI221_X1 g1007(.A(new_n404), .B1(new_n763), .B2(new_n748), .C1(new_n750), .C2(new_n808), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(G128), .B2(new_n760), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1209), .B1(new_n269), .B2(new_n745), .C1(new_n409), .C2(new_n735), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1204), .B1(new_n1207), .B2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1199), .B1(new_n1211), .B2(new_n727), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1130), .A2(new_n973), .B1(new_n1198), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1197), .A2(new_n1213), .ZN(G381));
  NAND4_X1  g1014(.A1(new_n1066), .A2(new_n974), .A3(new_n999), .A4(new_n1068), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n804), .A2(new_n1039), .A3(new_n1036), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1216), .A2(new_n853), .A3(new_n1218), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1169), .A2(new_n1143), .A3(new_n1115), .A4(new_n1193), .ZN(new_n1220));
  OR3_X1    g1020(.A1(new_n1219), .A2(new_n1220), .A3(G381), .ZN(G407));
  OAI211_X1 g1021(.A(G407), .B(G213), .C1(G343), .C2(new_n1220), .ZN(G409));
  NAND3_X1  g1022(.A1(new_n1169), .A2(G378), .A3(new_n1193), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1193), .ZN(new_n1224));
  NOR3_X1   g1024(.A1(new_n1166), .A2(new_n1167), .A3(new_n952), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1115), .B(new_n1143), .C1(new_n1224), .C2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1223), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(G213), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1228), .A2(G343), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT124), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1165), .A2(KEYINPUT60), .A3(new_n1127), .A4(new_n1129), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1232), .A2(new_n1138), .A3(new_n676), .ZN(new_n1233));
  AOI21_X1  g1033(.A(KEYINPUT60), .B1(new_n1195), .B2(new_n1165), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1231), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT60), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n1130), .B2(new_n1123), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1037), .B1(new_n1130), .B2(new_n1123), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1237), .A2(new_n1238), .A3(KEYINPUT124), .A4(new_n1232), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1235), .A2(new_n1213), .A3(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n853), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(G384), .A2(new_n1213), .A3(new_n1235), .A4(new_n1239), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(KEYINPUT125), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT125), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1241), .A2(new_n1245), .A3(new_n1242), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1227), .A2(new_n1230), .A3(new_n1244), .A4(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(KEYINPUT62), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1227), .A2(new_n1230), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1229), .A2(G2897), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1244), .A2(new_n1246), .A3(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1250), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1249), .A2(new_n1251), .A3(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT61), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1241), .A2(new_n1245), .A3(new_n1242), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1245), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1229), .B1(new_n1223), .B2(new_n1226), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT62), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1258), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1248), .A2(new_n1254), .A3(new_n1255), .A4(new_n1261), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n1066), .A2(new_n1068), .B1(new_n974), .B2(new_n999), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(G396), .A2(G393), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1217), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1264), .A2(KEYINPUT126), .A3(new_n1215), .A4(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT126), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1265), .A2(new_n1268), .A3(new_n1217), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1266), .A2(KEYINPUT126), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1269), .B(new_n1270), .C1(new_n1216), .C2(new_n1263), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1267), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1262), .A2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1252), .B1(new_n1258), .B2(new_n1250), .ZN(new_n1274));
  AOI21_X1  g1074(.A(KEYINPUT61), .B1(new_n1274), .B2(new_n1249), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1258), .A2(new_n1259), .A3(KEYINPUT63), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1272), .ZN(new_n1277));
  AND2_X1   g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT63), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1247), .A2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1275), .A2(new_n1278), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1273), .A2(new_n1281), .ZN(G405));
  NAND2_X1  g1082(.A1(G375), .A2(G378), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1220), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1284), .A2(KEYINPUT127), .A3(new_n1243), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1258), .A2(new_n1220), .A3(new_n1283), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT127), .B1(new_n1284), .B2(new_n1243), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1272), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1288), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1290), .A2(new_n1277), .A3(new_n1285), .A4(new_n1286), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1289), .A2(new_n1291), .ZN(G402));
endmodule


