//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 1 0 1 1 0 1 1 1 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 0 1 0 0 1 0 1 1 0 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n543,
    new_n544, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n567, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n612, new_n614, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT64), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT65), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT66), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT68), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n463), .A2(KEYINPUT3), .A3(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n465), .A2(G137), .A3(new_n466), .A4(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n463), .A2(new_n464), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n470), .A2(G101), .A3(new_n466), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  AND3_X1   g047(.A1(KEYINPUT67), .A2(G113), .A3(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(KEYINPUT67), .B1(G113), .B2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n468), .A2(new_n476), .A3(G125), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n466), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n472), .A2(new_n478), .ZN(G160));
  NAND2_X1  g054(.A1(new_n465), .A2(new_n468), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n480), .A2(new_n466), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n465), .A2(new_n468), .A3(new_n490), .ZN(new_n491));
  AND2_X1   g066(.A1(new_n468), .A2(new_n476), .ZN(new_n492));
  NOR3_X1   g067(.A1(new_n489), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n493));
  AOI22_X1  g068(.A1(new_n491), .A2(KEYINPUT4), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n465), .A2(G126), .A3(G2105), .A4(new_n468), .ZN(new_n495));
  OR2_X1    g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G114), .C2(new_n466), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n494), .A2(new_n498), .ZN(G164));
  XNOR2_X1  g074(.A(KEYINPUT6), .B(G651), .ZN(new_n500));
  AND2_X1   g075(.A1(new_n500), .A2(G543), .ZN(new_n501));
  AND3_X1   g076(.A1(KEYINPUT69), .A2(KEYINPUT5), .A3(G543), .ZN(new_n502));
  AOI21_X1  g077(.A(KEYINPUT5), .B1(KEYINPUT69), .B2(G543), .ZN(new_n503));
  AND2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  OAI22_X1  g080(.A1(new_n502), .A2(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(G50), .A2(new_n501), .B1(new_n507), .B2(G88), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT69), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(KEYINPUT69), .A2(KEYINPUT5), .A3(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G62), .ZN(new_n515));
  NAND2_X1  g090(.A1(G75), .A2(G543), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n509), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n508), .B1(KEYINPUT70), .B2(new_n517), .ZN(new_n518));
  AND2_X1   g093(.A1(new_n517), .A2(KEYINPUT70), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(G166));
  NAND3_X1  g095(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  INV_X1    g098(.A(G51), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n500), .A2(G543), .ZN(new_n525));
  OAI211_X1 g100(.A(new_n521), .B(new_n523), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n507), .A2(G89), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(G168));
  AOI22_X1  g103(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(new_n509), .ZN(new_n530));
  INV_X1    g105(.A(G52), .ZN(new_n531));
  INV_X1    g106(.A(G90), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n525), .A2(new_n531), .B1(new_n506), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n530), .A2(new_n533), .ZN(G171));
  INV_X1    g109(.A(G43), .ZN(new_n535));
  INV_X1    g110(.A(G81), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n525), .A2(new_n535), .B1(new_n506), .B2(new_n536), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT71), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(new_n509), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n538), .A2(G860), .A3(new_n540), .ZN(G153));
  NAND4_X1  g116(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g117(.A1(G1), .A2(G3), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT8), .ZN(new_n544));
  NAND4_X1  g119(.A1(G319), .A2(G483), .A3(G661), .A4(new_n544), .ZN(G188));
  NAND2_X1  g120(.A1(new_n506), .A2(KEYINPUT72), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT72), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n514), .A2(new_n547), .A3(new_n500), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n546), .A2(G91), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(KEYINPUT73), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT73), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n546), .A2(new_n548), .A3(new_n551), .A4(G91), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(G53), .ZN(new_n554));
  OAI21_X1  g129(.A(KEYINPUT9), .B1(new_n525), .B2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT9), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n501), .A2(new_n556), .A3(G53), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n514), .A2(G65), .ZN(new_n558));
  INV_X1    g133(.A(G78), .ZN(new_n559));
  INV_X1    g134(.A(G543), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n555), .A2(new_n557), .B1(new_n561), .B2(G651), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n553), .A2(new_n562), .ZN(G299));
  XNOR2_X1  g138(.A(G171), .B(KEYINPUT74), .ZN(G301));
  INV_X1    g139(.A(G168), .ZN(G286));
  INV_X1    g140(.A(G166), .ZN(G303));
  AND2_X1   g141(.A1(new_n546), .A2(new_n548), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G87), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n514), .A2(G74), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n569), .A2(G651), .B1(new_n501), .B2(G49), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(G288));
  NAND3_X1  g146(.A1(new_n546), .A2(G86), .A3(new_n548), .ZN(new_n572));
  OAI211_X1 g147(.A(G48), .B(G543), .C1(new_n504), .C2(new_n505), .ZN(new_n573));
  AND2_X1   g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g149(.A(G61), .B1(new_n502), .B2(new_n503), .ZN(new_n575));
  AND3_X1   g150(.A1(KEYINPUT75), .A2(G73), .A3(G543), .ZN(new_n576));
  AOI21_X1  g151(.A(KEYINPUT75), .B1(G73), .B2(G543), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g154(.A(KEYINPUT76), .B1(new_n579), .B2(G651), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT76), .ZN(new_n581));
  AOI211_X1 g156(.A(new_n581), .B(new_n509), .C1(new_n575), .C2(new_n578), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n574), .A2(new_n583), .ZN(G305));
  AOI22_X1  g159(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n509), .ZN(new_n586));
  INV_X1    g161(.A(G47), .ZN(new_n587));
  INV_X1    g162(.A(G85), .ZN(new_n588));
  OAI22_X1  g163(.A1(new_n525), .A2(new_n587), .B1(new_n506), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(KEYINPUT77), .ZN(new_n593));
  AND2_X1   g168(.A1(new_n592), .A2(KEYINPUT77), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n514), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G54), .ZN(new_n596));
  OAI22_X1  g171(.A1(new_n595), .A2(new_n509), .B1(new_n596), .B2(new_n525), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n567), .A2(G92), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT10), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n567), .A2(KEYINPUT10), .A3(G92), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n597), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n593), .B1(new_n594), .B2(new_n605), .ZN(G284));
  AOI21_X1  g181(.A(new_n593), .B1(new_n594), .B2(new_n605), .ZN(G321));
  NAND2_X1  g182(.A1(G286), .A2(G868), .ZN(new_n608));
  AND2_X1   g183(.A1(new_n553), .A2(new_n562), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(G868), .ZN(G297));
  OAI21_X1  g185(.A(new_n608), .B1(new_n609), .B2(G868), .ZN(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n602), .B1(new_n612), .B2(G860), .ZN(G148));
  NAND2_X1  g188(.A1(new_n538), .A2(new_n540), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(new_n604), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n603), .A2(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(new_n604), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g193(.A1(new_n492), .A2(new_n466), .A3(new_n470), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT78), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT13), .B(G2100), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n481), .A2(G135), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n483), .A2(G123), .ZN(new_n625));
  OR2_X1    g200(.A1(G99), .A2(G2105), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n626), .B(G2104), .C1(G111), .C2(new_n466), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n624), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n628), .A2(G2096), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(G2096), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n623), .A2(new_n629), .A3(new_n630), .ZN(G156));
  XNOR2_X1  g206(.A(G2427), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2430), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(KEYINPUT14), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT80), .ZN(new_n638));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2451), .B(G2454), .Z(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n640), .B(new_n643), .Z(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(G14), .A3(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(G401));
  INV_X1    g224(.A(KEYINPUT18), .ZN(new_n650));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(KEYINPUT17), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n651), .A2(new_n652), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n650), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2100), .ZN(new_n657));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  AOI21_X1  g233(.A(new_n658), .B1(new_n653), .B2(KEYINPUT18), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2096), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n657), .B(new_n660), .ZN(G227));
  XNOR2_X1  g236(.A(G1971), .B(G1976), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT19), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G1961), .B(G1966), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT81), .ZN(new_n666));
  XOR2_X1   g241(.A(G1956), .B(G2474), .Z(new_n667));
  NAND3_X1  g242(.A1(new_n664), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT20), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n664), .B1(new_n666), .B2(new_n667), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n666), .A2(new_n667), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OAI211_X1 g247(.A(new_n669), .B(new_n672), .C1(new_n663), .C2(new_n671), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1991), .B(G1996), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1981), .B(G1986), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n677), .B(new_n678), .Z(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(G229));
  INV_X1    g255(.A(G16), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(G23), .ZN(new_n682));
  INV_X1    g257(.A(G288), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n682), .B1(new_n683), .B2(new_n681), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT33), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G1976), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n681), .A2(G22), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(G166), .B2(new_n681), .ZN(new_n688));
  INV_X1    g263(.A(G1971), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  MUX2_X1   g265(.A(G6), .B(G305), .S(G16), .Z(new_n691));
  XOR2_X1   g266(.A(KEYINPUT32), .B(G1981), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n686), .A2(new_n690), .A3(new_n693), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n694), .A2(KEYINPUT34), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(KEYINPUT34), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT82), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(KEYINPUT36), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n590), .A2(G16), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G16), .B2(G24), .ZN(new_n700));
  INV_X1    g275(.A(G1986), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n698), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n481), .A2(G131), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n483), .A2(G119), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n466), .A2(G107), .ZN(new_n705));
  OAI21_X1  g280(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n703), .B(new_n704), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  MUX2_X1   g282(.A(G25), .B(new_n707), .S(G29), .Z(new_n708));
  XOR2_X1   g283(.A(KEYINPUT35), .B(G1991), .Z(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n708), .B(new_n710), .ZN(new_n711));
  AOI211_X1 g286(.A(new_n702), .B(new_n711), .C1(new_n701), .C2(new_n700), .ZN(new_n712));
  AND3_X1   g287(.A1(new_n695), .A2(new_n696), .A3(new_n712), .ZN(new_n713));
  OR3_X1    g288(.A1(new_n713), .A2(new_n697), .A3(KEYINPUT36), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n697), .B2(KEYINPUT36), .ZN(new_n715));
  INV_X1    g290(.A(G29), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G33), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n481), .A2(G139), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT85), .B(KEYINPUT25), .Z(new_n719));
  NAND3_X1  g294(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n492), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n718), .B(new_n721), .C1(new_n466), .C2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n717), .B1(new_n724), .B2(new_n716), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT86), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G2072), .ZN(new_n727));
  INV_X1    g302(.A(G1348), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n602), .A2(new_n681), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G4), .B2(new_n681), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n727), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT31), .B(G11), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT90), .Z(new_n733));
  INV_X1    g308(.A(KEYINPUT30), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n716), .B1(new_n734), .B2(G28), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n735), .A2(KEYINPUT91), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n734), .A2(G28), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n735), .B2(KEYINPUT91), .ZN(new_n738));
  OAI221_X1 g313(.A(new_n733), .B1(new_n736), .B2(new_n738), .C1(new_n628), .C2(new_n716), .ZN(new_n739));
  NOR2_X1   g314(.A1(G171), .A2(new_n681), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G5), .B2(new_n681), .ZN(new_n741));
  INV_X1    g316(.A(G1961), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n739), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n742), .B2(new_n741), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n481), .A2(G140), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n483), .A2(G128), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n466), .A2(G116), .ZN(new_n747));
  OAI21_X1  g322(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n745), .B(new_n746), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G29), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT83), .B(KEYINPUT28), .Z(new_n751));
  NAND2_X1  g326(.A1(new_n716), .A2(G26), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT84), .B(G2067), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n754), .A2(new_n755), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT24), .ZN(new_n758));
  INV_X1    g333(.A(G34), .ZN(new_n759));
  AOI21_X1  g334(.A(G29), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n758), .B2(new_n759), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G160), .B2(new_n716), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(G2084), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n762), .A2(G2084), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n756), .A2(new_n757), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G1341), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n681), .A2(G19), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n614), .B2(G16), .ZN(new_n768));
  AOI211_X1 g343(.A(new_n744), .B(new_n765), .C1(new_n766), .C2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n681), .A2(G20), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT23), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n609), .B2(new_n681), .ZN(new_n772));
  INV_X1    g347(.A(G1956), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n481), .A2(G141), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT87), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n483), .A2(G129), .ZN(new_n777));
  NAND3_X1  g352(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT26), .Z(new_n779));
  NAND3_X1  g354(.A1(new_n470), .A2(G105), .A3(new_n466), .ZN(new_n780));
  AND4_X1   g355(.A1(new_n776), .A2(new_n777), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n781), .A2(new_n716), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n716), .B2(G32), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT27), .B(G1996), .ZN(new_n784));
  OAI22_X1  g359(.A1(new_n783), .A2(new_n784), .B1(new_n766), .B2(new_n768), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n681), .A2(G21), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G168), .B2(new_n681), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT89), .ZN(new_n788));
  INV_X1    g363(.A(G1966), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n785), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n731), .A2(new_n769), .A3(new_n774), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n716), .A2(G35), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G162), .B2(new_n716), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT29), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n795), .A2(G2090), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT94), .Z(new_n797));
  INV_X1    g372(.A(new_n730), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n716), .A2(G27), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G164), .B2(new_n716), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT92), .Z(new_n801));
  AOI22_X1  g376(.A1(new_n798), .A2(G1348), .B1(G2078), .B2(new_n801), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n797), .B(new_n802), .C1(G2078), .C2(new_n801), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n783), .A2(new_n784), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT88), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n795), .A2(G2090), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT93), .Z(new_n807));
  NOR4_X1   g382(.A1(new_n792), .A2(new_n803), .A3(new_n805), .A4(new_n807), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n714), .A2(new_n715), .A3(new_n808), .ZN(G150));
  INV_X1    g384(.A(G150), .ZN(G311));
  INV_X1    g385(.A(G55), .ZN(new_n811));
  INV_X1    g386(.A(G93), .ZN(new_n812));
  OAI22_X1  g387(.A1(new_n525), .A2(new_n811), .B1(new_n506), .B2(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT95), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n814), .B1(new_n509), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(G860), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT37), .Z(new_n818));
  NAND2_X1  g393(.A1(new_n602), .A2(G559), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT38), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n816), .A2(new_n614), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n816), .A2(new_n614), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n820), .B(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(KEYINPUT39), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT96), .Z(new_n827));
  INV_X1    g402(.A(G860), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n825), .B2(KEYINPUT39), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n818), .B1(new_n827), .B2(new_n829), .ZN(G145));
  NAND2_X1  g405(.A1(new_n483), .A2(G130), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n466), .A2(G118), .ZN(new_n832));
  OAI21_X1  g407(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(G142), .B2(new_n481), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(new_n707), .Z(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(new_n621), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n749), .B(G164), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n781), .B(new_n838), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n839), .A2(new_n724), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT98), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n839), .A2(new_n724), .ZN(new_n842));
  AND3_X1   g417(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n841), .B1(new_n840), .B2(new_n842), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n837), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(KEYINPUT99), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT99), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n847), .B(new_n837), .C1(new_n843), .C2(new_n844), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(G160), .B(KEYINPUT97), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n487), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n628), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n840), .A2(new_n842), .ZN(new_n854));
  INV_X1    g429(.A(new_n837), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n849), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n854), .B(new_n855), .ZN(new_n858));
  AOI21_X1  g433(.A(G37), .B1(new_n858), .B2(new_n853), .ZN(new_n859));
  AND3_X1   g434(.A1(new_n857), .A2(KEYINPUT40), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(KEYINPUT40), .B1(new_n857), .B2(new_n859), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n860), .A2(new_n861), .ZN(G395));
  NAND2_X1  g437(.A1(new_n816), .A2(new_n604), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n609), .A2(KEYINPUT100), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT100), .ZN(new_n865));
  NAND2_X1  g440(.A1(G299), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n602), .A3(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n603), .A2(new_n865), .A3(G299), .ZN(new_n868));
  AND2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT41), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n867), .A2(new_n868), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(KEYINPUT41), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n823), .B(new_n616), .ZN(new_n875));
  MUX2_X1   g450(.A(new_n869), .B(new_n874), .S(new_n875), .Z(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT42), .ZN(new_n877));
  XOR2_X1   g452(.A(G166), .B(G305), .Z(new_n878));
  XNOR2_X1  g453(.A(G288), .B(new_n590), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n877), .B(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n863), .B1(new_n882), .B2(new_n604), .ZN(G295));
  OAI21_X1  g458(.A(new_n863), .B1(new_n882), .B2(new_n604), .ZN(G331));
  INV_X1    g459(.A(KEYINPUT44), .ZN(new_n885));
  NOR2_X1   g460(.A1(G301), .A2(G286), .ZN(new_n886));
  NOR2_X1   g461(.A1(G168), .A2(G171), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(new_n823), .ZN(new_n889));
  OAI211_X1 g464(.A(new_n821), .B(new_n822), .C1(new_n886), .C2(new_n887), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n874), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n889), .A2(new_n890), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(new_n869), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n892), .A2(new_n881), .A3(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(G37), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n893), .B1(new_n871), .B2(new_n873), .ZN(new_n898));
  INV_X1    g473(.A(new_n894), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n880), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  XOR2_X1   g475(.A(KEYINPUT101), .B(KEYINPUT43), .Z(new_n901));
  NAND3_X1  g476(.A1(new_n897), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n871), .A2(KEYINPUT102), .A3(new_n873), .ZN(new_n903));
  OAI211_X1 g478(.A(new_n903), .B(new_n891), .C1(KEYINPUT102), .C2(new_n873), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n881), .B1(new_n904), .B2(new_n894), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n895), .A2(new_n896), .ZN(new_n906));
  OAI21_X1  g481(.A(KEYINPUT43), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n885), .B1(new_n902), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT103), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT102), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n874), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n891), .B1(new_n873), .B2(KEYINPUT102), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n894), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(new_n880), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n897), .A2(new_n914), .A3(new_n901), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n900), .A2(new_n895), .A3(new_n896), .ZN(new_n916));
  INV_X1    g491(.A(new_n901), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n909), .B1(new_n915), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n905), .A2(new_n906), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT103), .B1(new_n920), .B2(new_n901), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n908), .B1(new_n922), .B2(new_n885), .ZN(G397));
  AND3_X1   g498(.A1(new_n468), .A2(new_n476), .A3(G125), .ZN(new_n924));
  NAND2_X1  g499(.A1(G113), .A2(G2104), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT67), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(KEYINPUT67), .A2(G113), .A3(G2104), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(G2105), .B1(new_n924), .B2(new_n929), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n930), .A2(G40), .A3(new_n471), .A4(new_n469), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT104), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n469), .A2(new_n471), .ZN(new_n934));
  INV_X1    g509(.A(G40), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n478), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n934), .A2(new_n936), .A3(KEYINPUT104), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n933), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(G1384), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(new_n494), .B2(new_n498), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(KEYINPUT50), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT50), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n942), .B(new_n939), .C1(new_n494), .C2(new_n498), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n938), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n773), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT45), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n940), .A2(new_n946), .ZN(new_n947));
  OAI211_X1 g522(.A(KEYINPUT45), .B(new_n939), .C1(new_n494), .C2(new_n498), .ZN(new_n948));
  XNOR2_X1  g523(.A(KEYINPUT56), .B(G2072), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n938), .A2(new_n947), .A3(new_n948), .A4(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n945), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n557), .A2(new_n555), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT115), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT57), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n955), .A2(new_n553), .A3(new_n562), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT57), .B1(new_n952), .B2(KEYINPUT115), .ZN(new_n957));
  NAND2_X1  g532(.A1(G299), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n951), .A2(new_n960), .A3(KEYINPUT117), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT117), .B1(new_n951), .B2(new_n960), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(G2067), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n940), .B1(new_n933), .B2(new_n937), .ZN(new_n966));
  AOI22_X1  g541(.A1(new_n944), .A2(new_n728), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n964), .B1(new_n603), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT116), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n938), .A2(new_n947), .A3(new_n948), .ZN(new_n970));
  AOI22_X1  g545(.A1(new_n970), .A2(new_n949), .B1(new_n944), .B2(new_n773), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n969), .B1(new_n971), .B2(new_n959), .ZN(new_n972));
  AND4_X1   g547(.A1(new_n969), .A2(new_n959), .A3(new_n945), .A4(new_n950), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n968), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n951), .A2(new_n960), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n975), .B1(new_n972), .B2(new_n973), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT61), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n614), .A2(KEYINPUT120), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n492), .A2(new_n493), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n498), .ZN(new_n983));
  AOI21_X1  g558(.A(G1384), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n931), .A2(new_n932), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT104), .B1(new_n934), .B2(new_n936), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n984), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n988), .B(G1341), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT119), .ZN(new_n991));
  INV_X1    g566(.A(G1996), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n938), .A2(new_n947), .A3(new_n992), .A4(new_n948), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n990), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n991), .B1(new_n990), .B2(new_n993), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n979), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT59), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT59), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n998), .B(new_n979), .C1(new_n994), .C2(new_n995), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n963), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n977), .B1(new_n971), .B2(new_n959), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1001), .A2(new_n961), .A3(new_n1002), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n978), .A2(new_n1000), .A3(KEYINPUT121), .A4(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n967), .B(new_n603), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n603), .A2(KEYINPUT60), .ZN(new_n1006));
  AOI22_X1  g581(.A1(new_n1005), .A2(KEYINPUT60), .B1(new_n967), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  AOI22_X1  g583(.A1(new_n964), .A2(new_n1002), .B1(new_n997), .B2(new_n999), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT121), .B1(new_n1009), .B2(new_n978), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n974), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n944), .A2(new_n742), .ZN(new_n1012));
  INV_X1    g587(.A(G2078), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n970), .A2(KEYINPUT53), .A3(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n938), .A2(new_n947), .A3(new_n948), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(KEYINPUT108), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT108), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n938), .A2(new_n947), .A3(new_n1017), .A4(new_n948), .ZN(new_n1018));
  AOI21_X1  g593(.A(G2078), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1012), .B(new_n1014), .C1(new_n1019), .C2(KEYINPUT53), .ZN(new_n1020));
  INV_X1    g595(.A(G301), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT54), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT123), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1023), .B1(new_n944), .B2(new_n742), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1012), .A2(KEYINPUT123), .ZN(new_n1025));
  INV_X1    g600(.A(new_n936), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n934), .A2(KEYINPUT124), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT124), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n472), .A2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1026), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n1030), .A2(new_n947), .A3(KEYINPUT125), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT125), .B1(new_n1030), .B2(new_n947), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  OR2_X1    g608(.A1(new_n1013), .A2(KEYINPUT126), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1035), .B1(KEYINPUT126), .B2(new_n1013), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n948), .A2(new_n1034), .A3(new_n1036), .ZN(new_n1037));
  OAI22_X1  g612(.A1(new_n1024), .A2(new_n1025), .B1(new_n1033), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT53), .B1(new_n1039), .B2(new_n1013), .ZN(new_n1040));
  OAI21_X1  g615(.A(G171), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT127), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT127), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1043), .B(G171), .C1(new_n1038), .C2(new_n1040), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1022), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n1046));
  INV_X1    g621(.A(G8), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n966), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n683), .A2(G1976), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1046), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1051));
  INV_X1    g626(.A(G1976), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT52), .B1(G288), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1050), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G61), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1055), .B1(new_n512), .B2(new_n513), .ZN(new_n1056));
  INV_X1    g631(.A(new_n577), .ZN(new_n1057));
  NAND3_X1  g632(.A1(KEYINPUT75), .A2(G73), .A3(G543), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(G651), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(new_n581), .ZN(new_n1061));
  INV_X1    g636(.A(G86), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n573), .B1(new_n506), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT111), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n579), .A2(KEYINPUT76), .A3(G651), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT111), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1066), .B(new_n573), .C1(new_n506), .C2(new_n1062), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1061), .A2(new_n1064), .A3(new_n1065), .A4(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(G1981), .ZN(new_n1069));
  XNOR2_X1  g644(.A(KEYINPUT110), .B(G1981), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n574), .A2(new_n583), .A3(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1069), .A2(new_n1071), .A3(KEYINPUT49), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT112), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1069), .A2(new_n1071), .A3(KEYINPUT112), .A4(KEYINPUT49), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n987), .A2(G8), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT49), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AND3_X1   g654(.A1(new_n1076), .A2(KEYINPUT113), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT113), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1054), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1016), .A2(new_n689), .A3(new_n1018), .ZN(new_n1083));
  OR2_X1    g658(.A1(new_n944), .A2(G2090), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(G8), .B1(new_n518), .B2(new_n519), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n1087));
  XNOR2_X1  g662(.A(new_n1086), .B(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1085), .A2(G8), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1082), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1085), .A2(G8), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1088), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n938), .A2(new_n941), .A3(new_n943), .ZN(new_n1095));
  INV_X1    g670(.A(G2084), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1095), .A2(new_n1096), .B1(new_n1015), .B2(new_n789), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1047), .B1(new_n1097), .B2(G168), .ZN(new_n1098));
  XOR2_X1   g673(.A(KEYINPUT122), .B(KEYINPUT51), .Z(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  OR3_X1    g675(.A1(new_n1097), .A2(new_n1047), .A3(G168), .ZN(new_n1101));
  NAND2_X1  g676(.A1(KEYINPUT122), .A2(KEYINPUT51), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1100), .B(new_n1101), .C1(new_n1098), .C2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1091), .A2(new_n1094), .A3(new_n1103), .ZN(new_n1104));
  OR3_X1    g679(.A1(new_n1038), .A2(new_n1040), .A3(new_n1021), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT54), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n1045), .A2(new_n1104), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1011), .A2(new_n1108), .ZN(new_n1109));
  XOR2_X1   g684(.A(new_n1103), .B(KEYINPUT62), .Z(new_n1110));
  INV_X1    g685(.A(new_n1106), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1110), .A2(new_n1094), .A3(new_n1091), .A4(new_n1111), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n1097), .A2(new_n1047), .A3(G286), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1091), .A2(KEYINPUT63), .A3(new_n1094), .A4(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1048), .A2(new_n1049), .A3(new_n1053), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(new_n1051), .B2(new_n1046), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1076), .A2(new_n1079), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT113), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1076), .A2(KEYINPUT113), .A3(new_n1079), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1116), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1121), .A2(new_n1094), .A3(new_n1089), .A4(new_n1113), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT63), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1114), .A2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n683), .A2(new_n1052), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1071), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n1128), .A2(new_n1048), .B1(new_n1121), .B2(new_n1090), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1125), .A2(KEYINPUT114), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(KEYINPUT114), .B1(new_n1125), .B2(new_n1129), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1109), .B(new_n1112), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n947), .B1(new_n937), .B2(new_n933), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n1134), .A2(new_n781), .A3(new_n992), .ZN(new_n1135));
  XOR2_X1   g710(.A(new_n1135), .B(KEYINPUT105), .Z(new_n1136));
  NOR2_X1   g711(.A1(new_n1134), .A2(G1996), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1136), .B1(new_n781), .B2(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n749), .B(G2067), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(KEYINPUT106), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1140), .A2(new_n1134), .ZN(new_n1141));
  XOR2_X1   g716(.A(new_n1141), .B(KEYINPUT107), .Z(new_n1142));
  AND2_X1   g717(.A1(new_n1138), .A2(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n707), .B(new_n709), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1143), .B1(new_n1134), .B2(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n590), .B(new_n701), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1145), .B1(new_n1133), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1132), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1134), .B1(new_n1140), .B2(new_n781), .ZN(new_n1149));
  OAI21_X1  g724(.A(KEYINPUT46), .B1(new_n1134), .B2(G1996), .ZN(new_n1150));
  OR3_X1    g725(.A1(new_n1134), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1149), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  XOR2_X1   g727(.A(new_n1152), .B(KEYINPUT47), .Z(new_n1153));
  NAND3_X1  g728(.A1(new_n1133), .A2(new_n701), .A3(new_n590), .ZN(new_n1154));
  XOR2_X1   g729(.A(new_n1154), .B(KEYINPUT48), .Z(new_n1155));
  OAI21_X1  g730(.A(new_n1153), .B1(new_n1145), .B2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n707), .A2(new_n710), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1143), .A2(new_n1157), .ZN(new_n1158));
  OR2_X1    g733(.A1(new_n749), .A2(G2067), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1134), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1156), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1148), .A2(new_n1161), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g737(.A1(G227), .A2(new_n459), .ZN(new_n1164));
  AND3_X1   g738(.A1(new_n679), .A2(new_n648), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g739(.A(new_n856), .ZN(new_n1166));
  AOI21_X1  g740(.A(new_n1166), .B1(new_n846), .B2(new_n848), .ZN(new_n1167));
  INV_X1    g741(.A(new_n859), .ZN(new_n1168));
  OAI21_X1  g742(.A(new_n1165), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g743(.A1(new_n922), .A2(new_n1169), .ZN(G308));
  OAI221_X1 g744(.A(new_n1165), .B1(new_n1167), .B2(new_n1168), .C1(new_n919), .C2(new_n921), .ZN(G225));
endmodule


