

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744;

  NOR2_X1 U362 ( .A1(n707), .A2(n716), .ZN(n708) );
  AND2_X1 U363 ( .A1(n620), .A2(n420), .ZN(n416) );
  XNOR2_X1 U364 ( .A(n514), .B(n513), .ZN(n741) );
  NAND2_X1 U365 ( .A1(n527), .A2(n584), .ZN(n463) );
  AND2_X1 U366 ( .A1(n399), .A2(n398), .ZN(n397) );
  XNOR2_X1 U367 ( .A(n572), .B(n448), .ZN(n519) );
  OR2_X1 U368 ( .A1(n611), .A2(G902), .ZN(n447) );
  XNOR2_X1 U369 ( .A(n414), .B(n724), .ZN(n704) );
  XNOR2_X1 U370 ( .A(n506), .B(n426), .ZN(n444) );
  XNOR2_X1 U371 ( .A(n679), .B(G128), .ZN(n466) );
  XNOR2_X1 U372 ( .A(n468), .B(KEYINPUT77), .ZN(n470) );
  NAND2_X1 U373 ( .A1(n717), .A2(G224), .ZN(n468) );
  INV_X2 U374 ( .A(G143), .ZN(n679) );
  NOR2_X2 U375 ( .A1(n662), .A2(n423), .ZN(n422) );
  XNOR2_X2 U376 ( .A(n524), .B(n523), .ZN(n662) );
  INV_X4 U377 ( .A(G953), .ZN(n717) );
  XNOR2_X1 U378 ( .A(KEYINPUT86), .B(KEYINPUT15), .ZN(n449) );
  BUF_X1 U379 ( .A(n569), .Z(n340) );
  NOR2_X1 U380 ( .A1(n563), .A2(n562), .ZN(n581) );
  XNOR2_X1 U381 ( .A(n435), .B(G472), .ZN(n569) );
  XNOR2_X2 U382 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n465) );
  XNOR2_X2 U383 ( .A(KEYINPUT18), .B(KEYINPUT78), .ZN(n464) );
  XNOR2_X2 U384 ( .A(n602), .B(n342), .ZN(n639) );
  NAND2_X1 U385 ( .A1(n386), .A2(n384), .ZN(n655) );
  AND2_X1 U386 ( .A1(n371), .A2(n370), .ZN(n369) );
  OR2_X1 U387 ( .A1(n661), .A2(n660), .ZN(n405) );
  XNOR2_X1 U388 ( .A(n545), .B(KEYINPUT108), .ZN(n546) );
  NAND2_X2 U389 ( .A1(n369), .A2(n365), .ZN(n602) );
  XNOR2_X2 U390 ( .A(n463), .B(KEYINPUT33), .ZN(n648) );
  NOR2_X1 U391 ( .A1(G953), .A2(G237), .ZN(n494) );
  XNOR2_X1 U392 ( .A(n466), .B(n425), .ZN(n506) );
  INV_X1 U393 ( .A(G134), .ZN(n425) );
  XNOR2_X1 U394 ( .A(G146), .B(G125), .ZN(n469) );
  XNOR2_X1 U395 ( .A(n349), .B(n344), .ZN(n538) );
  OR2_X1 U396 ( .A1(n671), .A2(G902), .ZN(n349) );
  XNOR2_X1 U397 ( .A(n469), .B(n393), .ZN(n731) );
  INV_X1 U398 ( .A(KEYINPUT10), .ZN(n393) );
  NOR2_X1 U399 ( .A1(n600), .A2(n599), .ZN(n601) );
  NAND2_X1 U400 ( .A1(n602), .A2(n638), .ZN(n586) );
  XNOR2_X1 U401 ( .A(n511), .B(n510), .ZN(n539) );
  XNOR2_X1 U402 ( .A(n352), .B(n351), .ZN(n363) );
  INV_X1 U403 ( .A(KEYINPUT107), .ZN(n351) );
  NAND2_X1 U404 ( .A1(n687), .A2(n691), .ZN(n352) );
  NOR2_X1 U405 ( .A1(n360), .A2(n699), .ZN(n592) );
  NAND2_X1 U406 ( .A1(n377), .A2(n519), .ZN(n376) );
  XNOR2_X1 U407 ( .A(n354), .B(n459), .ZN(n460) );
  XNOR2_X1 U408 ( .A(n358), .B(n434), .ZN(n665) );
  XNOR2_X1 U409 ( .A(n444), .B(n343), .ZN(n358) );
  BUF_X1 U410 ( .A(n619), .Z(n733) );
  XNOR2_X1 U411 ( .A(G110), .B(KEYINPUT90), .ZN(n453) );
  XNOR2_X1 U412 ( .A(n452), .B(n391), .ZN(n390) );
  XNOR2_X1 U413 ( .A(G128), .B(G119), .ZN(n391) );
  XNOR2_X1 U414 ( .A(G107), .B(KEYINPUT7), .ZN(n502) );
  XOR2_X1 U415 ( .A(KEYINPUT104), .B(KEYINPUT103), .Z(n503) );
  XNOR2_X1 U416 ( .A(n506), .B(n341), .ZN(n374) );
  XNOR2_X1 U417 ( .A(n350), .B(n500), .ZN(n671) );
  XNOR2_X1 U418 ( .A(n499), .B(n731), .ZN(n350) );
  XNOR2_X1 U419 ( .A(G122), .B(G113), .ZN(n492) );
  XNOR2_X1 U420 ( .A(n473), .B(n375), .ZN(n445) );
  XNOR2_X1 U421 ( .A(n442), .B(n439), .ZN(n375) );
  XOR2_X1 U422 ( .A(G146), .B(G101), .Z(n439) );
  INV_X1 U423 ( .A(KEYINPUT110), .ZN(n348) );
  NAND2_X1 U424 ( .A1(n383), .A2(n385), .ZN(n384) );
  AND2_X1 U425 ( .A1(n388), .A2(n387), .ZN(n386) );
  NOR2_X1 U426 ( .A1(n641), .A2(n345), .ZN(n385) );
  XNOR2_X1 U427 ( .A(n357), .B(KEYINPUT109), .ZN(n356) );
  NAND2_X1 U428 ( .A1(n368), .A2(n367), .ZN(n366) );
  XNOR2_X1 U429 ( .A(n538), .B(n410), .ZN(n540) );
  INV_X1 U430 ( .A(KEYINPUT102), .ZN(n410) );
  BUF_X1 U431 ( .A(n518), .Z(n629) );
  NAND2_X1 U432 ( .A1(n528), .A2(n516), .ZN(n400) );
  NOR2_X1 U433 ( .A1(n641), .A2(n515), .ZN(n516) );
  BUF_X1 U434 ( .A(n701), .Z(n712) );
  AND2_X1 U435 ( .A1(n616), .A2(G953), .ZN(n716) );
  NOR2_X1 U436 ( .A1(n624), .A2(n623), .ZN(n661) );
  XNOR2_X1 U437 ( .A(n362), .B(n590), .ZN(n361) );
  INV_X1 U438 ( .A(n682), .ZN(n378) );
  INV_X1 U439 ( .A(n363), .ZN(n643) );
  XNOR2_X1 U440 ( .A(n355), .B(KEYINPUT20), .ZN(n458) );
  INV_X1 U441 ( .A(G237), .ZN(n477) );
  NAND2_X1 U442 ( .A1(n458), .A2(G217), .ZN(n354) );
  XNOR2_X1 U443 ( .A(G131), .B(KEYINPUT4), .ZN(n426) );
  XNOR2_X1 U444 ( .A(G146), .B(G137), .ZN(n427) );
  XOR2_X1 U445 ( .A(KEYINPUT98), .B(KEYINPUT11), .Z(n497) );
  XNOR2_X1 U446 ( .A(G143), .B(G104), .ZN(n495) );
  XNOR2_X1 U447 ( .A(n407), .B(n406), .ZN(n493) );
  XNOR2_X1 U448 ( .A(KEYINPUT100), .B(KEYINPUT99), .ZN(n406) );
  XNOR2_X1 U449 ( .A(n408), .B(G140), .ZN(n407) );
  XNOR2_X1 U450 ( .A(G131), .B(KEYINPUT12), .ZN(n408) );
  XNOR2_X1 U451 ( .A(KEYINPUT3), .B(G119), .ZN(n431) );
  NAND2_X1 U452 ( .A1(n641), .A2(n345), .ZN(n387) );
  INV_X1 U453 ( .A(n476), .ZN(n368) );
  INV_X1 U454 ( .A(n479), .ZN(n367) );
  NAND2_X1 U455 ( .A1(n476), .A2(n479), .ZN(n370) );
  NOR2_X1 U456 ( .A1(n568), .A2(n630), .ZN(n585) );
  OR2_X2 U457 ( .A1(n518), .A2(n515), .ZN(n353) );
  INV_X1 U458 ( .A(G902), .ZN(n478) );
  NAND2_X1 U459 ( .A1(n396), .A2(n395), .ZN(n394) );
  NOR2_X1 U460 ( .A1(n489), .A2(n346), .ZN(n395) );
  XNOR2_X1 U461 ( .A(n438), .B(n437), .ZN(n723) );
  INV_X1 U462 ( .A(G104), .ZN(n437) );
  XNOR2_X1 U463 ( .A(n723), .B(KEYINPUT70), .ZN(n473) );
  NOR2_X1 U464 ( .A1(n621), .A2(KEYINPUT2), .ZN(n624) );
  XNOR2_X1 U465 ( .A(n565), .B(n564), .ZN(n412) );
  NAND2_X1 U466 ( .A1(n581), .A2(n639), .ZN(n565) );
  XNOR2_X1 U467 ( .A(n340), .B(n436), .ZN(n584) );
  XOR2_X1 U468 ( .A(n665), .B(n664), .Z(n666) );
  XNOR2_X1 U469 ( .A(n392), .B(n389), .ZN(n713) );
  XNOR2_X1 U470 ( .A(n455), .B(n390), .ZN(n389) );
  XNOR2_X1 U471 ( .A(n457), .B(n731), .ZN(n392) );
  XNOR2_X1 U472 ( .A(n505), .B(n374), .ZN(n509) );
  XNOR2_X1 U473 ( .A(KEYINPUT59), .B(n671), .ZN(n672) );
  AND2_X1 U474 ( .A1(n604), .A2(n603), .ZN(n663) );
  XNOR2_X1 U475 ( .A(n601), .B(n347), .ZN(n604) );
  XNOR2_X1 U476 ( .A(n348), .B(KEYINPUT43), .ZN(n347) );
  NAND2_X1 U477 ( .A1(n589), .A2(n655), .ZN(n576) );
  XNOR2_X1 U478 ( .A(n587), .B(KEYINPUT36), .ZN(n359) );
  XNOR2_X1 U479 ( .A(n541), .B(KEYINPUT106), .ZN(n687) );
  AND2_X1 U480 ( .A1(n525), .A2(n629), .ZN(n372) );
  XNOR2_X1 U481 ( .A(n615), .B(n614), .ZN(n618) );
  INV_X1 U482 ( .A(KEYINPUT53), .ZN(n401) );
  XNOR2_X1 U483 ( .A(n542), .B(G101), .ZN(G3) );
  XNOR2_X1 U484 ( .A(n449), .B(G902), .ZN(n607) );
  XOR2_X1 U485 ( .A(G116), .B(G122), .Z(n341) );
  XOR2_X1 U486 ( .A(KEYINPUT72), .B(KEYINPUT38), .Z(n342) );
  XOR2_X1 U487 ( .A(n428), .B(n427), .Z(n343) );
  XNOR2_X1 U488 ( .A(n586), .B(n481), .ZN(n588) );
  XOR2_X1 U489 ( .A(n501), .B(G475), .Z(n344) );
  BUF_X1 U490 ( .A(n519), .Z(n600) );
  XOR2_X1 U491 ( .A(KEYINPUT41), .B(KEYINPUT113), .Z(n345) );
  XNOR2_X1 U492 ( .A(n530), .B(n529), .ZN(n694) );
  XNOR2_X1 U493 ( .A(KEYINPUT67), .B(KEYINPUT0), .ZN(n346) );
  INV_X1 U494 ( .A(KEYINPUT46), .ZN(n380) );
  INV_X1 U495 ( .A(KEYINPUT2), .ZN(n420) );
  XNOR2_X2 U496 ( .A(n608), .B(KEYINPUT80), .ZN(n619) );
  NAND2_X1 U497 ( .A1(n605), .A2(n606), .ZN(n608) );
  NAND2_X1 U498 ( .A1(n356), .A2(n695), .ZN(n597) );
  NOR2_X1 U499 ( .A1(n413), .A2(n572), .ZN(n531) );
  XNOR2_X2 U500 ( .A(n353), .B(KEYINPUT68), .ZN(n413) );
  XNOR2_X1 U501 ( .A(n461), .B(n462), .ZN(n518) );
  NAND2_X1 U502 ( .A1(n607), .A2(G234), .ZN(n355) );
  NAND2_X1 U503 ( .A1(n585), .A2(n584), .ZN(n357) );
  AND2_X1 U504 ( .A1(n359), .A2(n600), .ZN(n699) );
  NAND2_X1 U505 ( .A1(n361), .A2(n591), .ZN(n360) );
  NAND2_X1 U506 ( .A1(n364), .A2(n363), .ZN(n362) );
  INV_X1 U507 ( .A(n692), .ZN(n364) );
  OR2_X1 U508 ( .A1(n704), .A2(n366), .ZN(n365) );
  NAND2_X1 U509 ( .A1(n704), .A2(n479), .ZN(n371) );
  NAND2_X1 U510 ( .A1(n535), .A2(n372), .ZN(n686) );
  NAND2_X1 U511 ( .A1(n535), .A2(n373), .ZN(n524) );
  AND2_X1 U512 ( .A1(n521), .A2(n629), .ZN(n373) );
  XNOR2_X1 U513 ( .A(n471), .B(n472), .ZN(n415) );
  NAND2_X1 U514 ( .A1(n550), .A2(KEYINPUT44), .ZN(n547) );
  NAND2_X1 U515 ( .A1(n526), .A2(n741), .ZN(n550) );
  XOR2_X1 U516 ( .A(n460), .B(KEYINPUT91), .Z(n461) );
  INV_X1 U517 ( .A(n382), .ZN(n742) );
  NAND2_X1 U518 ( .A1(n382), .A2(n379), .ZN(n577) );
  XNOR2_X2 U519 ( .A(n566), .B(KEYINPUT40), .ZN(n382) );
  INV_X1 U520 ( .A(n600), .ZN(n583) );
  XNOR2_X2 U521 ( .A(n376), .B(KEYINPUT73), .ZN(n527) );
  INV_X1 U522 ( .A(n413), .ZN(n377) );
  INV_X1 U523 ( .A(n340), .ZN(n627) );
  INV_X1 U524 ( .A(n584), .ZN(n520) );
  NAND2_X1 U525 ( .A1(n378), .A2(n542), .ZN(n537) );
  NAND2_X1 U526 ( .A1(n536), .A2(n535), .ZN(n542) );
  INV_X1 U527 ( .A(n744), .ZN(n379) );
  NAND2_X1 U528 ( .A1(n381), .A2(n382), .ZN(n578) );
  NOR2_X1 U529 ( .A1(n744), .A2(n380), .ZN(n381) );
  INV_X1 U530 ( .A(n644), .ZN(n383) );
  XNOR2_X2 U531 ( .A(n574), .B(KEYINPUT112), .ZN(n644) );
  NAND2_X1 U532 ( .A1(n644), .A2(n345), .ZN(n388) );
  NOR2_X1 U533 ( .A1(n668), .A2(n716), .ZN(n670) );
  NOR2_X1 U534 ( .A1(n417), .A2(n416), .ZN(n610) );
  NOR2_X1 U535 ( .A1(n674), .A2(n716), .ZN(n677) );
  NAND2_X1 U536 ( .A1(n418), .A2(n476), .ZN(n417) );
  NAND2_X2 U537 ( .A1(n397), .A2(n394), .ZN(n528) );
  INV_X1 U538 ( .A(n588), .ZN(n396) );
  NAND2_X1 U539 ( .A1(n489), .A2(n346), .ZN(n398) );
  NAND2_X1 U540 ( .A1(n588), .A2(n346), .ZN(n399) );
  XNOR2_X2 U541 ( .A(n400), .B(n517), .ZN(n535) );
  XNOR2_X1 U542 ( .A(n402), .B(n401), .ZN(G75) );
  NAND2_X1 U543 ( .A1(n403), .A2(n717), .ZN(n402) );
  XNOR2_X1 U544 ( .A(n405), .B(n404), .ZN(n403) );
  INV_X1 U545 ( .A(KEYINPUT122), .ZN(n404) );
  NAND2_X1 U546 ( .A1(n411), .A2(n409), .ZN(n541) );
  INV_X1 U547 ( .A(n540), .ZN(n409) );
  INV_X1 U548 ( .A(n539), .ZN(n411) );
  NAND2_X1 U549 ( .A1(n412), .A2(n695), .ZN(n566) );
  NAND2_X1 U550 ( .A1(n412), .A2(n697), .ZN(n596) );
  NAND2_X1 U551 ( .A1(n583), .A2(n413), .ZN(n626) );
  XNOR2_X1 U552 ( .A(n415), .B(n473), .ZN(n414) );
  XNOR2_X2 U553 ( .A(n554), .B(n553), .ZN(n620) );
  NAND2_X1 U554 ( .A1(n419), .A2(n420), .ZN(n418) );
  XNOR2_X1 U555 ( .A(n619), .B(KEYINPUT74), .ZN(n419) );
  XNOR2_X1 U556 ( .A(n422), .B(n421), .ZN(n526) );
  INV_X1 U557 ( .A(KEYINPUT83), .ZN(n421) );
  INV_X1 U558 ( .A(n686), .ZN(n423) );
  AND2_X1 U559 ( .A1(n618), .A2(n617), .ZN(G54) );
  INV_X1 U560 ( .A(KEYINPUT47), .ZN(n590) );
  INV_X1 U561 ( .A(KEYINPUT76), .ZN(n440) );
  INV_X1 U562 ( .A(KEYINPUT48), .ZN(n594) );
  XNOR2_X1 U563 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U564 ( .A(n445), .B(n732), .ZN(n611) );
  XNOR2_X1 U565 ( .A(n475), .B(n433), .ZN(n434) );
  XNOR2_X1 U566 ( .A(KEYINPUT111), .B(KEYINPUT28), .ZN(n570) );
  XNOR2_X1 U567 ( .A(KEYINPUT97), .B(KEYINPUT31), .ZN(n529) );
  INV_X1 U568 ( .A(n716), .ZN(n617) );
  INV_X1 U569 ( .A(KEYINPUT42), .ZN(n575) );
  XOR2_X1 U570 ( .A(KEYINPUT96), .B(KEYINPUT5), .Z(n428) );
  XNOR2_X1 U571 ( .A(G116), .B(G113), .ZN(n430) );
  XNOR2_X1 U572 ( .A(G101), .B(KEYINPUT69), .ZN(n429) );
  XNOR2_X1 U573 ( .A(n430), .B(n429), .ZN(n432) );
  XNOR2_X1 U574 ( .A(n432), .B(n431), .ZN(n475) );
  NAND2_X1 U575 ( .A1(G210), .A2(n494), .ZN(n433) );
  NAND2_X1 U576 ( .A1(n665), .A2(n478), .ZN(n435) );
  INV_X1 U577 ( .A(KEYINPUT6), .ZN(n436) );
  XNOR2_X1 U578 ( .A(G110), .B(G107), .ZN(n438) );
  NAND2_X1 U579 ( .A1(G227), .A2(n717), .ZN(n441) );
  XOR2_X1 U580 ( .A(G140), .B(G137), .Z(n452) );
  INV_X1 U581 ( .A(n452), .ZN(n443) );
  XNOR2_X1 U582 ( .A(n444), .B(n443), .ZN(n732) );
  INV_X1 U583 ( .A(G469), .ZN(n446) );
  XNOR2_X2 U584 ( .A(n447), .B(n446), .ZN(n572) );
  INV_X1 U585 ( .A(KEYINPUT1), .ZN(n448) );
  NAND2_X1 U586 ( .A1(n458), .A2(G221), .ZN(n451) );
  XOR2_X1 U587 ( .A(KEYINPUT93), .B(KEYINPUT21), .Z(n450) );
  XNOR2_X1 U588 ( .A(n451), .B(n450), .ZN(n630) );
  XNOR2_X1 U589 ( .A(n630), .B(KEYINPUT94), .ZN(n515) );
  XOR2_X1 U590 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n454) );
  XOR2_X1 U591 ( .A(n454), .B(n453), .Z(n455) );
  NAND2_X1 U592 ( .A1(G234), .A2(n717), .ZN(n456) );
  XOR2_X1 U593 ( .A(KEYINPUT8), .B(n456), .Z(n507) );
  NAND2_X1 U594 ( .A1(G221), .A2(n507), .ZN(n457) );
  NOR2_X1 U595 ( .A1(n713), .A2(G902), .ZN(n462) );
  XOR2_X1 U596 ( .A(KEYINPUT92), .B(KEYINPUT25), .Z(n459) );
  XNOR2_X1 U597 ( .A(n465), .B(n464), .ZN(n467) );
  XNOR2_X1 U598 ( .A(n466), .B(n467), .ZN(n472) );
  XNOR2_X1 U599 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U600 ( .A(KEYINPUT16), .B(G122), .ZN(n474) );
  XNOR2_X1 U601 ( .A(n475), .B(n474), .ZN(n724) );
  INV_X1 U602 ( .A(n607), .ZN(n476) );
  NAND2_X1 U603 ( .A1(n478), .A2(n477), .ZN(n480) );
  AND2_X1 U604 ( .A1(n480), .A2(G210), .ZN(n479) );
  NAND2_X1 U605 ( .A1(n480), .A2(G214), .ZN(n638) );
  XNOR2_X1 U606 ( .A(KEYINPUT75), .B(KEYINPUT19), .ZN(n481) );
  XOR2_X1 U607 ( .A(KEYINPUT14), .B(KEYINPUT87), .Z(n483) );
  NAND2_X1 U608 ( .A1(G237), .A2(G234), .ZN(n482) );
  XNOR2_X1 U609 ( .A(n483), .B(n482), .ZN(n485) );
  NAND2_X1 U610 ( .A1(G952), .A2(n485), .ZN(n484) );
  XNOR2_X1 U611 ( .A(n484), .B(KEYINPUT88), .ZN(n654) );
  NOR2_X1 U612 ( .A1(n654), .A2(G953), .ZN(n556) );
  NAND2_X1 U613 ( .A1(G902), .A2(n485), .ZN(n557) );
  INV_X1 U614 ( .A(n557), .ZN(n486) );
  NOR2_X1 U615 ( .A1(G898), .A2(n717), .ZN(n725) );
  NAND2_X1 U616 ( .A1(n486), .A2(n725), .ZN(n487) );
  XNOR2_X1 U617 ( .A(n487), .B(KEYINPUT89), .ZN(n488) );
  NOR2_X1 U618 ( .A1(n556), .A2(n488), .ZN(n489) );
  NAND2_X1 U619 ( .A1(n648), .A2(n528), .ZN(n491) );
  XNOR2_X1 U620 ( .A(KEYINPUT71), .B(KEYINPUT34), .ZN(n490) );
  XNOR2_X1 U621 ( .A(n491), .B(n490), .ZN(n512) );
  XNOR2_X1 U622 ( .A(n493), .B(n492), .ZN(n500) );
  NAND2_X1 U623 ( .A1(n494), .A2(G214), .ZN(n496) );
  XNOR2_X1 U624 ( .A(n496), .B(n495), .ZN(n498) );
  XNOR2_X1 U625 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U626 ( .A(KEYINPUT101), .B(KEYINPUT13), .ZN(n501) );
  XOR2_X1 U627 ( .A(KEYINPUT105), .B(G478), .Z(n511) );
  XNOR2_X1 U628 ( .A(n503), .B(n502), .ZN(n504) );
  XOR2_X1 U629 ( .A(n504), .B(KEYINPUT9), .Z(n505) );
  NAND2_X1 U630 ( .A1(G217), .A2(n507), .ZN(n508) );
  XNOR2_X1 U631 ( .A(n509), .B(n508), .ZN(n709) );
  NOR2_X1 U632 ( .A1(G902), .A2(n709), .ZN(n510) );
  NOR2_X1 U633 ( .A1(n538), .A2(n539), .ZN(n580) );
  NAND2_X1 U634 ( .A1(n512), .A2(n580), .ZN(n514) );
  INV_X1 U635 ( .A(KEYINPUT35), .ZN(n513) );
  NAND2_X1 U636 ( .A1(n538), .A2(n539), .ZN(n641) );
  XNOR2_X1 U637 ( .A(KEYINPUT65), .B(KEYINPUT22), .ZN(n517) );
  AND2_X1 U638 ( .A1(n600), .A2(n520), .ZN(n521) );
  XNOR2_X1 U639 ( .A(KEYINPUT79), .B(KEYINPUT32), .ZN(n522) );
  XNOR2_X1 U640 ( .A(n522), .B(KEYINPUT64), .ZN(n523) );
  NOR2_X1 U641 ( .A1(n600), .A2(n340), .ZN(n525) );
  NAND2_X1 U642 ( .A1(n527), .A2(n340), .ZN(n625) );
  INV_X1 U643 ( .A(n528), .ZN(n532) );
  NOR2_X1 U644 ( .A1(n625), .A2(n532), .ZN(n530) );
  XNOR2_X1 U645 ( .A(n531), .B(KEYINPUT95), .ZN(n563) );
  OR2_X1 U646 ( .A1(n563), .A2(n340), .ZN(n533) );
  NOR2_X1 U647 ( .A1(n533), .A2(n532), .ZN(n682) );
  OR2_X1 U648 ( .A1(n584), .A2(n629), .ZN(n534) );
  NOR2_X1 U649 ( .A1(n600), .A2(n534), .ZN(n536) );
  OR2_X1 U650 ( .A1(n694), .A2(n537), .ZN(n544) );
  AND2_X1 U651 ( .A1(n540), .A2(n539), .ZN(n695) );
  INV_X1 U652 ( .A(n695), .ZN(n691) );
  NAND2_X1 U653 ( .A1(n542), .A2(n643), .ZN(n543) );
  NAND2_X1 U654 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U655 ( .A1(n547), .A2(n546), .ZN(n549) );
  INV_X1 U656 ( .A(KEYINPUT82), .ZN(n548) );
  XNOR2_X1 U657 ( .A(n549), .B(n548), .ZN(n552) );
  OR2_X1 U658 ( .A1(n550), .A2(KEYINPUT44), .ZN(n551) );
  NAND2_X1 U659 ( .A1(n552), .A2(n551), .ZN(n554) );
  INV_X1 U660 ( .A(KEYINPUT45), .ZN(n553) );
  NAND2_X1 U661 ( .A1(n569), .A2(n638), .ZN(n555) );
  XOR2_X1 U662 ( .A(KEYINPUT30), .B(n555), .Z(n561) );
  INV_X1 U663 ( .A(n556), .ZN(n560) );
  NOR2_X1 U664 ( .A1(G900), .A2(n557), .ZN(n558) );
  NAND2_X1 U665 ( .A1(G953), .A2(n558), .ZN(n559) );
  NAND2_X1 U666 ( .A1(n560), .A2(n559), .ZN(n567) );
  NAND2_X1 U667 ( .A1(n561), .A2(n567), .ZN(n562) );
  XOR2_X1 U668 ( .A(KEYINPUT81), .B(KEYINPUT39), .Z(n564) );
  NAND2_X1 U669 ( .A1(n567), .A2(n629), .ZN(n568) );
  AND2_X1 U670 ( .A1(n340), .A2(n585), .ZN(n571) );
  XNOR2_X1 U671 ( .A(n571), .B(n570), .ZN(n573) );
  NOR2_X1 U672 ( .A1(n573), .A2(n572), .ZN(n589) );
  NAND2_X1 U673 ( .A1(n639), .A2(n638), .ZN(n574) );
  XNOR2_X2 U674 ( .A(n576), .B(n575), .ZN(n744) );
  NAND2_X1 U675 ( .A1(n577), .A2(n380), .ZN(n579) );
  NAND2_X1 U676 ( .A1(n579), .A2(n578), .ZN(n593) );
  AND2_X1 U677 ( .A1(n581), .A2(n580), .ZN(n582) );
  AND2_X1 U678 ( .A1(n602), .A2(n582), .ZN(n678) );
  INV_X1 U679 ( .A(n678), .ZN(n591) );
  NOR2_X1 U680 ( .A1(n597), .A2(n586), .ZN(n587) );
  NAND2_X1 U681 ( .A1(n589), .A2(n396), .ZN(n692) );
  NAND2_X1 U682 ( .A1(n593), .A2(n592), .ZN(n595) );
  XNOR2_X1 U683 ( .A(n595), .B(n594), .ZN(n606) );
  INV_X1 U684 ( .A(n687), .ZN(n697) );
  XOR2_X1 U685 ( .A(KEYINPUT114), .B(n596), .Z(n743) );
  INV_X1 U686 ( .A(n597), .ZN(n598) );
  NAND2_X1 U687 ( .A1(n598), .A2(n638), .ZN(n599) );
  INV_X1 U688 ( .A(n602), .ZN(n603) );
  NOR2_X1 U689 ( .A1(n743), .A2(n663), .ZN(n605) );
  INV_X1 U690 ( .A(n620), .ZN(n718) );
  NOR2_X1 U691 ( .A1(n608), .A2(n420), .ZN(n609) );
  NAND2_X1 U692 ( .A1(n718), .A2(n609), .ZN(n622) );
  AND2_X2 U693 ( .A1(n610), .A2(n622), .ZN(n701) );
  NAND2_X1 U694 ( .A1(n712), .A2(G469), .ZN(n615) );
  XOR2_X1 U695 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n613) );
  XNOR2_X1 U696 ( .A(n611), .B(KEYINPUT123), .ZN(n612) );
  XNOR2_X1 U697 ( .A(n613), .B(n612), .ZN(n614) );
  INV_X1 U698 ( .A(G952), .ZN(n616) );
  NOR2_X1 U699 ( .A1(n620), .A2(n733), .ZN(n621) );
  INV_X1 U700 ( .A(n622), .ZN(n623) );
  INV_X1 U701 ( .A(n625), .ZN(n635) );
  XNOR2_X1 U702 ( .A(n626), .B(KEYINPUT50), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n628), .A2(n627), .ZN(n633) );
  NAND2_X1 U704 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U705 ( .A(KEYINPUT49), .B(n631), .ZN(n632) );
  NOR2_X1 U706 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U707 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U708 ( .A(n636), .B(KEYINPUT51), .ZN(n637) );
  NAND2_X1 U709 ( .A1(n637), .A2(n655), .ZN(n651) );
  NOR2_X1 U710 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U711 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U712 ( .A(n642), .B(KEYINPUT118), .ZN(n646) );
  NOR2_X1 U713 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U714 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U715 ( .A(KEYINPUT119), .B(n647), .ZN(n649) );
  NAND2_X1 U716 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U717 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U718 ( .A(KEYINPUT52), .B(n652), .Z(n653) );
  NOR2_X1 U719 ( .A1(n654), .A2(n653), .ZN(n658) );
  NAND2_X1 U720 ( .A1(n655), .A2(n648), .ZN(n656) );
  XOR2_X1 U721 ( .A(KEYINPUT120), .B(n656), .Z(n657) );
  NOR2_X1 U722 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U723 ( .A(n659), .B(KEYINPUT121), .ZN(n660) );
  XOR2_X1 U724 ( .A(n662), .B(G119), .Z(G21) );
  XOR2_X1 U725 ( .A(n663), .B(G140), .Z(G42) );
  AND2_X1 U726 ( .A1(n701), .A2(G472), .ZN(n667) );
  XNOR2_X1 U727 ( .A(KEYINPUT85), .B(KEYINPUT62), .ZN(n664) );
  XNOR2_X1 U728 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U729 ( .A(KEYINPUT115), .B(KEYINPUT63), .ZN(n669) );
  XNOR2_X1 U730 ( .A(n670), .B(n669), .ZN(G57) );
  AND2_X1 U731 ( .A1(n701), .A2(G475), .ZN(n673) );
  XNOR2_X1 U732 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U733 ( .A(KEYINPUT124), .B(KEYINPUT60), .ZN(n675) );
  XNOR2_X1 U734 ( .A(n675), .B(KEYINPUT66), .ZN(n676) );
  XNOR2_X1 U735 ( .A(n677), .B(n676), .ZN(G60) );
  XNOR2_X1 U736 ( .A(n679), .B(n678), .ZN(G45) );
  NAND2_X1 U737 ( .A1(n682), .A2(n695), .ZN(n680) );
  XNOR2_X1 U738 ( .A(n680), .B(KEYINPUT116), .ZN(n681) );
  XNOR2_X1 U739 ( .A(G104), .B(n681), .ZN(G6) );
  XOR2_X1 U740 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n684) );
  NAND2_X1 U741 ( .A1(n682), .A2(n697), .ZN(n683) );
  XNOR2_X1 U742 ( .A(n684), .B(n683), .ZN(n685) );
  XNOR2_X1 U743 ( .A(G107), .B(n685), .ZN(G9) );
  XNOR2_X1 U744 ( .A(G110), .B(n686), .ZN(G12) );
  NOR2_X1 U745 ( .A1(n692), .A2(n687), .ZN(n689) );
  XNOR2_X1 U746 ( .A(KEYINPUT117), .B(KEYINPUT29), .ZN(n688) );
  XNOR2_X1 U747 ( .A(n689), .B(n688), .ZN(n690) );
  XOR2_X1 U748 ( .A(G128), .B(n690), .Z(G30) );
  NOR2_X1 U749 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U750 ( .A(G146), .B(n693), .Z(G48) );
  NAND2_X1 U751 ( .A1(n694), .A2(n695), .ZN(n696) );
  XNOR2_X1 U752 ( .A(n696), .B(G113), .ZN(G15) );
  NAND2_X1 U753 ( .A1(n697), .A2(n694), .ZN(n698) );
  XNOR2_X1 U754 ( .A(n698), .B(G116), .ZN(G18) );
  XNOR2_X1 U755 ( .A(G125), .B(n699), .ZN(n700) );
  XNOR2_X1 U756 ( .A(n700), .B(KEYINPUT37), .ZN(G27) );
  NAND2_X1 U757 ( .A1(n701), .A2(G210), .ZN(n706) );
  XNOR2_X1 U758 ( .A(KEYINPUT55), .B(KEYINPUT84), .ZN(n702) );
  XOR2_X1 U759 ( .A(n702), .B(KEYINPUT54), .Z(n703) );
  XNOR2_X1 U760 ( .A(n704), .B(n703), .ZN(n705) );
  XNOR2_X1 U761 ( .A(n706), .B(n705), .ZN(n707) );
  XNOR2_X1 U762 ( .A(n708), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U763 ( .A1(n712), .A2(G478), .ZN(n710) );
  XNOR2_X1 U764 ( .A(n710), .B(n709), .ZN(n711) );
  NOR2_X1 U765 ( .A1(n716), .A2(n711), .ZN(G63) );
  NAND2_X1 U766 ( .A1(n712), .A2(G217), .ZN(n714) );
  XNOR2_X1 U767 ( .A(n714), .B(n713), .ZN(n715) );
  NOR2_X1 U768 ( .A1(n716), .A2(n715), .ZN(G66) );
  NAND2_X1 U769 ( .A1(n718), .A2(n717), .ZN(n722) );
  NAND2_X1 U770 ( .A1(G953), .A2(G224), .ZN(n719) );
  XNOR2_X1 U771 ( .A(KEYINPUT61), .B(n719), .ZN(n720) );
  NAND2_X1 U772 ( .A1(n720), .A2(G898), .ZN(n721) );
  NAND2_X1 U773 ( .A1(n722), .A2(n721), .ZN(n729) );
  XNOR2_X1 U774 ( .A(n724), .B(n723), .ZN(n726) );
  NOR2_X1 U775 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U776 ( .A(KEYINPUT126), .B(n727), .Z(n728) );
  XNOR2_X1 U777 ( .A(n729), .B(n728), .ZN(n730) );
  XNOR2_X1 U778 ( .A(KEYINPUT125), .B(n730), .ZN(G69) );
  XNOR2_X1 U779 ( .A(n732), .B(n731), .ZN(n736) );
  XOR2_X1 U780 ( .A(n733), .B(n736), .Z(n734) );
  NOR2_X1 U781 ( .A1(G953), .A2(n734), .ZN(n735) );
  XNOR2_X1 U782 ( .A(n735), .B(KEYINPUT127), .ZN(n740) );
  XNOR2_X1 U783 ( .A(G227), .B(n736), .ZN(n737) );
  NAND2_X1 U784 ( .A1(n737), .A2(G900), .ZN(n738) );
  NAND2_X1 U785 ( .A1(n738), .A2(G953), .ZN(n739) );
  NAND2_X1 U786 ( .A1(n740), .A2(n739), .ZN(G72) );
  XNOR2_X1 U787 ( .A(n741), .B(G122), .ZN(G24) );
  XOR2_X1 U788 ( .A(n742), .B(G131), .Z(G33) );
  XOR2_X1 U789 ( .A(G134), .B(n743), .Z(G36) );
  XOR2_X1 U790 ( .A(G137), .B(n744), .Z(G39) );
endmodule

