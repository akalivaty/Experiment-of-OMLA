//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 0 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 1 1 1 1 0 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1201,
    new_n1202, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  AND2_X1   g0009(.A1(G116), .A2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G77), .ZN(new_n211));
  INV_X1    g0011(.A(G244), .ZN(new_n212));
  INV_X1    g0012(.A(G97), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  OAI22_X1  g0014(.A1(new_n211), .A2(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n210), .B(new_n215), .C1(G87), .C2(G250), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G58), .A2(G232), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G107), .A2(G264), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G50), .A2(G226), .ZN(new_n219));
  NAND4_X1  g0019(.A1(new_n216), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n206), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(G50), .B1(G58), .B2(G68), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n209), .B(new_n225), .C1(new_n228), .C2(new_n230), .ZN(G361));
  XOR2_X1   g0031(.A(KEYINPUT64), .B(KEYINPUT2), .Z(new_n232));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G226), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n237), .B(new_n238), .Z(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  NAND2_X1  g0047(.A1(new_n203), .A2(G20), .ZN(new_n248));
  INV_X1    g0048(.A(G150), .ZN(new_n249));
  NOR2_X1   g0049(.A1(G20), .A2(G33), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(G20), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT8), .B(G58), .ZN(new_n255));
  OAI221_X1 g0055(.A(new_n248), .B1(new_n249), .B2(new_n251), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n226), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(G13), .A3(G20), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n202), .ZN(new_n263));
  INV_X1    g0063(.A(new_n258), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n264), .B1(G1), .B2(new_n227), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n259), .B(new_n263), .C1(new_n202), .C2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT67), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n266), .A2(new_n267), .ZN(new_n270));
  OAI21_X1  g0070(.A(KEYINPUT9), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  OR2_X1    g0071(.A1(new_n266), .A2(new_n267), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT9), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n272), .A2(new_n273), .A3(new_n268), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT3), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n252), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G222), .A2(G1698), .ZN(new_n279));
  INV_X1    g0079(.A(G1698), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(G223), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n278), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G41), .ZN(new_n283));
  OAI211_X1 g0083(.A(G1), .B(G13), .C1(new_n252), .C2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n282), .B(new_n285), .C1(G77), .C2(new_n278), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n260), .B1(G41), .B2(G45), .ZN(new_n287));
  INV_X1    g0087(.A(G274), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G226), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n284), .A2(new_n287), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n286), .B(new_n290), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G200), .ZN(new_n294));
  INV_X1    g0094(.A(G190), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n271), .A2(new_n274), .A3(new_n294), .A4(new_n296), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n297), .B(KEYINPUT10), .ZN(new_n298));
  XNOR2_X1  g0098(.A(KEYINPUT65), .B(G179), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n293), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n293), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n300), .A2(new_n266), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n299), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n278), .A2(G232), .A3(new_n280), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n278), .A2(G238), .A3(G1698), .ZN(new_n306));
  INV_X1    g0106(.A(G107), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n305), .B(new_n306), .C1(new_n307), .C2(new_n278), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n289), .B1(new_n308), .B2(new_n285), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n284), .A2(new_n287), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G244), .ZN(new_n311));
  AND3_X1   g0111(.A1(new_n309), .A2(KEYINPUT66), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(KEYINPUT66), .B1(new_n309), .B2(new_n311), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n304), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n308), .A2(new_n285), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n315), .A2(new_n290), .A3(new_n311), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT66), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n309), .A2(KEYINPUT66), .A3(new_n311), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n318), .A2(new_n301), .A3(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n265), .A2(new_n211), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n261), .A2(G77), .ZN(new_n322));
  INV_X1    g0122(.A(new_n255), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n323), .A2(new_n250), .B1(G20), .B2(G77), .ZN(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT15), .B(G87), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n324), .B1(new_n254), .B2(new_n325), .ZN(new_n326));
  AOI211_X1 g0126(.A(new_n321), .B(new_n322), .C1(new_n326), .C2(new_n258), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n314), .A2(new_n320), .A3(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(G190), .B1(new_n312), .B2(new_n313), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n318), .A2(G200), .A3(new_n319), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n330), .A2(new_n327), .A3(new_n331), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n298), .A2(new_n303), .A3(new_n329), .A4(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT16), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n276), .A2(new_n227), .A3(new_n277), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT7), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n276), .A2(KEYINPUT7), .A3(new_n227), .A4(new_n277), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n221), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G58), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n340), .A2(new_n221), .ZN(new_n341));
  OAI21_X1  g0141(.A(G20), .B1(new_n341), .B2(new_n201), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n250), .A2(G159), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n334), .B1(new_n339), .B2(new_n344), .ZN(new_n345));
  AND2_X1   g0145(.A1(KEYINPUT3), .A2(G33), .ZN(new_n346));
  NOR2_X1   g0146(.A1(KEYINPUT3), .A2(G33), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(KEYINPUT7), .B1(new_n348), .B2(new_n227), .ZN(new_n349));
  INV_X1    g0149(.A(new_n338), .ZN(new_n350));
  OAI21_X1  g0150(.A(G68), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n344), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(KEYINPUT16), .A3(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n345), .A2(new_n353), .A3(new_n258), .ZN(new_n354));
  MUX2_X1   g0154(.A(new_n261), .B(new_n265), .S(new_n323), .Z(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n291), .A2(G1698), .ZN(new_n357));
  OAI221_X1 g0157(.A(new_n357), .B1(G223), .B2(G1698), .C1(new_n346), .C2(new_n347), .ZN(new_n358));
  NAND2_X1  g0158(.A1(G33), .A2(G87), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n285), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n289), .B1(new_n310), .B2(G232), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(G169), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(new_n363), .B2(new_n304), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n356), .A2(KEYINPUT18), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(KEYINPUT18), .B1(new_n356), .B2(new_n365), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n361), .A2(new_n362), .A3(new_n295), .ZN(new_n369));
  INV_X1    g0169(.A(G200), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n284), .B1(new_n358), .B2(new_n359), .ZN(new_n371));
  INV_X1    g0171(.A(G232), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n290), .B1(new_n292), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n370), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n369), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n354), .A2(new_n355), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT17), .ZN(new_n377));
  XNOR2_X1  g0177(.A(new_n376), .B(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n368), .A2(new_n378), .ZN(new_n379));
  OR2_X1    g0179(.A1(new_n379), .A2(KEYINPUT69), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT13), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n372), .A2(G1698), .ZN(new_n382));
  OAI221_X1 g0182(.A(new_n382), .B1(G226), .B2(G1698), .C1(new_n346), .C2(new_n347), .ZN(new_n383));
  NAND2_X1  g0183(.A1(G33), .A2(G97), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n289), .B1(new_n385), .B2(new_n285), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n284), .A2(G238), .A3(new_n287), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n381), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n284), .B1(new_n383), .B2(new_n384), .ZN(new_n390));
  NOR4_X1   g0190(.A1(new_n390), .A2(KEYINPUT13), .A3(new_n387), .A4(new_n289), .ZN(new_n391));
  OAI21_X1  g0191(.A(G169), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(KEYINPUT14), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n389), .A2(new_n391), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(G179), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT14), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n396), .B(G169), .C1(new_n389), .C2(new_n391), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n393), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n253), .A2(G77), .B1(G20), .B2(new_n221), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n250), .A2(G50), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n264), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  XOR2_X1   g0201(.A(new_n401), .B(KEYINPUT11), .Z(new_n402));
  NOR2_X1   g0202(.A1(new_n261), .A2(G68), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT12), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n405), .B(KEYINPUT68), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(new_n404), .B2(new_n403), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n402), .B(new_n407), .C1(new_n221), .C2(new_n265), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n398), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n408), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n394), .A2(G190), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n410), .B(new_n411), .C1(new_n370), .C2(new_n394), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n379), .A2(KEYINPUT69), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n380), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  OAI211_X1 g0215(.A(G257), .B(new_n280), .C1(new_n346), .C2(new_n347), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT75), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n278), .A2(KEYINPUT75), .A3(G257), .A4(new_n280), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n278), .A2(G264), .A3(G1698), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n348), .A2(G303), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n418), .A2(new_n419), .A3(new_n420), .A4(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n285), .ZN(new_n423));
  INV_X1    g0223(.A(G45), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n424), .A2(G1), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n283), .A2(KEYINPUT5), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT5), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(G41), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n425), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n429), .A2(G270), .A3(new_n284), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n425), .A2(new_n426), .A3(new_n428), .A4(G274), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n423), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n261), .A2(G116), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n260), .A2(G33), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n261), .A2(new_n436), .A3(new_n226), .A4(new_n257), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n435), .B1(new_n438), .B2(G116), .ZN(new_n439));
  AOI21_X1  g0239(.A(G20), .B1(G33), .B2(G283), .ZN(new_n440));
  OR2_X1    g0240(.A1(KEYINPUT71), .A2(G97), .ZN(new_n441));
  NAND2_X1  g0241(.A1(KEYINPUT71), .A2(G97), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n440), .B1(new_n443), .B2(G33), .ZN(new_n444));
  INV_X1    g0244(.A(G116), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n257), .A2(new_n226), .B1(G20), .B2(new_n445), .ZN(new_n446));
  AND3_X1   g0246(.A1(new_n444), .A2(KEYINPUT20), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(KEYINPUT20), .B1(new_n444), .B2(new_n446), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n439), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n434), .A2(KEYINPUT21), .A3(new_n449), .A4(G169), .ZN(new_n450));
  INV_X1    g0250(.A(G179), .ZN(new_n451));
  AOI211_X1 g0251(.A(new_n451), .B(new_n432), .C1(new_n422), .C2(new_n285), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n449), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT76), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n253), .A2(G116), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n227), .A2(G107), .ZN(new_n457));
  XNOR2_X1  g0257(.A(new_n457), .B(KEYINPUT23), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n227), .B(G87), .C1(new_n346), .C2(new_n347), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n459), .A2(KEYINPUT22), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n459), .A2(KEYINPUT22), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n456), .B(new_n458), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT24), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g0264(.A(new_n459), .B(KEYINPUT22), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n465), .A2(KEYINPUT24), .A3(new_n456), .A4(new_n458), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n464), .A2(new_n258), .A3(new_n466), .ZN(new_n467));
  OR3_X1    g0267(.A1(new_n261), .A2(KEYINPUT25), .A3(G107), .ZN(new_n468));
  OAI21_X1  g0268(.A(KEYINPUT25), .B1(new_n261), .B2(G107), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n468), .B(new_n469), .C1(new_n307), .C2(new_n437), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT77), .ZN(new_n471));
  XNOR2_X1  g0271(.A(new_n470), .B(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  OAI211_X1 g0273(.A(G257), .B(G1698), .C1(new_n346), .C2(new_n347), .ZN(new_n474));
  OAI211_X1 g0274(.A(G250), .B(new_n280), .C1(new_n346), .C2(new_n347), .ZN(new_n475));
  INV_X1    g0275(.A(G294), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n474), .B(new_n475), .C1(new_n252), .C2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n285), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n429), .A2(new_n284), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(G264), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n478), .A2(new_n431), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n301), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n481), .A2(G179), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n473), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n434), .A2(G169), .A3(new_n449), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT21), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT76), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n450), .A2(new_n453), .A3(new_n489), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n455), .A2(new_n485), .A3(new_n488), .A4(new_n490), .ZN(new_n491));
  NOR4_X1   g0291(.A1(new_n211), .A2(KEYINPUT70), .A3(G20), .A4(G33), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT70), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n493), .B1(new_n250), .B2(G77), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT6), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n496), .B1(new_n441), .B2(new_n442), .ZN(new_n497));
  OAI21_X1  g0297(.A(G107), .B1(new_n213), .B2(KEYINPUT6), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n496), .A2(new_n307), .A3(G97), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n495), .B1(new_n501), .B2(G20), .ZN(new_n502));
  OAI21_X1  g0302(.A(G107), .B1(new_n349), .B2(new_n350), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n264), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n437), .A2(G97), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n261), .A2(new_n213), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n505), .A2(KEYINPUT72), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(KEYINPUT72), .B1(new_n505), .B2(new_n506), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(KEYINPUT73), .B1(new_n504), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n442), .ZN(new_n511));
  NOR2_X1   g0311(.A1(KEYINPUT71), .A2(G97), .ZN(new_n512));
  OAI21_X1  g0312(.A(KEYINPUT6), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n513), .A2(G20), .A3(new_n498), .A4(new_n499), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n514), .B1(new_n494), .B2(new_n492), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n307), .B1(new_n337), .B2(new_n338), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n258), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n505), .A2(new_n506), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT72), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n505), .A2(KEYINPUT72), .A3(new_n506), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT73), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n517), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n510), .A2(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(G244), .B(new_n280), .C1(new_n346), .C2(new_n347), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT4), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n278), .A2(KEYINPUT4), .A3(G244), .A4(new_n280), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n278), .A2(G250), .A3(G1698), .ZN(new_n531));
  NAND2_X1  g0331(.A1(G33), .A2(G283), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n285), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n429), .A2(new_n284), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n431), .B1(new_n535), .B2(new_n214), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n534), .A2(new_n299), .A3(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n528), .A2(new_n529), .A3(new_n532), .A4(new_n531), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n536), .B1(new_n539), .B2(new_n285), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n538), .B1(new_n301), .B2(new_n540), .ZN(new_n541));
  AOI211_X1 g0341(.A(new_n295), .B(new_n536), .C1(new_n285), .C2(new_n539), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n370), .B1(new_n534), .B2(new_n537), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n504), .A2(new_n509), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n525), .A2(new_n541), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n481), .A2(new_n370), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n477), .A2(new_n285), .B1(new_n479), .B2(G264), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n548), .A2(new_n295), .A3(new_n431), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n550), .A2(new_n472), .A3(new_n467), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n325), .A2(new_n262), .ZN(new_n552));
  INV_X1    g0352(.A(G87), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n553), .B(new_n307), .C1(new_n511), .C2(new_n512), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT19), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n227), .B1(new_n384), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n555), .B1(new_n443), .B2(new_n254), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n278), .A2(new_n227), .A3(G68), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n552), .B1(new_n560), .B2(new_n258), .ZN(new_n561));
  XNOR2_X1  g0361(.A(new_n325), .B(KEYINPUT74), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n438), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n260), .A2(G45), .ZN(new_n564));
  AND2_X1   g0364(.A1(G33), .A2(G41), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n564), .B(G250), .C1(new_n565), .C2(new_n226), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n222), .A2(new_n280), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n212), .A2(G1698), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n568), .B(new_n569), .C1(new_n346), .C2(new_n347), .ZN(new_n570));
  NAND2_X1  g0370(.A1(G33), .A2(G116), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n567), .B1(new_n572), .B2(new_n285), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n564), .A2(new_n288), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n561), .A2(new_n563), .B1(new_n576), .B2(new_n301), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n284), .B1(new_n570), .B2(new_n571), .ZN(new_n578));
  NOR3_X1   g0378(.A1(new_n578), .A2(new_n574), .A3(new_n567), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n304), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n370), .B1(new_n573), .B2(new_n575), .ZN(new_n581));
  NOR4_X1   g0381(.A1(new_n578), .A2(new_n295), .A3(new_n567), .A4(new_n574), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n437), .A2(new_n553), .ZN(new_n584));
  AOI211_X1 g0384(.A(new_n552), .B(new_n584), .C1(new_n560), .C2(new_n258), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n577), .A2(new_n580), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n449), .B1(new_n434), .B2(G200), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(new_n295), .B2(new_n434), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n546), .A2(new_n551), .A3(new_n586), .A4(new_n588), .ZN(new_n589));
  NOR4_X1   g0389(.A1(new_n333), .A2(new_n415), .A3(new_n491), .A4(new_n589), .ZN(G372));
  NOR2_X1   g0390(.A1(new_n333), .A2(new_n415), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n517), .A2(new_n522), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n541), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT80), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n541), .A2(KEYINPUT80), .A3(new_n592), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n595), .A2(new_n586), .A3(new_n596), .ZN(new_n597));
  OR2_X1    g0397(.A1(new_n597), .A2(KEYINPUT26), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n577), .A2(new_n580), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n586), .A2(new_n541), .A3(new_n525), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n600), .B1(new_n601), .B2(KEYINPUT26), .ZN(new_n602));
  NOR3_X1   g0402(.A1(new_n504), .A2(new_n509), .A3(KEYINPUT73), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n523), .B1(new_n517), .B2(new_n522), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n541), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n540), .A2(G190), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n545), .B(new_n606), .C1(new_n370), .C2(new_n540), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n605), .A2(new_n586), .A3(new_n551), .A4(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(KEYINPUT78), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT78), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n546), .A2(new_n610), .A3(new_n551), .A4(new_n586), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT79), .ZN(new_n613));
  AOI221_X4 g0413(.A(new_n483), .B1(new_n301), .B2(new_n481), .C1(new_n467), .C2(new_n472), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n488), .A2(new_n450), .A3(new_n453), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n454), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n617), .A2(new_n485), .A3(KEYINPUT79), .A4(new_n488), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n598), .B(new_n602), .C1(new_n612), .C2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n591), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g0421(.A(new_n621), .B(KEYINPUT81), .Z(new_n622));
  NAND2_X1  g0422(.A1(new_n409), .A2(new_n329), .ZN(new_n623));
  XNOR2_X1  g0423(.A(new_n376), .B(KEYINPUT17), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n623), .A2(new_n412), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n356), .A2(new_n365), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT18), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n356), .A2(new_n365), .A3(KEYINPUT18), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n625), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT10), .ZN(new_n632));
  XNOR2_X1  g0432(.A(new_n297), .B(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n303), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT82), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI211_X1 g0436(.A(KEYINPUT82), .B(new_n303), .C1(new_n631), .C2(new_n633), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n622), .A2(new_n638), .ZN(G369));
  INV_X1    g0439(.A(G13), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(G20), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  OR3_X1    g0442(.A1(new_n642), .A2(KEYINPUT27), .A3(G1), .ZN(new_n643));
  OAI21_X1  g0443(.A(KEYINPUT27), .B1(new_n642), .B2(G1), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(G213), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(G343), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n449), .A2(new_n647), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n615), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n588), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n455), .A2(new_n488), .A3(new_n490), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n650), .B1(new_n651), .B2(new_n648), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(G330), .ZN(new_n653));
  INV_X1    g0453(.A(new_n551), .ZN(new_n654));
  INV_X1    g0454(.A(new_n647), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n655), .B1(new_n467), .B2(new_n472), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n485), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n614), .A2(new_n655), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n653), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n657), .A2(new_n651), .A3(new_n485), .A4(new_n655), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n658), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n661), .A2(new_n664), .ZN(G399));
  NOR2_X1   g0465(.A1(new_n554), .A2(G116), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n207), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(G41), .ZN(new_n669));
  NOR3_X1   g0469(.A1(new_n667), .A2(new_n260), .A3(new_n669), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT83), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n669), .A2(new_n230), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n670), .A2(KEYINPUT83), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n674), .B(KEYINPUT28), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n589), .A2(new_n491), .A3(new_n647), .ZN(new_n676));
  AND3_X1   g0476(.A1(new_n534), .A2(new_n548), .A3(new_n537), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n677), .A2(KEYINPUT30), .A3(new_n452), .A4(new_n579), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT30), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n423), .A2(G179), .A3(new_n579), .A4(new_n433), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n534), .A2(new_n548), .A3(new_n537), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n679), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT84), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n299), .B1(new_n579), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n576), .A2(KEYINPUT84), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n534), .A2(new_n537), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n685), .A2(new_n434), .A3(new_n686), .A4(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n481), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n647), .B1(new_n683), .B2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT31), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OAI211_X1 g0493(.A(KEYINPUT31), .B(new_n647), .C1(new_n683), .C2(new_n690), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n676), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n620), .A2(new_n655), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT29), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n583), .A2(new_n585), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n599), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n605), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT26), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n600), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n597), .A2(KEYINPUT26), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n455), .A2(new_n488), .A3(new_n490), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n608), .B1(new_n709), .B2(new_n485), .ZN(new_n710));
  OAI211_X1 g0510(.A(KEYINPUT29), .B(new_n655), .C1(new_n708), .C2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n697), .B1(new_n701), .B2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n675), .B1(new_n714), .B2(G1), .ZN(G364));
  NAND2_X1  g0515(.A1(new_n299), .A2(G20), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(G190), .A2(G200), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n295), .A2(new_n370), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n227), .A2(G179), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT87), .ZN(new_n724));
  AOI22_X1  g0524(.A1(new_n720), .A2(G311), .B1(new_n724), .B2(G303), .ZN(new_n725));
  INV_X1    g0525(.A(G283), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n370), .A2(G190), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n722), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n295), .A2(G200), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n451), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(G20), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  OAI221_X1 g0532(.A(new_n725), .B1(new_n726), .B2(new_n728), .C1(new_n476), .C2(new_n732), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n716), .A2(G190), .A3(new_n370), .ZN(new_n734));
  XNOR2_X1  g0534(.A(KEYINPUT33), .B(G317), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n717), .A2(new_n729), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G322), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n722), .A2(new_n718), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n278), .B1(new_n741), .B2(G329), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n716), .A2(new_n295), .A3(new_n370), .ZN(new_n743));
  XNOR2_X1  g0543(.A(KEYINPUT86), .B(G326), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n736), .A2(new_n739), .A3(new_n742), .A4(new_n745), .ZN(new_n746));
  AOI22_X1  g0546(.A1(new_n738), .A2(G58), .B1(G50), .B2(new_n743), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n747), .B1(new_n211), .B2(new_n719), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT85), .ZN(new_n749));
  INV_X1    g0549(.A(new_n723), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n749), .B1(G87), .B2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n728), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G107), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n732), .A2(new_n213), .ZN(new_n754));
  AOI211_X1 g0554(.A(new_n348), .B(new_n754), .C1(new_n734), .C2(G68), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n751), .A2(new_n753), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n741), .A2(G159), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT32), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n746), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT88), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n226), .B1(G20), .B2(new_n301), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G13), .A2(G33), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G20), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n761), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n230), .A2(new_n424), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n668), .A2(new_n278), .ZN(new_n767));
  OAI211_X1 g0567(.A(new_n766), .B(new_n767), .C1(new_n246), .C2(new_n424), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n278), .A2(G355), .A3(new_n207), .ZN(new_n769));
  OAI211_X1 g0569(.A(new_n768), .B(new_n769), .C1(G116), .C2(new_n207), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n760), .A2(new_n761), .B1(new_n765), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n260), .B1(new_n641), .B2(G45), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n669), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n764), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n771), .B(new_n774), .C1(new_n652), .C2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n652), .A2(G330), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n653), .B1(new_n669), .B2(new_n773), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(G396));
  INV_X1    g0579(.A(KEYINPUT94), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(new_n327), .B2(new_n655), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n328), .A2(KEYINPUT94), .A3(new_n647), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n329), .A2(new_n332), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n314), .A2(new_n320), .A3(new_n328), .A4(new_n647), .ZN(new_n784));
  AND2_X1   g0584(.A1(new_n784), .A2(KEYINPUT95), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(KEYINPUT95), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n783), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n698), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n620), .A2(new_n655), .A3(new_n787), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(new_n697), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT96), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n793), .B1(new_n669), .B2(new_n773), .C1(new_n697), .C2(new_n791), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n278), .B1(new_n724), .B2(G107), .ZN(new_n795));
  INV_X1    g0595(.A(G303), .ZN(new_n796));
  INV_X1    g0596(.A(new_n743), .ZN(new_n797));
  INV_X1    g0597(.A(G311), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n795), .B1(new_n796), .B2(new_n797), .C1(new_n798), .C2(new_n740), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n754), .B1(new_n738), .B2(G294), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT90), .Z(new_n801));
  XNOR2_X1  g0601(.A(KEYINPUT89), .B(G283), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n799), .B(new_n801), .C1(new_n734), .C2(new_n802), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n803), .B1(new_n553), .B2(new_n728), .C1(new_n445), .C2(new_n719), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT91), .ZN(new_n805));
  XOR2_X1   g0605(.A(KEYINPUT92), .B(G143), .Z(new_n806));
  AOI22_X1  g0606(.A1(new_n720), .A2(G159), .B1(new_n738), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G137), .ZN(new_n808));
  INV_X1    g0608(.A(new_n734), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n807), .B1(new_n808), .B2(new_n797), .C1(new_n249), .C2(new_n809), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT34), .Z(new_n811));
  NOR2_X1   g0611(.A1(new_n728), .A2(new_n221), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(G132), .B2(new_n741), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n813), .B(new_n278), .C1(new_n340), .C2(new_n732), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(G50), .B2(new_n724), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT93), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n805), .B1(new_n811), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n761), .A2(new_n762), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n817), .A2(new_n761), .B1(new_n211), .B2(new_n818), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n819), .B(new_n774), .C1(new_n763), .C2(new_n787), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n794), .A2(new_n820), .ZN(G384));
  INV_X1    g0621(.A(KEYINPUT38), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT37), .ZN(new_n823));
  AND3_X1   g0623(.A1(new_n354), .A2(new_n355), .A3(new_n375), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n645), .B1(new_n354), .B2(new_n355), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n823), .B1(new_n826), .B2(new_n626), .ZN(new_n827));
  INV_X1    g0627(.A(new_n645), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n356), .A2(new_n828), .ZN(new_n829));
  AND4_X1   g0629(.A1(new_n823), .A2(new_n626), .A3(new_n829), .A4(new_n376), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n829), .B1(new_n630), .B2(new_n624), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n822), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n825), .B1(new_n368), .B2(new_n378), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n626), .A2(new_n829), .A3(new_n376), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(KEYINPUT37), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n826), .A2(new_n823), .A3(new_n626), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n834), .A2(new_n838), .A3(KEYINPUT38), .ZN(new_n839));
  AND3_X1   g0639(.A1(new_n833), .A2(KEYINPUT98), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(KEYINPUT98), .B1(new_n833), .B2(new_n839), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n408), .A2(new_n647), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n409), .A2(new_n412), .A3(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n398), .A2(new_n408), .A3(new_n647), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n787), .B(new_n845), .C1(new_n676), .C2(new_n695), .ZN(new_n846));
  NOR3_X1   g0646(.A1(new_n840), .A2(new_n841), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(KEYINPUT99), .B1(new_n847), .B2(KEYINPUT40), .ZN(new_n848));
  INV_X1    g0648(.A(new_n846), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT98), .ZN(new_n850));
  AND3_X1   g0650(.A1(new_n834), .A2(new_n838), .A3(KEYINPUT38), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT38), .B1(new_n834), .B2(new_n838), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n833), .A2(KEYINPUT98), .A3(new_n839), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n849), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT99), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT40), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n848), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n833), .A2(new_n839), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n849), .A2(KEYINPUT40), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n862), .B(KEYINPUT100), .Z(new_n863));
  NAND2_X1  g0663(.A1(new_n591), .A2(new_n696), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n863), .B(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(G330), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT39), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n860), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n833), .A2(KEYINPUT39), .A3(new_n839), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n409), .A2(new_n647), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n870), .A2(new_n871), .B1(new_n368), .B2(new_n645), .ZN(new_n872));
  INV_X1    g0672(.A(new_n845), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n329), .A2(new_n647), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n873), .B1(new_n790), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n876), .A2(new_n853), .A3(new_n854), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n872), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n591), .A2(new_n700), .A3(new_n711), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n638), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n878), .B(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  OAI22_X1  g0682(.A1(new_n866), .A2(new_n882), .B1(new_n260), .B2(new_n641), .ZN(new_n883));
  OR2_X1    g0683(.A1(new_n883), .A2(KEYINPUT101), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n866), .A2(new_n882), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n883), .A2(KEYINPUT101), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n501), .B(KEYINPUT97), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n445), .B1(new_n888), .B2(KEYINPUT35), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n889), .B(new_n228), .C1(KEYINPUT35), .C2(new_n888), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n890), .B(KEYINPUT36), .ZN(new_n891));
  OAI21_X1  g0691(.A(G77), .B1(new_n340), .B2(new_n221), .ZN(new_n892));
  OAI22_X1  g0692(.A1(new_n892), .A2(new_n229), .B1(G50), .B2(new_n221), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n893), .A2(G1), .A3(new_n640), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n887), .A2(new_n891), .A3(new_n894), .ZN(G367));
  INV_X1    g0695(.A(new_n767), .ZN(new_n896));
  OAI221_X1 g0696(.A(new_n765), .B1(new_n207), .B2(new_n325), .C1(new_n239), .C2(new_n896), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n738), .A2(G303), .B1(G107), .B2(new_n731), .ZN(new_n898));
  INV_X1    g0698(.A(new_n802), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n898), .B(new_n348), .C1(new_n719), .C2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(G317), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n740), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n723), .A2(new_n445), .ZN(new_n903));
  OAI22_X1  g0703(.A1(new_n903), .A2(KEYINPUT46), .B1(new_n443), .B2(new_n728), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n809), .A2(new_n476), .ZN(new_n905));
  NOR4_X1   g0705(.A1(new_n900), .A2(new_n902), .A3(new_n904), .A4(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n724), .A2(KEYINPUT46), .A3(G116), .ZN(new_n907));
  XOR2_X1   g0707(.A(new_n907), .B(KEYINPUT108), .Z(new_n908));
  OAI211_X1 g0708(.A(new_n906), .B(new_n908), .C1(new_n798), .C2(new_n797), .ZN(new_n909));
  XOR2_X1   g0709(.A(new_n909), .B(KEYINPUT109), .Z(new_n910));
  AOI22_X1  g0710(.A1(G50), .A2(new_n720), .B1(new_n738), .B2(G150), .ZN(new_n911));
  INV_X1    g0711(.A(new_n806), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n911), .B1(new_n797), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n731), .A2(G68), .ZN(new_n914));
  INV_X1    g0714(.A(G159), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n914), .B1(new_n809), .B2(new_n915), .ZN(new_n916));
  OAI221_X1 g0716(.A(new_n278), .B1(new_n728), .B2(new_n211), .C1(new_n340), .C2(new_n723), .ZN(new_n917));
  NOR3_X1   g0717(.A1(new_n913), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n808), .B2(new_n740), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n910), .A2(new_n919), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n920), .B(KEYINPUT47), .Z(new_n921));
  INV_X1    g0721(.A(new_n761), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n774), .B(new_n897), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n923), .B(KEYINPUT110), .Z(new_n924));
  NOR2_X1   g0724(.A1(new_n585), .A2(new_n655), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT102), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n703), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n600), .B2(new_n926), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n928), .A2(new_n764), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n924), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT107), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n669), .B(KEYINPUT41), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n659), .B1(new_n709), .B2(new_n647), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n652), .A2(G330), .B1(new_n934), .B2(new_n662), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n660), .A2(new_n935), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n936), .B(new_n697), .C1(new_n701), .C2(new_n712), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n546), .B1(new_n545), .B2(new_n655), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n541), .A2(new_n592), .A3(new_n647), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(KEYINPUT105), .B1(new_n664), .B2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT105), .ZN(new_n942));
  INV_X1    g0742(.A(new_n940), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n663), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT44), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n941), .A2(new_n944), .A3(KEYINPUT44), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT104), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n664), .A2(new_n950), .A3(new_n940), .ZN(new_n951));
  OAI21_X1  g0751(.A(KEYINPUT104), .B1(new_n663), .B2(new_n943), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n953), .B(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n937), .B1(new_n949), .B2(new_n956), .ZN(new_n957));
  OAI211_X1 g0757(.A(KEYINPUT106), .B(new_n933), .C1(new_n957), .C2(new_n713), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT106), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n953), .A2(new_n955), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n954), .B1(new_n951), .B2(new_n952), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n947), .B(new_n948), .C1(new_n960), .C2(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n713), .B1(new_n962), .B2(new_n936), .ZN(new_n963));
  INV_X1    g0763(.A(new_n933), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n959), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n958), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n772), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n660), .A2(new_n940), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT43), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n928), .A2(new_n969), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n968), .B(new_n970), .Z(new_n971));
  NOR2_X1   g0771(.A1(new_n662), .A2(new_n938), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT42), .Z(new_n973));
  NAND2_X1  g0773(.A1(new_n940), .A2(new_n614), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n647), .B1(new_n974), .B2(new_n605), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n973), .A2(new_n975), .B1(new_n969), .B2(new_n928), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n971), .B(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n932), .B1(new_n967), .B2(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n773), .B1(new_n958), .B2(new_n965), .ZN(new_n980));
  NOR3_X1   g0780(.A1(new_n980), .A2(KEYINPUT107), .A3(new_n977), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n931), .B1(new_n979), .B2(new_n981), .ZN(G387));
  NAND2_X1  g0782(.A1(new_n659), .A2(new_n764), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n323), .A2(new_n202), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT50), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n666), .B1(new_n221), .B2(new_n211), .ZN(new_n986));
  NOR3_X1   g0786(.A1(new_n985), .A2(G45), .A3(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n236), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n767), .B1(new_n988), .B2(new_n424), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n667), .A2(new_n207), .A3(new_n278), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n987), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n207), .A2(G107), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n765), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n983), .A2(new_n774), .A3(new_n993), .ZN(new_n994));
  AOI22_X1  g0794(.A1(G311), .A2(new_n734), .B1(new_n743), .B2(G322), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n995), .B1(new_n796), .B2(new_n719), .C1(new_n901), .C2(new_n737), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT48), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n997), .B1(new_n476), .B2(new_n723), .C1(new_n732), .C2(new_n899), .ZN(new_n998));
  XOR2_X1   g0798(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n999));
  XNOR2_X1  g0799(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n741), .A2(new_n744), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n278), .B1(new_n752), .B2(G116), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n740), .A2(new_n249), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n797), .A2(new_n915), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n720), .A2(G68), .B1(new_n323), .B2(new_n734), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT111), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n737), .A2(new_n202), .B1(new_n211), .B2(new_n723), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n562), .A2(new_n731), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n1009), .B(new_n278), .C1(new_n213), .C2(new_n728), .ZN(new_n1010));
  OR4_X1    g0810(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .A4(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1003), .B1(new_n1004), .B2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT113), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n994), .B1(new_n1013), .B2(new_n761), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(new_n773), .B2(new_n936), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n713), .B1(new_n660), .B2(new_n935), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1016), .A2(new_n937), .A3(new_n669), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1015), .A2(new_n1017), .ZN(G393));
  INV_X1    g0818(.A(new_n957), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n962), .B(new_n661), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n937), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n669), .B(new_n1019), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1020), .A2(new_n773), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n943), .A2(new_n764), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n765), .B1(new_n207), .B2(new_n443), .C1(new_n243), .C2(new_n896), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n732), .A2(new_n211), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(G50), .B2(new_n734), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n255), .B2(new_n719), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT114), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n912), .A2(new_n740), .B1(new_n728), .B2(new_n553), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n348), .B(new_n1030), .C1(G68), .C2(new_n750), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n797), .A2(new_n249), .B1(new_n915), .B2(new_n737), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT51), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1029), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n719), .A2(new_n476), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n797), .A2(new_n901), .B1(new_n798), .B2(new_n737), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT52), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n809), .A2(new_n796), .B1(new_n723), .B2(new_n899), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(G107), .A2(new_n752), .B1(new_n741), .B2(G322), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n278), .B1(new_n731), .B2(G116), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1037), .A2(new_n1039), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1034), .B1(new_n1035), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n761), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1024), .A2(new_n774), .A3(new_n1025), .A4(new_n1044), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1022), .A2(new_n1023), .A3(new_n1045), .ZN(G390));
  INV_X1    g0846(.A(KEYINPUT116), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n696), .A2(G330), .A3(new_n787), .A4(new_n845), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n868), .A2(new_n869), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n876), .B2(new_n871), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n655), .B1(new_n708), .B2(new_n710), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n875), .B1(new_n1051), .B2(new_n788), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n845), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n871), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1053), .A2(new_n860), .A3(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1048), .B1(new_n1050), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1050), .A2(new_n1055), .A3(new_n1048), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1047), .B1(new_n1059), .B2(new_n772), .ZN(new_n1060));
  AND3_X1   g0860(.A1(new_n1050), .A2(new_n1048), .A3(new_n1055), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1061), .A2(new_n1056), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1062), .A2(KEYINPUT116), .A3(new_n773), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n591), .A2(G330), .A3(new_n696), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n638), .A2(new_n879), .A3(new_n1065), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n787), .B(G330), .C1(new_n676), .C2(new_n695), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n873), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n1048), .A2(new_n1068), .B1(new_n790), .B2(new_n875), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT115), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1048), .A2(new_n1068), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n1069), .A2(new_n1070), .B1(new_n1071), .B2(new_n1052), .ZN(new_n1072));
  OR3_X1    g0872(.A1(new_n1071), .A2(new_n1070), .A3(new_n1052), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1066), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n1059), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1074), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1076), .A2(new_n1077), .A3(new_n669), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n723), .A2(new_n249), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT53), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n741), .A2(G125), .ZN(new_n1081));
  INV_X1    g0881(.A(G132), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1080), .B(new_n1081), .C1(new_n1082), .C2(new_n737), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n743), .A2(G128), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(KEYINPUT54), .B(G143), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT117), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1087), .A2(new_n719), .ZN(new_n1088));
  NOR4_X1   g0888(.A1(new_n1083), .A2(new_n348), .A3(new_n1084), .A4(new_n1088), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n1089), .B1(new_n202), .B2(new_n728), .C1(new_n915), .C2(new_n732), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(G137), .B2(new_n734), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT118), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n809), .A2(new_n307), .B1(new_n443), .B2(new_n719), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT119), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n797), .A2(new_n726), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n1026), .B(new_n1095), .C1(G87), .C2(new_n724), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n348), .B1(new_n740), .B2(new_n476), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n812), .B(new_n1097), .C1(new_n738), .C2(G116), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1094), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1092), .A2(new_n1099), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT120), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n761), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1049), .A2(new_n762), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n818), .A2(new_n255), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1102), .A2(new_n1103), .A3(new_n774), .A4(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1064), .A2(new_n1078), .A3(new_n1105), .ZN(G378));
  NAND2_X1  g0906(.A1(new_n1066), .A2(KEYINPUT123), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT123), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n638), .A2(new_n879), .A3(new_n1108), .A4(new_n1065), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1077), .A2(new_n1111), .ZN(new_n1112));
  AND3_X1   g0912(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n856), .B1(new_n855), .B2(new_n857), .ZN(new_n1114));
  OAI211_X1 g0914(.A(G330), .B(new_n861), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n298), .A2(new_n303), .ZN(new_n1116));
  NOR3_X1   g0916(.A1(new_n269), .A2(new_n270), .A3(new_n645), .ZN(new_n1117));
  OR2_X1    g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1118), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1115), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n859), .A2(G330), .A3(new_n861), .A4(new_n1125), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n1127), .A2(new_n1128), .A3(new_n878), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n878), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1112), .B(KEYINPUT57), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT122), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(new_n872), .B2(new_n877), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n1127), .A2(new_n1128), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1110), .B1(new_n1062), .B2(new_n1074), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1133), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1136));
  NOR3_X1   g0936(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n669), .B(new_n1131), .C1(new_n1137), .C2(KEYINPUT57), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1126), .A2(new_n762), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n202), .B1(new_n346), .B2(G41), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n719), .A2(new_n808), .B1(new_n249), .B2(new_n732), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(G125), .A2(new_n743), .B1(new_n1086), .B2(new_n750), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n1082), .B2(new_n809), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n1141), .B(new_n1143), .C1(G128), .C2(new_n738), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT59), .ZN(new_n1145));
  OR2_X1    g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n752), .A2(G159), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(KEYINPUT121), .B(G124), .ZN(new_n1148));
  AOI21_X1  g0948(.A(G41), .B1(new_n741), .B2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1146), .A2(new_n252), .A3(new_n1147), .A4(new_n1149), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1140), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n728), .A2(new_n340), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n720), .A2(new_n562), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n743), .A2(G116), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(G77), .A2(new_n750), .B1(new_n741), .B2(G283), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1154), .A2(new_n1155), .A3(new_n914), .A4(new_n1156), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1153), .B(new_n1157), .C1(G107), .C2(new_n738), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n734), .A2(G97), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1158), .A2(new_n283), .A3(new_n348), .A4(new_n1159), .ZN(new_n1160));
  XOR2_X1   g0960(.A(new_n1160), .B(KEYINPUT58), .Z(new_n1161));
  OAI21_X1  g0961(.A(new_n761), .B1(new_n1152), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n818), .A2(new_n202), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1139), .A2(new_n774), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1165), .B1(new_n1166), .B2(new_n773), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1138), .A2(new_n1167), .ZN(G375));
  NAND2_X1  g0968(.A1(new_n873), .A2(new_n762), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1153), .B1(G50), .B2(new_n731), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n348), .B1(new_n743), .B2(G132), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n724), .A2(G159), .B1(G128), .B2(new_n741), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1170), .B(new_n1171), .C1(new_n1172), .C2(KEYINPUT124), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1172), .A2(KEYINPUT124), .B1(G137), .B2(new_n738), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n809), .B2(new_n1087), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1173), .B(new_n1175), .C1(G150), .C2(new_n720), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n724), .A2(G97), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n734), .A2(G116), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n278), .B1(new_n741), .B2(G303), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1177), .A2(new_n1009), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n797), .A2(new_n476), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n719), .A2(new_n307), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n737), .A2(new_n726), .B1(new_n211), .B2(new_n728), .ZN(new_n1183));
  NOR4_X1   g0983(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n761), .B1(new_n1176), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n818), .A2(new_n221), .ZN(new_n1186));
  AND4_X1   g0986(.A1(new_n774), .A2(new_n1169), .A3(new_n1185), .A4(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1187), .B1(new_n1188), .B2(new_n773), .ZN(new_n1189));
  AND3_X1   g0989(.A1(new_n1072), .A2(new_n1073), .A3(new_n1066), .ZN(new_n1190));
  OR2_X1    g0990(.A1(new_n1190), .A2(new_n964), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1189), .B1(new_n1191), .B2(new_n1074), .ZN(G381));
  NOR4_X1   g0992(.A1(G375), .A2(G384), .A3(G378), .A4(G381), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n967), .A2(new_n932), .A3(new_n978), .ZN(new_n1194));
  OAI21_X1  g0994(.A(KEYINPUT107), .B1(new_n980), .B2(new_n977), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(G390), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1196), .A2(new_n931), .A3(new_n1197), .ZN(new_n1198));
  NOR3_X1   g0998(.A1(new_n1198), .A2(G396), .A3(G393), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1193), .A2(new_n1199), .ZN(G407));
  INV_X1    g1000(.A(G378), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1138), .A2(new_n1201), .A3(new_n646), .A4(new_n1167), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(G407), .A2(G213), .A3(new_n1202), .ZN(G409));
  XOR2_X1   g1003(.A(G393), .B(G396), .Z(new_n1204));
  AOI21_X1  g1004(.A(new_n1197), .B1(new_n1196), .B2(new_n931), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n930), .B(G390), .C1(new_n1194), .C2(new_n1195), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1204), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(G387), .A2(G390), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1204), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1208), .A2(new_n1198), .A3(new_n1209), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n1207), .A2(new_n1210), .A3(KEYINPUT127), .ZN(new_n1211));
  AOI21_X1  g1011(.A(KEYINPUT127), .B1(new_n1207), .B2(new_n1210), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1138), .A2(G378), .A3(new_n1167), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1166), .A2(new_n933), .A3(new_n1112), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n773), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1215), .A2(new_n1164), .A3(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n1201), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1214), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n646), .A2(G213), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1190), .A2(KEYINPUT60), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1221), .A2(new_n669), .A3(new_n1075), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1190), .A2(KEYINPUT60), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1189), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1224), .B(G384), .ZN(new_n1225));
  AND4_X1   g1025(.A1(KEYINPUT62), .A2(new_n1219), .A3(new_n1220), .A4(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT125), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1219), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1214), .A2(new_n1218), .A3(KEYINPUT125), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1228), .A2(new_n1220), .A3(new_n1225), .A4(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT62), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1226), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT61), .ZN(new_n1233));
  AND2_X1   g1033(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n646), .A2(G213), .A3(G2897), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1225), .B(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1233), .B1(new_n1234), .B2(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1213), .B1(new_n1232), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT63), .ZN(new_n1239));
  AOI21_X1  g1039(.A(KEYINPUT61), .B1(new_n1230), .B2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1228), .A2(new_n1220), .A3(new_n1229), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1236), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1207), .A2(new_n1210), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT126), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1219), .A2(KEYINPUT63), .A3(new_n1220), .A4(new_n1225), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1244), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  OR2_X1    g1047(.A1(new_n1246), .A2(new_n1245), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1240), .A2(new_n1243), .A3(new_n1247), .A4(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1238), .A2(new_n1249), .ZN(G405));
  XNOR2_X1  g1050(.A(G375), .B(G378), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n1251), .A2(new_n1225), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1251), .A2(new_n1225), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n1213), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n1252), .A2(new_n1253), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(G402));
endmodule


