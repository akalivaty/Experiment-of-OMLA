

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U560 ( .A(KEYINPUT101), .ZN(n697) );
  INV_X1 U561 ( .A(KEYINPUT31), .ZN(n706) );
  NAND2_X1 U562 ( .A1(n769), .A2(n771), .ZN(n743) );
  NAND2_X1 U563 ( .A1(G8), .A2(n743), .ZN(n825) );
  NOR2_X1 U564 ( .A1(G651), .A2(n656), .ZN(n650) );
  XOR2_X1 U565 ( .A(KEYINPUT0), .B(G543), .Z(n656) );
  INV_X1 U566 ( .A(G651), .ZN(n529) );
  NOR2_X1 U567 ( .A1(n656), .A2(n529), .ZN(n644) );
  NAND2_X1 U568 ( .A1(G72), .A2(n644), .ZN(n528) );
  NOR2_X1 U569 ( .A1(G651), .A2(G543), .ZN(n641) );
  NAND2_X1 U570 ( .A1(G85), .A2(n641), .ZN(n527) );
  NAND2_X1 U571 ( .A1(n528), .A2(n527), .ZN(n536) );
  NAND2_X1 U572 ( .A1(n650), .A2(G47), .ZN(n534) );
  NOR2_X1 U573 ( .A1(G543), .A2(n529), .ZN(n531) );
  XNOR2_X1 U574 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n530) );
  XNOR2_X1 U575 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U576 ( .A(KEYINPUT65), .B(n532), .ZN(n654) );
  NAND2_X1 U577 ( .A1(G60), .A2(n654), .ZN(n533) );
  NAND2_X1 U578 ( .A1(n534), .A2(n533), .ZN(n535) );
  OR2_X1 U579 ( .A1(n536), .A2(n535), .ZN(G290) );
  NOR2_X1 U580 ( .A1(G2105), .A2(G2104), .ZN(n537) );
  XOR2_X2 U581 ( .A(KEYINPUT17), .B(n537), .Z(n895) );
  NAND2_X1 U582 ( .A1(G137), .A2(n895), .ZN(n539) );
  AND2_X1 U583 ( .A1(G2105), .A2(G2104), .ZN(n901) );
  NAND2_X1 U584 ( .A1(G113), .A2(n901), .ZN(n538) );
  NAND2_X1 U585 ( .A1(n539), .A2(n538), .ZN(n541) );
  INV_X1 U586 ( .A(KEYINPUT64), .ZN(n540) );
  XNOR2_X1 U587 ( .A(n541), .B(n540), .ZN(n543) );
  INV_X1 U588 ( .A(G2105), .ZN(n544) );
  NOR2_X1 U589 ( .A1(G2104), .A2(n544), .ZN(n900) );
  NAND2_X1 U590 ( .A1(n900), .A2(G125), .ZN(n542) );
  AND2_X1 U591 ( .A1(n543), .A2(n542), .ZN(n691) );
  AND2_X1 U592 ( .A1(n544), .A2(G2104), .ZN(n896) );
  NAND2_X1 U593 ( .A1(G101), .A2(n896), .ZN(n545) );
  XOR2_X1 U594 ( .A(KEYINPUT23), .B(n545), .Z(n689) );
  AND2_X1 U595 ( .A1(n691), .A2(n689), .ZN(n688) );
  BUF_X1 U596 ( .A(n688), .Z(G160) );
  NAND2_X1 U597 ( .A1(n650), .A2(G52), .ZN(n547) );
  NAND2_X1 U598 ( .A1(G64), .A2(n654), .ZN(n546) );
  NAND2_X1 U599 ( .A1(n547), .A2(n546), .ZN(n553) );
  NAND2_X1 U600 ( .A1(n641), .A2(G90), .ZN(n548) );
  XOR2_X1 U601 ( .A(KEYINPUT67), .B(n548), .Z(n550) );
  NAND2_X1 U602 ( .A1(n644), .A2(G77), .ZN(n549) );
  NAND2_X1 U603 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U604 ( .A(KEYINPUT9), .B(n551), .Z(n552) );
  NOR2_X1 U605 ( .A1(n553), .A2(n552), .ZN(G171) );
  AND2_X1 U606 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U607 ( .A(G57), .ZN(G237) );
  INV_X1 U608 ( .A(G69), .ZN(G235) );
  INV_X1 U609 ( .A(G108), .ZN(G238) );
  INV_X1 U610 ( .A(G120), .ZN(G236) );
  INV_X1 U611 ( .A(G82), .ZN(G220) );
  NAND2_X1 U612 ( .A1(G126), .A2(n900), .ZN(n555) );
  NAND2_X1 U613 ( .A1(G138), .A2(n895), .ZN(n554) );
  NAND2_X1 U614 ( .A1(n555), .A2(n554), .ZN(n559) );
  NAND2_X1 U615 ( .A1(G114), .A2(n901), .ZN(n557) );
  NAND2_X1 U616 ( .A1(G102), .A2(n896), .ZN(n556) );
  NAND2_X1 U617 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U618 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U619 ( .A(KEYINPUT88), .B(n560), .ZN(G164) );
  NAND2_X1 U620 ( .A1(G7), .A2(G661), .ZN(n561) );
  XNOR2_X1 U621 ( .A(n561), .B(KEYINPUT10), .ZN(n562) );
  XNOR2_X1 U622 ( .A(KEYINPUT70), .B(n562), .ZN(G223) );
  XOR2_X1 U623 ( .A(KEYINPUT72), .B(KEYINPUT11), .Z(n564) );
  XNOR2_X1 U624 ( .A(KEYINPUT71), .B(G223), .ZN(n851) );
  NAND2_X1 U625 ( .A1(n851), .A2(G567), .ZN(n563) );
  XNOR2_X1 U626 ( .A(n564), .B(n563), .ZN(G234) );
  NAND2_X1 U627 ( .A1(n650), .A2(G43), .ZN(n565) );
  XNOR2_X1 U628 ( .A(KEYINPUT75), .B(n565), .ZN(n576) );
  NAND2_X1 U629 ( .A1(G56), .A2(n654), .ZN(n566) );
  XOR2_X1 U630 ( .A(KEYINPUT14), .B(n566), .Z(n573) );
  NAND2_X1 U631 ( .A1(n644), .A2(G68), .ZN(n567) );
  XNOR2_X1 U632 ( .A(KEYINPUT73), .B(n567), .ZN(n570) );
  NAND2_X1 U633 ( .A1(n641), .A2(G81), .ZN(n568) );
  XOR2_X1 U634 ( .A(KEYINPUT12), .B(n568), .Z(n569) );
  NOR2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n571), .B(KEYINPUT13), .ZN(n572) );
  NOR2_X1 U637 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U638 ( .A(KEYINPUT74), .B(n574), .Z(n575) );
  NOR2_X1 U639 ( .A1(n576), .A2(n575), .ZN(n1018) );
  NAND2_X1 U640 ( .A1(G860), .A2(n1018), .ZN(n577) );
  XNOR2_X1 U641 ( .A(n577), .B(KEYINPUT76), .ZN(G153) );
  INV_X1 U642 ( .A(G171), .ZN(G301) );
  NAND2_X1 U643 ( .A1(n650), .A2(G54), .ZN(n579) );
  NAND2_X1 U644 ( .A1(G66), .A2(n654), .ZN(n578) );
  NAND2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n583) );
  NAND2_X1 U646 ( .A1(G79), .A2(n644), .ZN(n581) );
  NAND2_X1 U647 ( .A1(G92), .A2(n641), .ZN(n580) );
  NAND2_X1 U648 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U649 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n584), .B(KEYINPUT15), .ZN(n1042) );
  INV_X1 U651 ( .A(n1042), .ZN(n919) );
  NOR2_X1 U652 ( .A1(n919), .A2(G868), .ZN(n585) );
  XNOR2_X1 U653 ( .A(n585), .B(KEYINPUT77), .ZN(n587) );
  NAND2_X1 U654 ( .A1(G868), .A2(G301), .ZN(n586) );
  NAND2_X1 U655 ( .A1(n587), .A2(n586), .ZN(G284) );
  NAND2_X1 U656 ( .A1(n650), .A2(G51), .ZN(n589) );
  NAND2_X1 U657 ( .A1(G63), .A2(n654), .ZN(n588) );
  NAND2_X1 U658 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U659 ( .A(KEYINPUT6), .B(n590), .ZN(n596) );
  NAND2_X1 U660 ( .A1(n641), .A2(G89), .ZN(n591) );
  XNOR2_X1 U661 ( .A(n591), .B(KEYINPUT4), .ZN(n593) );
  NAND2_X1 U662 ( .A1(G76), .A2(n644), .ZN(n592) );
  NAND2_X1 U663 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U664 ( .A(n594), .B(KEYINPUT5), .Z(n595) );
  NOR2_X1 U665 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U666 ( .A(KEYINPUT7), .B(n597), .Z(n598) );
  XNOR2_X1 U667 ( .A(KEYINPUT78), .B(n598), .ZN(G168) );
  XOR2_X1 U668 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U669 ( .A1(G91), .A2(n641), .ZN(n600) );
  NAND2_X1 U670 ( .A1(G65), .A2(n654), .ZN(n599) );
  NAND2_X1 U671 ( .A1(n600), .A2(n599), .ZN(n603) );
  NAND2_X1 U672 ( .A1(n644), .A2(G78), .ZN(n601) );
  XOR2_X1 U673 ( .A(KEYINPUT68), .B(n601), .Z(n602) );
  NOR2_X1 U674 ( .A1(n603), .A2(n602), .ZN(n605) );
  NAND2_X1 U675 ( .A1(n650), .A2(G53), .ZN(n604) );
  NAND2_X1 U676 ( .A1(n605), .A2(n604), .ZN(G299) );
  INV_X1 U677 ( .A(G868), .ZN(n668) );
  NOR2_X1 U678 ( .A1(G286), .A2(n668), .ZN(n606) );
  XOR2_X1 U679 ( .A(KEYINPUT79), .B(n606), .Z(n608) );
  NOR2_X1 U680 ( .A1(G868), .A2(G299), .ZN(n607) );
  NOR2_X1 U681 ( .A1(n608), .A2(n607), .ZN(G297) );
  INV_X1 U682 ( .A(G860), .ZN(n609) );
  NAND2_X1 U683 ( .A1(n609), .A2(G559), .ZN(n610) );
  NAND2_X1 U684 ( .A1(n610), .A2(n919), .ZN(n611) );
  XNOR2_X1 U685 ( .A(n611), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U686 ( .A1(n919), .A2(G868), .ZN(n612) );
  NOR2_X1 U687 ( .A1(G559), .A2(n612), .ZN(n614) );
  AND2_X1 U688 ( .A1(n668), .A2(n1018), .ZN(n613) );
  NOR2_X1 U689 ( .A1(n614), .A2(n613), .ZN(G282) );
  XOR2_X1 U690 ( .A(G2100), .B(KEYINPUT80), .Z(n623) );
  NAND2_X1 U691 ( .A1(n900), .A2(G123), .ZN(n615) );
  XNOR2_X1 U692 ( .A(n615), .B(KEYINPUT18), .ZN(n617) );
  NAND2_X1 U693 ( .A1(G111), .A2(n901), .ZN(n616) );
  NAND2_X1 U694 ( .A1(n617), .A2(n616), .ZN(n621) );
  NAND2_X1 U695 ( .A1(G135), .A2(n895), .ZN(n619) );
  NAND2_X1 U696 ( .A1(G99), .A2(n896), .ZN(n618) );
  NAND2_X1 U697 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U698 ( .A1(n621), .A2(n620), .ZN(n1002) );
  XNOR2_X1 U699 ( .A(G2096), .B(n1002), .ZN(n622) );
  NAND2_X1 U700 ( .A1(n623), .A2(n622), .ZN(G156) );
  NAND2_X1 U701 ( .A1(G80), .A2(n644), .ZN(n625) );
  NAND2_X1 U702 ( .A1(G93), .A2(n641), .ZN(n624) );
  NAND2_X1 U703 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U704 ( .A(KEYINPUT81), .B(n626), .ZN(n631) );
  NAND2_X1 U705 ( .A1(n650), .A2(G55), .ZN(n628) );
  NAND2_X1 U706 ( .A1(G67), .A2(n654), .ZN(n627) );
  NAND2_X1 U707 ( .A1(n628), .A2(n627), .ZN(n629) );
  XOR2_X1 U708 ( .A(KEYINPUT82), .B(n629), .Z(n630) );
  NAND2_X1 U709 ( .A1(n631), .A2(n630), .ZN(n667) );
  NAND2_X1 U710 ( .A1(G559), .A2(n919), .ZN(n632) );
  XOR2_X1 U711 ( .A(n1018), .B(n632), .Z(n664) );
  NOR2_X1 U712 ( .A1(n664), .A2(G860), .ZN(n633) );
  XNOR2_X1 U713 ( .A(n633), .B(KEYINPUT83), .ZN(n634) );
  XNOR2_X1 U714 ( .A(n667), .B(n634), .ZN(G145) );
  NAND2_X1 U715 ( .A1(G75), .A2(n644), .ZN(n636) );
  NAND2_X1 U716 ( .A1(G88), .A2(n641), .ZN(n635) );
  NAND2_X1 U717 ( .A1(n636), .A2(n635), .ZN(n640) );
  NAND2_X1 U718 ( .A1(n650), .A2(G50), .ZN(n638) );
  NAND2_X1 U719 ( .A1(G62), .A2(n654), .ZN(n637) );
  NAND2_X1 U720 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U721 ( .A1(n640), .A2(n639), .ZN(G166) );
  NAND2_X1 U722 ( .A1(G86), .A2(n641), .ZN(n643) );
  NAND2_X1 U723 ( .A1(G61), .A2(n654), .ZN(n642) );
  NAND2_X1 U724 ( .A1(n643), .A2(n642), .ZN(n647) );
  NAND2_X1 U725 ( .A1(n644), .A2(G73), .ZN(n645) );
  XOR2_X1 U726 ( .A(KEYINPUT2), .B(n645), .Z(n646) );
  NOR2_X1 U727 ( .A1(n647), .A2(n646), .ZN(n649) );
  NAND2_X1 U728 ( .A1(n650), .A2(G48), .ZN(n648) );
  NAND2_X1 U729 ( .A1(n649), .A2(n648), .ZN(G305) );
  NAND2_X1 U730 ( .A1(G49), .A2(n650), .ZN(n652) );
  NAND2_X1 U731 ( .A1(G74), .A2(G651), .ZN(n651) );
  NAND2_X1 U732 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U733 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U734 ( .A(n655), .B(KEYINPUT84), .ZN(n658) );
  NAND2_X1 U735 ( .A1(G87), .A2(n656), .ZN(n657) );
  NAND2_X1 U736 ( .A1(n658), .A2(n657), .ZN(G288) );
  XNOR2_X1 U737 ( .A(G166), .B(G305), .ZN(n659) );
  XNOR2_X1 U738 ( .A(n659), .B(n667), .ZN(n660) );
  XNOR2_X1 U739 ( .A(KEYINPUT19), .B(n660), .ZN(n662) );
  INV_X1 U740 ( .A(G299), .ZN(n1038) );
  XNOR2_X1 U741 ( .A(G290), .B(n1038), .ZN(n661) );
  XNOR2_X1 U742 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U743 ( .A(n663), .B(G288), .ZN(n918) );
  XNOR2_X1 U744 ( .A(KEYINPUT85), .B(n664), .ZN(n665) );
  XNOR2_X1 U745 ( .A(n918), .B(n665), .ZN(n666) );
  NAND2_X1 U746 ( .A1(n666), .A2(G868), .ZN(n670) );
  NAND2_X1 U747 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U748 ( .A1(n670), .A2(n669), .ZN(G295) );
  NAND2_X1 U749 ( .A1(G2078), .A2(G2084), .ZN(n671) );
  XOR2_X1 U750 ( .A(KEYINPUT20), .B(n671), .Z(n672) );
  NAND2_X1 U751 ( .A1(G2090), .A2(n672), .ZN(n673) );
  XNOR2_X1 U752 ( .A(KEYINPUT21), .B(n673), .ZN(n674) );
  NAND2_X1 U753 ( .A1(n674), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U754 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U755 ( .A(KEYINPUT69), .B(G132), .ZN(G219) );
  NOR2_X1 U756 ( .A1(G220), .A2(G219), .ZN(n675) );
  XOR2_X1 U757 ( .A(KEYINPUT22), .B(n675), .Z(n676) );
  NOR2_X1 U758 ( .A1(G218), .A2(n676), .ZN(n677) );
  NAND2_X1 U759 ( .A1(G96), .A2(n677), .ZN(n855) );
  NAND2_X1 U760 ( .A1(G2106), .A2(n855), .ZN(n678) );
  XOR2_X1 U761 ( .A(KEYINPUT86), .B(n678), .Z(n683) );
  NOR2_X1 U762 ( .A1(G236), .A2(G238), .ZN(n680) );
  NOR2_X1 U763 ( .A1(G235), .A2(G237), .ZN(n679) );
  NAND2_X1 U764 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U765 ( .A(KEYINPUT87), .B(n681), .Z(n856) );
  AND2_X1 U766 ( .A1(n856), .A2(G567), .ZN(n682) );
  NOR2_X1 U767 ( .A1(n683), .A2(n682), .ZN(G319) );
  INV_X1 U768 ( .A(G319), .ZN(n685) );
  NAND2_X1 U769 ( .A1(G483), .A2(G661), .ZN(n684) );
  NOR2_X1 U770 ( .A1(n685), .A2(n684), .ZN(n854) );
  NAND2_X1 U771 ( .A1(n854), .A2(G36), .ZN(G176) );
  INV_X1 U772 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U773 ( .A(KEYINPUT40), .B(KEYINPUT110), .ZN(n850) );
  AND2_X1 U774 ( .A1(G288), .A2(G1976), .ZN(n1027) );
  INV_X1 U775 ( .A(n1027), .ZN(n757) );
  INV_X1 U776 ( .A(KEYINPUT89), .ZN(n686) );
  AND2_X1 U777 ( .A1(G40), .A2(n686), .ZN(n687) );
  NAND2_X1 U778 ( .A1(n688), .A2(n687), .ZN(n694) );
  AND2_X1 U779 ( .A1(G40), .A2(n689), .ZN(n690) );
  NAND2_X1 U780 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U781 ( .A1(KEYINPUT89), .A2(n692), .ZN(n693) );
  NAND2_X1 U782 ( .A1(n694), .A2(n693), .ZN(n769) );
  NOR2_X1 U783 ( .A1(G1384), .A2(G164), .ZN(n771) );
  NOR2_X1 U784 ( .A1(G2084), .A2(n743), .ZN(n696) );
  NAND2_X1 U785 ( .A1(G8), .A2(n696), .ZN(n741) );
  NOR2_X1 U786 ( .A1(G1966), .A2(n825), .ZN(n695) );
  XOR2_X1 U787 ( .A(KEYINPUT97), .B(n695), .Z(n739) );
  NOR2_X1 U788 ( .A1(n739), .A2(n696), .ZN(n698) );
  XNOR2_X1 U789 ( .A(n698), .B(n697), .ZN(n699) );
  NAND2_X1 U790 ( .A1(n699), .A2(G8), .ZN(n700) );
  XNOR2_X1 U791 ( .A(KEYINPUT30), .B(n700), .ZN(n701) );
  NOR2_X1 U792 ( .A1(G168), .A2(n701), .ZN(n705) );
  INV_X1 U793 ( .A(G1961), .ZN(n967) );
  NAND2_X1 U794 ( .A1(n743), .A2(n967), .ZN(n703) );
  AND2_X1 U795 ( .A1(n771), .A2(n769), .ZN(n720) );
  XNOR2_X1 U796 ( .A(G2078), .B(KEYINPUT25), .ZN(n941) );
  NAND2_X1 U797 ( .A1(n720), .A2(n941), .ZN(n702) );
  NAND2_X1 U798 ( .A1(n703), .A2(n702), .ZN(n708) );
  NOR2_X1 U799 ( .A1(G171), .A2(n708), .ZN(n704) );
  NOR2_X1 U800 ( .A1(n705), .A2(n704), .ZN(n707) );
  XNOR2_X1 U801 ( .A(n707), .B(n706), .ZN(n737) );
  NAND2_X1 U802 ( .A1(n708), .A2(G171), .ZN(n735) );
  NAND2_X1 U803 ( .A1(n720), .A2(G2072), .ZN(n709) );
  XNOR2_X1 U804 ( .A(KEYINPUT27), .B(n709), .ZN(n712) );
  NAND2_X1 U805 ( .A1(G1956), .A2(n743), .ZN(n710) );
  XOR2_X1 U806 ( .A(KEYINPUT98), .B(n710), .Z(n711) );
  NOR2_X1 U807 ( .A1(n712), .A2(n711), .ZN(n715) );
  NOR2_X1 U808 ( .A1(n1038), .A2(n715), .ZN(n714) );
  XNOR2_X1 U809 ( .A(KEYINPUT99), .B(KEYINPUT28), .ZN(n713) );
  XNOR2_X1 U810 ( .A(n714), .B(n713), .ZN(n732) );
  NAND2_X1 U811 ( .A1(n1038), .A2(n715), .ZN(n730) );
  AND2_X1 U812 ( .A1(n720), .A2(G1996), .ZN(n717) );
  XOR2_X1 U813 ( .A(KEYINPUT26), .B(KEYINPUT100), .Z(n716) );
  XNOR2_X1 U814 ( .A(n717), .B(n716), .ZN(n719) );
  NAND2_X1 U815 ( .A1(n743), .A2(G1341), .ZN(n718) );
  NAND2_X1 U816 ( .A1(n719), .A2(n718), .ZN(n725) );
  NAND2_X1 U817 ( .A1(G1348), .A2(n743), .ZN(n722) );
  NAND2_X1 U818 ( .A1(G2067), .A2(n720), .ZN(n721) );
  NAND2_X1 U819 ( .A1(n722), .A2(n721), .ZN(n726) );
  NAND2_X1 U820 ( .A1(n1042), .A2(n726), .ZN(n723) );
  NAND2_X1 U821 ( .A1(n1018), .A2(n723), .ZN(n724) );
  NOR2_X1 U822 ( .A1(n725), .A2(n724), .ZN(n728) );
  NOR2_X1 U823 ( .A1(n726), .A2(n1042), .ZN(n727) );
  NOR2_X1 U824 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U825 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U826 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U827 ( .A(KEYINPUT29), .B(n733), .Z(n734) );
  NAND2_X1 U828 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U829 ( .A1(n737), .A2(n736), .ZN(n742) );
  INV_X1 U830 ( .A(n742), .ZN(n738) );
  NOR2_X1 U831 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U832 ( .A1(n741), .A2(n740), .ZN(n754) );
  NAND2_X1 U833 ( .A1(G286), .A2(n742), .ZN(n750) );
  NOR2_X1 U834 ( .A1(G2090), .A2(n743), .ZN(n744) );
  XOR2_X1 U835 ( .A(KEYINPUT103), .B(n744), .Z(n747) );
  NOR2_X1 U836 ( .A1(G1971), .A2(n825), .ZN(n745) );
  XNOR2_X1 U837 ( .A(KEYINPUT102), .B(n745), .ZN(n746) );
  NOR2_X1 U838 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U839 ( .A1(n748), .A2(G303), .ZN(n749) );
  NAND2_X1 U840 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U841 ( .A1(n751), .A2(G8), .ZN(n752) );
  XNOR2_X1 U842 ( .A(n752), .B(KEYINPUT32), .ZN(n753) );
  NAND2_X1 U843 ( .A1(n754), .A2(n753), .ZN(n819) );
  NOR2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n755) );
  XOR2_X1 U845 ( .A(KEYINPUT104), .B(n755), .Z(n1045) );
  INV_X1 U846 ( .A(n1045), .ZN(n807) );
  NOR2_X1 U847 ( .A1(G1971), .A2(G303), .ZN(n1039) );
  NOR2_X1 U848 ( .A1(n807), .A2(n1039), .ZN(n756) );
  NAND2_X1 U849 ( .A1(n819), .A2(n756), .ZN(n806) );
  AND2_X1 U850 ( .A1(n757), .A2(n806), .ZN(n794) );
  INV_X1 U851 ( .A(n825), .ZN(n802) );
  NAND2_X1 U852 ( .A1(G140), .A2(n895), .ZN(n759) );
  NAND2_X1 U853 ( .A1(G104), .A2(n896), .ZN(n758) );
  NAND2_X1 U854 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U855 ( .A(KEYINPUT34), .B(n760), .ZN(n766) );
  NAND2_X1 U856 ( .A1(n900), .A2(G128), .ZN(n761) );
  XNOR2_X1 U857 ( .A(n761), .B(KEYINPUT90), .ZN(n763) );
  NAND2_X1 U858 ( .A1(G116), .A2(n901), .ZN(n762) );
  NAND2_X1 U859 ( .A1(n763), .A2(n762), .ZN(n764) );
  XOR2_X1 U860 ( .A(n764), .B(KEYINPUT35), .Z(n765) );
  NOR2_X1 U861 ( .A1(n766), .A2(n765), .ZN(n767) );
  XOR2_X1 U862 ( .A(KEYINPUT36), .B(n767), .Z(n768) );
  XNOR2_X1 U863 ( .A(KEYINPUT91), .B(n768), .ZN(n915) );
  XNOR2_X1 U864 ( .A(G2067), .B(KEYINPUT37), .ZN(n843) );
  NOR2_X1 U865 ( .A1(n915), .A2(n843), .ZN(n999) );
  INV_X1 U866 ( .A(n769), .ZN(n770) );
  NOR2_X1 U867 ( .A1(n771), .A2(n770), .ZN(n845) );
  NAND2_X1 U868 ( .A1(n999), .A2(n845), .ZN(n772) );
  XNOR2_X1 U869 ( .A(n772), .B(KEYINPUT92), .ZN(n841) );
  NAND2_X1 U870 ( .A1(n895), .A2(G131), .ZN(n773) );
  XOR2_X1 U871 ( .A(KEYINPUT93), .B(n773), .Z(n775) );
  NAND2_X1 U872 ( .A1(n896), .A2(G95), .ZN(n774) );
  NAND2_X1 U873 ( .A1(n775), .A2(n774), .ZN(n776) );
  XOR2_X1 U874 ( .A(KEYINPUT94), .B(n776), .Z(n780) );
  NAND2_X1 U875 ( .A1(G119), .A2(n900), .ZN(n778) );
  NAND2_X1 U876 ( .A1(G107), .A2(n901), .ZN(n777) );
  AND2_X1 U877 ( .A1(n778), .A2(n777), .ZN(n779) );
  NAND2_X1 U878 ( .A1(n780), .A2(n779), .ZN(n911) );
  NAND2_X1 U879 ( .A1(G1991), .A2(n911), .ZN(n781) );
  XOR2_X1 U880 ( .A(KEYINPUT95), .B(n781), .Z(n790) );
  NAND2_X1 U881 ( .A1(G129), .A2(n900), .ZN(n783) );
  NAND2_X1 U882 ( .A1(G141), .A2(n895), .ZN(n782) );
  NAND2_X1 U883 ( .A1(n783), .A2(n782), .ZN(n786) );
  NAND2_X1 U884 ( .A1(n896), .A2(G105), .ZN(n784) );
  XOR2_X1 U885 ( .A(KEYINPUT38), .B(n784), .Z(n785) );
  NOR2_X1 U886 ( .A1(n786), .A2(n785), .ZN(n788) );
  NAND2_X1 U887 ( .A1(n901), .A2(G117), .ZN(n787) );
  NAND2_X1 U888 ( .A1(n788), .A2(n787), .ZN(n907) );
  NAND2_X1 U889 ( .A1(G1996), .A2(n907), .ZN(n789) );
  NAND2_X1 U890 ( .A1(n790), .A2(n789), .ZN(n1010) );
  NAND2_X1 U891 ( .A1(n1010), .A2(n845), .ZN(n791) );
  XOR2_X1 U892 ( .A(KEYINPUT96), .B(n791), .Z(n837) );
  INV_X1 U893 ( .A(n837), .ZN(n792) );
  NAND2_X1 U894 ( .A1(n841), .A2(n792), .ZN(n796) );
  INV_X1 U895 ( .A(n796), .ZN(n827) );
  AND2_X1 U896 ( .A1(n802), .A2(n827), .ZN(n793) );
  NAND2_X1 U897 ( .A1(n794), .A2(n793), .ZN(n798) );
  NOR2_X1 U898 ( .A1(KEYINPUT105), .A2(KEYINPUT33), .ZN(n795) );
  OR2_X1 U899 ( .A1(n796), .A2(n795), .ZN(n797) );
  NAND2_X1 U900 ( .A1(n798), .A2(n797), .ZN(n816) );
  INV_X1 U901 ( .A(KEYINPUT105), .ZN(n799) );
  OR2_X1 U902 ( .A1(n799), .A2(n1027), .ZN(n804) );
  XNOR2_X1 U903 ( .A(G1981), .B(G305), .ZN(n1031) );
  INV_X1 U904 ( .A(n1031), .ZN(n801) );
  NAND2_X1 U905 ( .A1(KEYINPUT105), .A2(KEYINPUT33), .ZN(n800) );
  AND2_X1 U906 ( .A1(n801), .A2(n800), .ZN(n809) );
  INV_X1 U907 ( .A(n809), .ZN(n803) );
  NOR2_X1 U908 ( .A1(n803), .A2(n802), .ZN(n812) );
  NOR2_X1 U909 ( .A1(n804), .A2(n812), .ZN(n805) );
  NAND2_X1 U910 ( .A1(n806), .A2(n805), .ZN(n814) );
  NAND2_X1 U911 ( .A1(KEYINPUT33), .A2(n807), .ZN(n808) );
  XNOR2_X1 U912 ( .A(n808), .B(KEYINPUT106), .ZN(n810) );
  AND2_X1 U913 ( .A1(n810), .A2(n809), .ZN(n811) );
  OR2_X1 U914 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U915 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U916 ( .A1(n816), .A2(n815), .ZN(n831) );
  NOR2_X1 U917 ( .A1(G2090), .A2(G303), .ZN(n817) );
  XOR2_X1 U918 ( .A(KEYINPUT107), .B(n817), .Z(n818) );
  NAND2_X1 U919 ( .A1(n818), .A2(G8), .ZN(n820) );
  NAND2_X1 U920 ( .A1(n820), .A2(n819), .ZN(n822) );
  AND2_X1 U921 ( .A1(n825), .A2(n827), .ZN(n821) );
  AND2_X1 U922 ( .A1(n822), .A2(n821), .ZN(n829) );
  NOR2_X1 U923 ( .A1(G1981), .A2(G305), .ZN(n823) );
  XOR2_X1 U924 ( .A(n823), .B(KEYINPUT24), .Z(n824) );
  NOR2_X1 U925 ( .A1(n825), .A2(n824), .ZN(n826) );
  AND2_X1 U926 ( .A1(n827), .A2(n826), .ZN(n828) );
  NOR2_X1 U927 ( .A1(n829), .A2(n828), .ZN(n830) );
  NAND2_X1 U928 ( .A1(n831), .A2(n830), .ZN(n833) );
  XNOR2_X1 U929 ( .A(G1986), .B(G290), .ZN(n1021) );
  NAND2_X1 U930 ( .A1(n1021), .A2(n845), .ZN(n832) );
  NAND2_X1 U931 ( .A1(n833), .A2(n832), .ZN(n848) );
  NOR2_X1 U932 ( .A1(n907), .A2(G1996), .ZN(n834) );
  XNOR2_X1 U933 ( .A(n834), .B(KEYINPUT108), .ZN(n994) );
  NOR2_X1 U934 ( .A1(G1991), .A2(n911), .ZN(n1003) );
  NOR2_X1 U935 ( .A1(G1986), .A2(G290), .ZN(n835) );
  XOR2_X1 U936 ( .A(n835), .B(KEYINPUT109), .Z(n836) );
  NOR2_X1 U937 ( .A1(n1003), .A2(n836), .ZN(n838) );
  NOR2_X1 U938 ( .A1(n838), .A2(n837), .ZN(n839) );
  NOR2_X1 U939 ( .A1(n994), .A2(n839), .ZN(n840) );
  XNOR2_X1 U940 ( .A(n840), .B(KEYINPUT39), .ZN(n842) );
  NAND2_X1 U941 ( .A1(n842), .A2(n841), .ZN(n844) );
  NAND2_X1 U942 ( .A1(n915), .A2(n843), .ZN(n1000) );
  NAND2_X1 U943 ( .A1(n844), .A2(n1000), .ZN(n846) );
  NAND2_X1 U944 ( .A1(n846), .A2(n845), .ZN(n847) );
  NAND2_X1 U945 ( .A1(n848), .A2(n847), .ZN(n849) );
  XNOR2_X1 U946 ( .A(n850), .B(n849), .ZN(G329) );
  NAND2_X1 U947 ( .A1(G2106), .A2(n851), .ZN(G217) );
  AND2_X1 U948 ( .A1(G15), .A2(G2), .ZN(n852) );
  NAND2_X1 U949 ( .A1(G661), .A2(n852), .ZN(G259) );
  NAND2_X1 U950 ( .A1(G3), .A2(G1), .ZN(n853) );
  NAND2_X1 U951 ( .A1(n854), .A2(n853), .ZN(G188) );
  INV_X1 U953 ( .A(G96), .ZN(G221) );
  NOR2_X1 U954 ( .A1(n856), .A2(n855), .ZN(G325) );
  INV_X1 U955 ( .A(G325), .ZN(G261) );
  XOR2_X1 U956 ( .A(KEYINPUT43), .B(KEYINPUT112), .Z(n858) );
  XNOR2_X1 U957 ( .A(KEYINPUT111), .B(G2678), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U959 ( .A(KEYINPUT42), .B(G2090), .Z(n860) );
  XNOR2_X1 U960 ( .A(G2067), .B(G2072), .ZN(n859) );
  XNOR2_X1 U961 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U962 ( .A(n862), .B(n861), .Z(n864) );
  XNOR2_X1 U963 ( .A(G2100), .B(G2096), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n864), .B(n863), .ZN(n866) );
  XOR2_X1 U965 ( .A(G2078), .B(G2084), .Z(n865) );
  XNOR2_X1 U966 ( .A(n866), .B(n865), .ZN(G227) );
  XOR2_X1 U967 ( .A(G1971), .B(G1956), .Z(n868) );
  XNOR2_X1 U968 ( .A(G1991), .B(G1961), .ZN(n867) );
  XNOR2_X1 U969 ( .A(n868), .B(n867), .ZN(n872) );
  XOR2_X1 U970 ( .A(G1976), .B(G1981), .Z(n870) );
  XNOR2_X1 U971 ( .A(G1986), .B(G1966), .ZN(n869) );
  XNOR2_X1 U972 ( .A(n870), .B(n869), .ZN(n871) );
  XOR2_X1 U973 ( .A(n872), .B(n871), .Z(n874) );
  XNOR2_X1 U974 ( .A(KEYINPUT113), .B(KEYINPUT41), .ZN(n873) );
  XNOR2_X1 U975 ( .A(n874), .B(n873), .ZN(n875) );
  XNOR2_X1 U976 ( .A(G2474), .B(n875), .ZN(n876) );
  XOR2_X1 U977 ( .A(n876), .B(G1996), .Z(G229) );
  NAND2_X1 U978 ( .A1(n900), .A2(G124), .ZN(n877) );
  XNOR2_X1 U979 ( .A(n877), .B(KEYINPUT44), .ZN(n879) );
  NAND2_X1 U980 ( .A1(G112), .A2(n901), .ZN(n878) );
  NAND2_X1 U981 ( .A1(n879), .A2(n878), .ZN(n883) );
  NAND2_X1 U982 ( .A1(G136), .A2(n895), .ZN(n881) );
  NAND2_X1 U983 ( .A1(G100), .A2(n896), .ZN(n880) );
  NAND2_X1 U984 ( .A1(n881), .A2(n880), .ZN(n882) );
  NOR2_X1 U985 ( .A1(n883), .A2(n882), .ZN(G162) );
  NAND2_X1 U986 ( .A1(G130), .A2(n900), .ZN(n885) );
  NAND2_X1 U987 ( .A1(G118), .A2(n901), .ZN(n884) );
  NAND2_X1 U988 ( .A1(n885), .A2(n884), .ZN(n890) );
  NAND2_X1 U989 ( .A1(G142), .A2(n895), .ZN(n887) );
  NAND2_X1 U990 ( .A1(G106), .A2(n896), .ZN(n886) );
  NAND2_X1 U991 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U992 ( .A(KEYINPUT45), .B(n888), .Z(n889) );
  NOR2_X1 U993 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U994 ( .A(G160), .B(n891), .ZN(n914) );
  XOR2_X1 U995 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n893) );
  XNOR2_X1 U996 ( .A(n1002), .B(KEYINPUT114), .ZN(n892) );
  XNOR2_X1 U997 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U998 ( .A(G162), .B(n894), .ZN(n909) );
  NAND2_X1 U999 ( .A1(G139), .A2(n895), .ZN(n898) );
  NAND2_X1 U1000 ( .A1(G103), .A2(n896), .ZN(n897) );
  NAND2_X1 U1001 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U1002 ( .A(KEYINPUT115), .B(n899), .Z(n906) );
  NAND2_X1 U1003 ( .A1(G127), .A2(n900), .ZN(n903) );
  NAND2_X1 U1004 ( .A1(G115), .A2(n901), .ZN(n902) );
  NAND2_X1 U1005 ( .A1(n903), .A2(n902), .ZN(n904) );
  XOR2_X1 U1006 ( .A(KEYINPUT47), .B(n904), .Z(n905) );
  NOR2_X1 U1007 ( .A1(n906), .A2(n905), .ZN(n989) );
  XNOR2_X1 U1008 ( .A(n907), .B(n989), .ZN(n908) );
  XNOR2_X1 U1009 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1010 ( .A(n910), .B(G164), .ZN(n912) );
  XNOR2_X1 U1011 ( .A(n912), .B(n911), .ZN(n913) );
  XNOR2_X1 U1012 ( .A(n914), .B(n913), .ZN(n916) );
  XOR2_X1 U1013 ( .A(n916), .B(n915), .Z(n917) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n917), .ZN(G395) );
  XNOR2_X1 U1015 ( .A(G286), .B(n918), .ZN(n921) );
  XNOR2_X1 U1016 ( .A(G171), .B(n919), .ZN(n920) );
  XNOR2_X1 U1017 ( .A(n921), .B(n920), .ZN(n922) );
  XOR2_X1 U1018 ( .A(n1018), .B(n922), .Z(n923) );
  NOR2_X1 U1019 ( .A1(G37), .A2(n923), .ZN(G397) );
  XOR2_X1 U1020 ( .A(G2451), .B(G2430), .Z(n925) );
  XNOR2_X1 U1021 ( .A(G2438), .B(G2443), .ZN(n924) );
  XNOR2_X1 U1022 ( .A(n925), .B(n924), .ZN(n931) );
  XOR2_X1 U1023 ( .A(G2435), .B(G2454), .Z(n927) );
  XNOR2_X1 U1024 ( .A(G1348), .B(G1341), .ZN(n926) );
  XNOR2_X1 U1025 ( .A(n927), .B(n926), .ZN(n929) );
  XOR2_X1 U1026 ( .A(G2446), .B(G2427), .Z(n928) );
  XNOR2_X1 U1027 ( .A(n929), .B(n928), .ZN(n930) );
  XOR2_X1 U1028 ( .A(n931), .B(n930), .Z(n932) );
  NAND2_X1 U1029 ( .A1(G14), .A2(n932), .ZN(n938) );
  NAND2_X1 U1030 ( .A1(G319), .A2(n938), .ZN(n935) );
  NOR2_X1 U1031 ( .A1(G227), .A2(G229), .ZN(n933) );
  XNOR2_X1 U1032 ( .A(KEYINPUT49), .B(n933), .ZN(n934) );
  NOR2_X1 U1033 ( .A1(n935), .A2(n934), .ZN(n937) );
  NOR2_X1 U1034 ( .A1(G395), .A2(G397), .ZN(n936) );
  NAND2_X1 U1035 ( .A1(n937), .A2(n936), .ZN(G225) );
  INV_X1 U1036 ( .A(G225), .ZN(G308) );
  INV_X1 U1037 ( .A(n938), .ZN(G401) );
  XNOR2_X1 U1038 ( .A(G2084), .B(G34), .ZN(n939) );
  XNOR2_X1 U1039 ( .A(n939), .B(KEYINPUT54), .ZN(n956) );
  XNOR2_X1 U1040 ( .A(G2090), .B(G35), .ZN(n953) );
  XOR2_X1 U1041 ( .A(G2072), .B(G33), .Z(n940) );
  NAND2_X1 U1042 ( .A1(n940), .A2(G28), .ZN(n950) );
  XNOR2_X1 U1043 ( .A(n941), .B(G27), .ZN(n943) );
  XOR2_X1 U1044 ( .A(G1996), .B(G32), .Z(n942) );
  NAND2_X1 U1045 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1046 ( .A(KEYINPUT119), .B(n944), .ZN(n948) );
  XNOR2_X1 U1047 ( .A(G2067), .B(G26), .ZN(n946) );
  XNOR2_X1 U1048 ( .A(G1991), .B(G25), .ZN(n945) );
  NOR2_X1 U1049 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1050 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1051 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1052 ( .A(KEYINPUT53), .B(n951), .ZN(n952) );
  NOR2_X1 U1053 ( .A1(n953), .A2(n952), .ZN(n954) );
  XOR2_X1 U1054 ( .A(KEYINPUT120), .B(n954), .Z(n955) );
  NOR2_X1 U1055 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1056 ( .A(KEYINPUT55), .B(n957), .Z(n958) );
  NOR2_X1 U1057 ( .A1(G29), .A2(n958), .ZN(n988) );
  XOR2_X1 U1058 ( .A(G1348), .B(KEYINPUT59), .Z(n959) );
  XNOR2_X1 U1059 ( .A(G4), .B(n959), .ZN(n961) );
  XNOR2_X1 U1060 ( .A(G20), .B(G1956), .ZN(n960) );
  NOR2_X1 U1061 ( .A1(n961), .A2(n960), .ZN(n965) );
  XNOR2_X1 U1062 ( .A(G1341), .B(G19), .ZN(n963) );
  XNOR2_X1 U1063 ( .A(G1981), .B(G6), .ZN(n962) );
  NOR2_X1 U1064 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1065 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1066 ( .A(n966), .B(KEYINPUT60), .ZN(n981) );
  XNOR2_X1 U1067 ( .A(G5), .B(n967), .ZN(n979) );
  XNOR2_X1 U1068 ( .A(G1966), .B(G21), .ZN(n977) );
  XNOR2_X1 U1069 ( .A(G1971), .B(G22), .ZN(n969) );
  XNOR2_X1 U1070 ( .A(G1976), .B(G23), .ZN(n968) );
  NOR2_X1 U1071 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1072 ( .A(KEYINPUT124), .B(n970), .ZN(n973) );
  XNOR2_X1 U1073 ( .A(G1986), .B(KEYINPUT125), .ZN(n971) );
  XNOR2_X1 U1074 ( .A(n971), .B(G24), .ZN(n972) );
  NAND2_X1 U1075 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1076 ( .A(n974), .B(KEYINPUT58), .ZN(n975) );
  XNOR2_X1 U1077 ( .A(KEYINPUT126), .B(n975), .ZN(n976) );
  NOR2_X1 U1078 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1079 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1080 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1081 ( .A(KEYINPUT127), .B(n982), .Z(n983) );
  XNOR2_X1 U1082 ( .A(n983), .B(KEYINPUT61), .ZN(n985) );
  XNOR2_X1 U1083 ( .A(G16), .B(KEYINPUT123), .ZN(n984) );
  NAND2_X1 U1084 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1085 ( .A1(G11), .A2(n986), .ZN(n987) );
  NOR2_X1 U1086 ( .A1(n988), .A2(n987), .ZN(n1017) );
  XOR2_X1 U1087 ( .A(G2072), .B(n989), .Z(n991) );
  XOR2_X1 U1088 ( .A(G164), .B(G2078), .Z(n990) );
  NOR2_X1 U1089 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1090 ( .A(KEYINPUT50), .B(n992), .ZN(n1008) );
  XNOR2_X1 U1091 ( .A(G160), .B(G2084), .ZN(n997) );
  XOR2_X1 U1092 ( .A(G2090), .B(G162), .Z(n993) );
  NOR2_X1 U1093 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1094 ( .A(KEYINPUT51), .B(n995), .Z(n996) );
  NAND2_X1 U1095 ( .A1(n997), .A2(n996), .ZN(n998) );
  NOR2_X1 U1096 ( .A1(n999), .A2(n998), .ZN(n1001) );
  NAND2_X1 U1097 ( .A1(n1001), .A2(n1000), .ZN(n1006) );
  NOR2_X1 U1098 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1099 ( .A(KEYINPUT116), .B(n1004), .Z(n1005) );
  NOR2_X1 U1100 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1101 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1102 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XNOR2_X1 U1103 ( .A(KEYINPUT117), .B(KEYINPUT52), .ZN(n1011) );
  XNOR2_X1 U1104 ( .A(n1012), .B(n1011), .ZN(n1013) );
  NOR2_X1 U1105 ( .A1(KEYINPUT55), .A2(n1013), .ZN(n1014) );
  XOR2_X1 U1106 ( .A(KEYINPUT118), .B(n1014), .Z(n1015) );
  NAND2_X1 U1107 ( .A1(G29), .A2(n1015), .ZN(n1016) );
  NAND2_X1 U1108 ( .A1(n1017), .A2(n1016), .ZN(n1052) );
  XOR2_X1 U1109 ( .A(KEYINPUT56), .B(G16), .Z(n1050) );
  XNOR2_X1 U1110 ( .A(n1018), .B(G1341), .ZN(n1037) );
  NAND2_X1 U1111 ( .A1(G1971), .A2(G303), .ZN(n1022) );
  INV_X1 U1112 ( .A(KEYINPUT122), .ZN(n1019) );
  NOR2_X1 U1113 ( .A1(n1022), .A2(n1019), .ZN(n1020) );
  NOR2_X1 U1114 ( .A1(n1021), .A2(n1020), .ZN(n1029) );
  XNOR2_X1 U1115 ( .A(G171), .B(G1961), .ZN(n1025) );
  NOR2_X1 U1116 ( .A1(n1039), .A2(KEYINPUT122), .ZN(n1023) );
  NAND2_X1 U1117 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1118 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1119 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1120 ( .A1(n1029), .A2(n1028), .ZN(n1035) );
  XOR2_X1 U1121 ( .A(G168), .B(G1966), .Z(n1030) );
  NOR2_X1 U1122 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XOR2_X1 U1123 ( .A(KEYINPUT57), .B(n1032), .Z(n1033) );
  XNOR2_X1 U1124 ( .A(n1033), .B(KEYINPUT121), .ZN(n1034) );
  NOR2_X1 U1125 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NAND2_X1 U1126 ( .A1(n1037), .A2(n1036), .ZN(n1048) );
  XNOR2_X1 U1127 ( .A(n1038), .B(G1956), .ZN(n1041) );
  NAND2_X1 U1128 ( .A1(KEYINPUT122), .A2(n1039), .ZN(n1040) );
  NAND2_X1 U1129 ( .A1(n1041), .A2(n1040), .ZN(n1044) );
  XNOR2_X1 U1130 ( .A(G1348), .B(n1042), .ZN(n1043) );
  NOR2_X1 U1131 ( .A1(n1044), .A2(n1043), .ZN(n1046) );
  NAND2_X1 U1132 ( .A1(n1046), .A2(n1045), .ZN(n1047) );
  NOR2_X1 U1133 ( .A1(n1048), .A2(n1047), .ZN(n1049) );
  NOR2_X1 U1134 ( .A1(n1050), .A2(n1049), .ZN(n1051) );
  NOR2_X1 U1135 ( .A1(n1052), .A2(n1051), .ZN(n1053) );
  XNOR2_X1 U1136 ( .A(n1053), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1137 ( .A(G311), .ZN(G150) );
endmodule

