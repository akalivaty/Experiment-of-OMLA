

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755;

  OR2_X1 U372 ( .A1(n647), .A2(G902), .ZN(n393) );
  XNOR2_X1 U373 ( .A(n378), .B(n448), .ZN(n722) );
  XNOR2_X1 U374 ( .A(n506), .B(KEYINPUT4), .ZN(n421) );
  XNOR2_X2 U375 ( .A(n471), .B(KEYINPUT76), .ZN(n514) );
  AND2_X2 U376 ( .A1(n376), .A2(n375), .ZN(n374) );
  OR2_X2 U377 ( .A1(n551), .A2(KEYINPUT44), .ZN(n355) );
  NOR2_X1 U378 ( .A1(n677), .A2(n517), .ZN(n482) );
  XNOR2_X1 U379 ( .A(n385), .B(KEYINPUT33), .ZN(n677) );
  XNOR2_X1 U380 ( .A(n608), .B(KEYINPUT85), .ZN(n616) );
  INV_X2 U381 ( .A(G953), .ZN(n749) );
  XNOR2_X2 U382 ( .A(n377), .B(G143), .ZN(n506) );
  XNOR2_X2 U383 ( .A(n426), .B(n425), .ZN(n553) );
  XNOR2_X2 U384 ( .A(n421), .B(n440), .ZN(n743) );
  NOR2_X1 U385 ( .A1(n754), .A2(n631), .ZN(n544) );
  INV_X1 U386 ( .A(n572), .ZN(n690) );
  NAND2_X1 U387 ( .A1(n379), .A2(n607), .ZN(n608) );
  XNOR2_X1 U388 ( .A(n544), .B(KEYINPUT90), .ZN(n403) );
  NOR2_X1 U389 ( .A1(n595), .A2(n753), .ZN(n596) );
  XNOR2_X1 U390 ( .A(n367), .B(n579), .ZN(n629) );
  XNOR2_X1 U391 ( .A(n404), .B(KEYINPUT0), .ZN(n522) );
  NAND2_X1 U392 ( .A1(n582), .A2(n437), .ZN(n404) );
  NAND2_X1 U393 ( .A1(n669), .A2(n666), .ZN(n700) );
  NAND2_X1 U394 ( .A1(n390), .A2(n387), .ZN(n582) );
  AND2_X1 U395 ( .A1(n392), .A2(n391), .ZN(n390) );
  XNOR2_X1 U396 ( .A(n572), .B(KEYINPUT6), .ZN(n597) );
  XNOR2_X1 U397 ( .A(n366), .B(n414), .ZN(n416) );
  XNOR2_X1 U398 ( .A(KEYINPUT91), .B(KEYINPUT18), .ZN(n417) );
  XOR2_X1 U399 ( .A(G122), .B(G107), .Z(n501) );
  XNOR2_X1 U400 ( .A(n365), .B(KEYINPUT45), .ZN(n350) );
  INV_X1 U401 ( .A(n537), .ZN(n351) );
  XNOR2_X1 U402 ( .A(n365), .B(KEYINPUT45), .ZN(n730) );
  XNOR2_X1 U403 ( .A(n528), .B(KEYINPUT22), .ZN(n540) );
  XOR2_X1 U404 ( .A(KEYINPUT62), .B(n647), .Z(n648) );
  AND2_X2 U405 ( .A1(n543), .A2(n542), .ZN(n631) );
  NAND2_X1 U406 ( .A1(n382), .A2(n381), .ZN(n380) );
  AND2_X1 U407 ( .A1(n602), .A2(n601), .ZN(n382) );
  XNOR2_X1 U408 ( .A(n581), .B(n360), .ZN(n381) );
  NAND2_X2 U409 ( .A1(n374), .A2(n370), .ZN(n362) );
  NAND2_X1 U410 ( .A1(n373), .A2(n372), .ZN(n371) );
  NOR2_X1 U411 ( .A1(n688), .A2(n409), .ZN(n683) );
  NAND2_X1 U412 ( .A1(n749), .A2(G224), .ZN(n366) );
  XNOR2_X1 U413 ( .A(G125), .B(G146), .ZN(n451) );
  NOR2_X1 U414 ( .A1(n605), .A2(n571), .ZN(n398) );
  INV_X1 U415 ( .A(KEYINPUT79), .ZN(n429) );
  XNOR2_X1 U416 ( .A(n362), .B(n449), .ZN(n529) );
  XNOR2_X1 U417 ( .A(n405), .B(n412), .ZN(n478) );
  XNOR2_X1 U418 ( .A(n411), .B(n410), .ZN(n405) );
  INV_X1 U419 ( .A(G116), .ZN(n410) );
  XOR2_X1 U420 ( .A(G113), .B(G104), .Z(n488) );
  XNOR2_X1 U421 ( .A(G128), .B(G119), .ZN(n454) );
  XNOR2_X1 U422 ( .A(n380), .B(n359), .ZN(n379) );
  XNOR2_X1 U423 ( .A(n494), .B(n493), .ZN(n633) );
  XNOR2_X1 U424 ( .A(n492), .B(n491), .ZN(n493) );
  NAND2_X1 U425 ( .A1(n592), .A2(n703), .ZN(n384) );
  INV_X1 U426 ( .A(KEYINPUT36), .ZN(n399) );
  XNOR2_X1 U427 ( .A(n467), .B(n466), .ZN(n688) );
  BUF_X1 U428 ( .A(n529), .Z(n682) );
  AND2_X1 U429 ( .A1(n626), .A2(G953), .ZN(n727) );
  AND2_X1 U430 ( .A1(n717), .A2(n678), .ZN(n402) );
  INV_X1 U431 ( .A(G469), .ZN(n373) );
  NAND2_X1 U432 ( .A1(G902), .A2(G469), .ZN(n375) );
  XNOR2_X1 U433 ( .A(G101), .B(KEYINPUT70), .ZN(n411) );
  OR2_X1 U434 ( .A1(n545), .A2(KEYINPUT44), .ZN(n546) );
  AND2_X1 U435 ( .A1(n550), .A2(n534), .ZN(n368) );
  XNOR2_X1 U436 ( .A(G143), .B(G122), .ZN(n484) );
  XOR2_X1 U437 ( .A(KEYINPUT11), .B(KEYINPUT104), .Z(n485) );
  XNOR2_X1 U438 ( .A(G137), .B(G134), .ZN(n439) );
  XNOR2_X1 U439 ( .A(G131), .B(KEYINPUT69), .ZN(n438) );
  INV_X1 U440 ( .A(KEYINPUT17), .ZN(n414) );
  NOR2_X1 U441 ( .A1(n514), .A2(n386), .ZN(n385) );
  INV_X1 U442 ( .A(n597), .ZN(n386) );
  NAND2_X1 U443 ( .A1(G237), .A2(G234), .ZN(n431) );
  OR2_X1 U444 ( .A1(G902), .A2(G237), .ZN(n427) );
  XNOR2_X1 U445 ( .A(G113), .B(KEYINPUT102), .ZN(n472) );
  INV_X1 U446 ( .A(KEYINPUT7), .ZN(n502) );
  AND2_X1 U447 ( .A1(n616), .A2(n352), .ZN(n364) );
  XNOR2_X1 U448 ( .A(KEYINPUT71), .B(G110), .ZN(n442) );
  XNOR2_X1 U449 ( .A(G140), .B(G107), .ZN(n444) );
  XNOR2_X1 U450 ( .A(G104), .B(G101), .ZN(n445) );
  XNOR2_X1 U451 ( .A(n516), .B(KEYINPUT31), .ZN(n665) );
  NOR2_X1 U452 ( .A1(n681), .A2(n517), .ZN(n516) );
  BUF_X1 U453 ( .A(n553), .Z(n605) );
  AND2_X1 U454 ( .A1(n574), .A2(n575), .ZN(n592) );
  NAND2_X1 U455 ( .A1(n389), .A2(n388), .ZN(n387) );
  NOR2_X1 U456 ( .A1(n571), .A2(n354), .ZN(n388) );
  XNOR2_X1 U457 ( .A(n497), .B(n496), .ZN(n524) );
  XNOR2_X1 U458 ( .A(n495), .B(G475), .ZN(n496) );
  XNOR2_X1 U459 ( .A(n406), .B(n478), .ZN(n737) );
  XNOR2_X1 U460 ( .A(n413), .B(n407), .ZN(n406) );
  INV_X1 U461 ( .A(n488), .ZN(n407) );
  XNOR2_X1 U462 ( .A(n461), .B(n460), .ZN(n623) );
  NAND2_X1 U463 ( .A1(n578), .A2(n577), .ZN(n367) );
  NAND2_X1 U464 ( .A1(n395), .A2(n394), .ZN(n671) );
  NAND2_X1 U465 ( .A1(n682), .A2(n356), .ZN(n396) );
  XNOR2_X1 U466 ( .A(n539), .B(n538), .ZN(n754) );
  XNOR2_X1 U467 ( .A(KEYINPUT65), .B(KEYINPUT32), .ZN(n538) );
  XNOR2_X1 U468 ( .A(n724), .B(n723), .ZN(n369) );
  XNOR2_X1 U469 ( .A(n401), .B(n400), .ZN(G75) );
  XNOR2_X1 U470 ( .A(n718), .B(KEYINPUT53), .ZN(n400) );
  NAND2_X1 U471 ( .A1(n679), .A2(n402), .ZN(n401) );
  INV_X1 U472 ( .A(n628), .ZN(n609) );
  XNOR2_X1 U473 ( .A(n384), .B(n358), .ZN(n578) );
  AND2_X1 U474 ( .A1(n609), .A2(KEYINPUT82), .ZN(n352) );
  AND2_X1 U475 ( .A1(n621), .A2(G478), .ZN(n353) );
  XOR2_X1 U476 ( .A(n430), .B(n429), .Z(n354) );
  OR2_X1 U477 ( .A1(n398), .A2(n399), .ZN(n356) );
  AND2_X1 U478 ( .A1(n398), .A2(n399), .ZN(n357) );
  XOR2_X1 U479 ( .A(n576), .B(KEYINPUT39), .Z(n358) );
  INV_X1 U480 ( .A(G902), .ZN(n372) );
  XOR2_X1 U481 ( .A(KEYINPUT86), .B(KEYINPUT48), .Z(n359) );
  XOR2_X1 U482 ( .A(n580), .B(KEYINPUT46), .Z(n360) );
  AND2_X1 U483 ( .A1(n621), .A2(G475), .ZN(n361) );
  NAND2_X1 U484 ( .A1(n362), .A2(n683), .ZN(n570) );
  AND2_X1 U485 ( .A1(n564), .A2(n362), .ZN(n583) );
  NAND2_X1 U486 ( .A1(n363), .A2(n610), .ZN(n619) );
  NAND2_X1 U487 ( .A1(n730), .A2(n364), .ZN(n363) );
  NAND2_X1 U488 ( .A1(n552), .A2(n355), .ZN(n365) );
  NAND2_X1 U489 ( .A1(n533), .A2(n532), .ZN(n545) );
  NAND2_X1 U490 ( .A1(n368), .A2(n403), .ZN(n547) );
  NOR2_X1 U491 ( .A1(n369), .A2(n727), .ZN(G54) );
  INV_X1 U492 ( .A(n622), .ZN(n676) );
  AND2_X2 U493 ( .A1(n622), .A2(n621), .ZN(n646) );
  AND2_X2 U494 ( .A1(n619), .A2(n618), .ZN(n622) );
  OR2_X1 U495 ( .A1(n722), .A2(n371), .ZN(n370) );
  NAND2_X1 U496 ( .A1(n722), .A2(G469), .ZN(n376) );
  NAND2_X1 U497 ( .A1(n529), .A2(n683), .ZN(n471) );
  XNOR2_X2 U498 ( .A(G128), .B(KEYINPUT64), .ZN(n377) );
  XNOR2_X1 U499 ( .A(n378), .B(n480), .ZN(n647) );
  XNOR2_X2 U500 ( .A(n743), .B(G146), .ZN(n378) );
  NAND2_X1 U501 ( .A1(n616), .A2(n609), .ZN(n383) );
  XNOR2_X1 U502 ( .A(n383), .B(n748), .ZN(n750) );
  NAND2_X1 U503 ( .A1(n553), .A2(n354), .ZN(n392) );
  INV_X1 U504 ( .A(n553), .ZN(n389) );
  NAND2_X1 U505 ( .A1(n571), .A2(n354), .ZN(n391) );
  NAND2_X1 U506 ( .A1(n577), .A2(n597), .ZN(n598) );
  XNOR2_X2 U507 ( .A(n393), .B(n481), .ZN(n572) );
  OR2_X1 U508 ( .A1(n600), .A2(n399), .ZN(n394) );
  NOR2_X1 U509 ( .A1(n397), .A2(n396), .ZN(n395) );
  AND2_X1 U510 ( .A1(n600), .A2(n357), .ZN(n397) );
  NAND2_X1 U511 ( .A1(n600), .A2(n699), .ZN(n603) );
  NAND2_X1 U512 ( .A1(n403), .A2(n630), .ZN(n551) );
  AND2_X1 U513 ( .A1(n622), .A2(n361), .ZN(n635) );
  AND2_X1 U514 ( .A1(n622), .A2(n353), .ZN(n726) );
  NOR2_X1 U515 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U516 ( .A(n464), .B(n463), .Z(n408) );
  XOR2_X1 U517 ( .A(n687), .B(n470), .Z(n409) );
  XNOR2_X1 U518 ( .A(n416), .B(n415), .ZN(n420) );
  XNOR2_X1 U519 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U520 ( .A(n453), .B(n483), .ZN(n461) );
  XNOR2_X1 U521 ( .A(n465), .B(n408), .ZN(n466) );
  BUF_X1 U522 ( .A(n665), .Z(n668) );
  XNOR2_X1 U523 ( .A(n625), .B(n624), .ZN(n627) );
  BUF_X1 U524 ( .A(n550), .Z(n630) );
  XOR2_X1 U525 ( .A(KEYINPUT3), .B(G119), .Z(n412) );
  XNOR2_X1 U526 ( .A(n501), .B(KEYINPUT16), .ZN(n413) );
  INV_X1 U527 ( .A(n451), .ZN(n415) );
  XNOR2_X1 U528 ( .A(n417), .B(KEYINPUT81), .ZN(n418) );
  XNOR2_X1 U529 ( .A(n418), .B(n442), .ZN(n419) );
  XNOR2_X1 U530 ( .A(n420), .B(n419), .ZN(n423) );
  INV_X1 U531 ( .A(n421), .ZN(n422) );
  XNOR2_X1 U532 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U533 ( .A(n424), .B(n737), .ZN(n640) );
  XNOR2_X1 U534 ( .A(KEYINPUT15), .B(G902), .ZN(n620) );
  NAND2_X1 U535 ( .A1(n640), .A2(n620), .ZN(n426) );
  NAND2_X1 U536 ( .A1(G210), .A2(n427), .ZN(n425) );
  NAND2_X1 U537 ( .A1(n427), .A2(G214), .ZN(n428) );
  XNOR2_X1 U538 ( .A(n428), .B(KEYINPUT92), .ZN(n699) );
  INV_X1 U539 ( .A(n699), .ZN(n571) );
  XNOR2_X1 U540 ( .A(KEYINPUT19), .B(KEYINPUT67), .ZN(n430) );
  XNOR2_X1 U541 ( .A(n431), .B(KEYINPUT14), .ZN(n433) );
  NAND2_X1 U542 ( .A1(G952), .A2(n433), .ZN(n715) );
  NOR2_X1 U543 ( .A1(n715), .A2(G953), .ZN(n432) );
  XNOR2_X1 U544 ( .A(n432), .B(KEYINPUT93), .ZN(n558) );
  NAND2_X1 U545 ( .A1(G902), .A2(n433), .ZN(n555) );
  INV_X1 U546 ( .A(n555), .ZN(n434) );
  NOR2_X1 U547 ( .A1(G898), .A2(n749), .ZN(n739) );
  NAND2_X1 U548 ( .A1(n434), .A2(n739), .ZN(n435) );
  XNOR2_X1 U549 ( .A(n435), .B(KEYINPUT94), .ZN(n436) );
  NAND2_X1 U550 ( .A1(n558), .A2(n436), .ZN(n437) );
  BUF_X1 U551 ( .A(n522), .Z(n517) );
  XNOR2_X1 U552 ( .A(n439), .B(n438), .ZN(n440) );
  NAND2_X1 U553 ( .A1(n749), .A2(G227), .ZN(n441) );
  XNOR2_X1 U554 ( .A(n441), .B(KEYINPUT95), .ZN(n443) );
  XNOR2_X1 U555 ( .A(n443), .B(n442), .ZN(n447) );
  XNOR2_X1 U556 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U557 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U558 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n449) );
  NAND2_X1 U559 ( .A1(G234), .A2(n749), .ZN(n450) );
  XOR2_X1 U560 ( .A(KEYINPUT8), .B(n450), .Z(n498) );
  NAND2_X1 U561 ( .A1(G221), .A2(n498), .ZN(n453) );
  XNOR2_X1 U562 ( .A(G140), .B(KEYINPUT10), .ZN(n452) );
  XNOR2_X1 U563 ( .A(n452), .B(n451), .ZN(n483) );
  XOR2_X1 U564 ( .A(G137), .B(G110), .Z(n455) );
  XNOR2_X1 U565 ( .A(n455), .B(n454), .ZN(n459) );
  XOR2_X1 U566 ( .A(KEYINPUT24), .B(KEYINPUT96), .Z(n457) );
  XNOR2_X1 U567 ( .A(KEYINPUT97), .B(KEYINPUT23), .ZN(n456) );
  XNOR2_X1 U568 ( .A(n457), .B(n456), .ZN(n458) );
  XOR2_X1 U569 ( .A(n459), .B(n458), .Z(n460) );
  NOR2_X1 U570 ( .A1(G902), .A2(n623), .ZN(n467) );
  NAND2_X1 U571 ( .A1(G234), .A2(n620), .ZN(n462) );
  XNOR2_X1 U572 ( .A(KEYINPUT20), .B(n462), .ZN(n468) );
  NAND2_X1 U573 ( .A1(G217), .A2(n468), .ZN(n465) );
  XOR2_X1 U574 ( .A(KEYINPUT98), .B(KEYINPUT25), .Z(n464) );
  XNOR2_X1 U575 ( .A(KEYINPUT80), .B(KEYINPUT99), .ZN(n463) );
  NAND2_X1 U576 ( .A1(n468), .A2(G221), .ZN(n469) );
  XNOR2_X1 U577 ( .A(n469), .B(KEYINPUT21), .ZN(n687) );
  INV_X1 U578 ( .A(KEYINPUT100), .ZN(n470) );
  XNOR2_X1 U579 ( .A(n472), .B(KEYINPUT5), .ZN(n474) );
  XOR2_X1 U580 ( .A(KEYINPUT101), .B(KEYINPUT77), .Z(n473) );
  XNOR2_X1 U581 ( .A(n474), .B(n473), .ZN(n477) );
  NOR2_X1 U582 ( .A1(G237), .A2(G953), .ZN(n475) );
  XNOR2_X1 U583 ( .A(n475), .B(KEYINPUT78), .ZN(n487) );
  NAND2_X1 U584 ( .A1(n487), .A2(G210), .ZN(n476) );
  XNOR2_X1 U585 ( .A(n477), .B(n476), .ZN(n479) );
  XNOR2_X1 U586 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U587 ( .A(G472), .B(KEYINPUT73), .ZN(n481) );
  XNOR2_X1 U588 ( .A(n482), .B(KEYINPUT34), .ZN(n510) );
  INV_X1 U589 ( .A(n483), .ZN(n742) );
  XNOR2_X1 U590 ( .A(G131), .B(n742), .ZN(n494) );
  XNOR2_X1 U591 ( .A(n485), .B(n484), .ZN(n486) );
  XOR2_X1 U592 ( .A(KEYINPUT12), .B(n486), .Z(n492) );
  NAND2_X1 U593 ( .A1(n487), .A2(G214), .ZN(n490) );
  XNOR2_X1 U594 ( .A(n488), .B(KEYINPUT105), .ZN(n489) );
  XNOR2_X1 U595 ( .A(n490), .B(n489), .ZN(n491) );
  NOR2_X1 U596 ( .A1(G902), .A2(n633), .ZN(n497) );
  XNOR2_X1 U597 ( .A(KEYINPUT13), .B(KEYINPUT106), .ZN(n495) );
  XOR2_X1 U598 ( .A(KEYINPUT9), .B(G134), .Z(n500) );
  NAND2_X1 U599 ( .A1(G217), .A2(n498), .ZN(n499) );
  XNOR2_X1 U600 ( .A(n500), .B(n499), .ZN(n505) );
  XNOR2_X1 U601 ( .A(n501), .B(G116), .ZN(n503) );
  XNOR2_X1 U602 ( .A(n505), .B(n504), .ZN(n507) );
  XNOR2_X1 U603 ( .A(n506), .B(n507), .ZN(n725) );
  NAND2_X1 U604 ( .A1(n725), .A2(n372), .ZN(n508) );
  XNOR2_X1 U605 ( .A(n508), .B(G478), .ZN(n523) );
  NAND2_X1 U606 ( .A1(n524), .A2(n523), .ZN(n591) );
  INV_X1 U607 ( .A(n591), .ZN(n509) );
  NAND2_X1 U608 ( .A1(n510), .A2(n509), .ZN(n513) );
  INV_X1 U609 ( .A(KEYINPUT84), .ZN(n511) );
  XNOR2_X1 U610 ( .A(n511), .B(KEYINPUT35), .ZN(n512) );
  XNOR2_X1 U611 ( .A(n513), .B(n512), .ZN(n550) );
  NOR2_X1 U612 ( .A1(n514), .A2(n572), .ZN(n515) );
  XNOR2_X1 U613 ( .A(n515), .B(KEYINPUT103), .ZN(n681) );
  INV_X1 U614 ( .A(n517), .ZN(n519) );
  NOR2_X1 U615 ( .A1(n570), .A2(n690), .ZN(n518) );
  NAND2_X1 U616 ( .A1(n519), .A2(n518), .ZN(n655) );
  NAND2_X1 U617 ( .A1(n665), .A2(n655), .ZN(n521) );
  INV_X1 U618 ( .A(n523), .ZN(n520) );
  OR2_X1 U619 ( .A1(n524), .A2(n520), .ZN(n669) );
  NAND2_X1 U620 ( .A1(n524), .A2(n520), .ZN(n666) );
  NAND2_X1 U621 ( .A1(n521), .A2(n700), .ZN(n533) );
  INV_X1 U622 ( .A(n522), .ZN(n527) );
  NOR2_X1 U623 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U624 ( .A(n525), .B(KEYINPUT107), .ZN(n701) );
  NOR2_X1 U625 ( .A1(n701), .A2(n409), .ZN(n526) );
  NAND2_X1 U626 ( .A1(n527), .A2(n526), .ZN(n528) );
  OR2_X1 U627 ( .A1(n682), .A2(n688), .ZN(n530) );
  OR2_X1 U628 ( .A1(n530), .A2(n597), .ZN(n531) );
  NOR2_X1 U629 ( .A1(n351), .A2(n531), .ZN(n653) );
  INV_X1 U630 ( .A(n653), .ZN(n532) );
  INV_X1 U631 ( .A(n545), .ZN(n534) );
  INV_X1 U632 ( .A(n540), .ZN(n537) );
  NAND2_X1 U633 ( .A1(n682), .A2(n688), .ZN(n535) );
  NOR2_X1 U634 ( .A1(n535), .A2(n597), .ZN(n536) );
  NAND2_X1 U635 ( .A1(n537), .A2(n536), .ZN(n539) );
  NOR2_X1 U636 ( .A1(n540), .A2(n682), .ZN(n541) );
  XNOR2_X1 U637 ( .A(n541), .B(KEYINPUT108), .ZN(n543) );
  AND2_X1 U638 ( .A1(n572), .A2(n688), .ZN(n542) );
  NAND2_X1 U639 ( .A1(n547), .A2(n546), .ZN(n549) );
  INV_X1 U640 ( .A(KEYINPUT89), .ZN(n548) );
  XNOR2_X1 U641 ( .A(n549), .B(n548), .ZN(n552) );
  NOR2_X1 U642 ( .A1(n571), .A2(n701), .ZN(n705) );
  XNOR2_X1 U643 ( .A(n605), .B(KEYINPUT38), .ZN(n703) );
  NAND2_X1 U644 ( .A1(n705), .A2(n703), .ZN(n554) );
  XNOR2_X1 U645 ( .A(n554), .B(KEYINPUT41), .ZN(n698) );
  NOR2_X1 U646 ( .A1(G900), .A2(n555), .ZN(n556) );
  NAND2_X1 U647 ( .A1(n556), .A2(G953), .ZN(n557) );
  NAND2_X1 U648 ( .A1(n558), .A2(n557), .ZN(n568) );
  INV_X1 U649 ( .A(n687), .ZN(n559) );
  AND2_X1 U650 ( .A1(n559), .A2(n688), .ZN(n560) );
  NAND2_X1 U651 ( .A1(n568), .A2(n560), .ZN(n599) );
  INV_X1 U652 ( .A(n599), .ZN(n561) );
  NAND2_X1 U653 ( .A1(n690), .A2(n561), .ZN(n563) );
  INV_X1 U654 ( .A(KEYINPUT28), .ZN(n562) );
  XNOR2_X1 U655 ( .A(n563), .B(n562), .ZN(n564) );
  NAND2_X1 U656 ( .A1(n698), .A2(n583), .ZN(n567) );
  INV_X1 U657 ( .A(KEYINPUT111), .ZN(n565) );
  XNOR2_X1 U658 ( .A(n565), .B(KEYINPUT42), .ZN(n566) );
  XNOR2_X1 U659 ( .A(n567), .B(n566), .ZN(n755) );
  INV_X1 U660 ( .A(n568), .ZN(n569) );
  NOR2_X1 U661 ( .A1(n570), .A2(n569), .ZN(n575) );
  XNOR2_X1 U662 ( .A(n573), .B(KEYINPUT30), .ZN(n574) );
  INV_X1 U663 ( .A(KEYINPUT72), .ZN(n576) );
  INV_X1 U664 ( .A(n666), .ZN(n577) );
  XNOR2_X1 U665 ( .A(KEYINPUT110), .B(KEYINPUT40), .ZN(n579) );
  NAND2_X1 U666 ( .A1(n755), .A2(n629), .ZN(n581) );
  INV_X1 U667 ( .A(KEYINPUT87), .ZN(n580) );
  AND2_X2 U668 ( .A1(n583), .A2(n582), .ZN(n663) );
  NAND2_X1 U669 ( .A1(n663), .A2(n700), .ZN(n584) );
  NAND2_X1 U670 ( .A1(n584), .A2(KEYINPUT47), .ZN(n590) );
  INV_X1 U671 ( .A(n700), .ZN(n586) );
  XNOR2_X1 U672 ( .A(KEYINPUT68), .B(KEYINPUT47), .ZN(n585) );
  NOR2_X1 U673 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U674 ( .A(KEYINPUT75), .B(n587), .Z(n588) );
  NAND2_X1 U675 ( .A1(n588), .A2(n663), .ZN(n589) );
  NAND2_X1 U676 ( .A1(n590), .A2(n589), .ZN(n595) );
  NOR2_X1 U677 ( .A1(n591), .A2(n605), .ZN(n593) );
  NAND2_X1 U678 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U679 ( .A(n594), .B(KEYINPUT109), .ZN(n753) );
  XNOR2_X1 U680 ( .A(n596), .B(KEYINPUT74), .ZN(n602) );
  NOR2_X1 U681 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U682 ( .A(n671), .B(KEYINPUT88), .ZN(n601) );
  OR2_X1 U683 ( .A1(n682), .A2(n603), .ZN(n604) );
  XNOR2_X1 U684 ( .A(n604), .B(KEYINPUT43), .ZN(n606) );
  AND2_X1 U685 ( .A1(n606), .A2(n605), .ZN(n673) );
  INV_X1 U686 ( .A(n673), .ZN(n607) );
  INV_X1 U687 ( .A(n669), .ZN(n659) );
  AND2_X1 U688 ( .A1(n578), .A2(n659), .ZN(n628) );
  INV_X1 U689 ( .A(KEYINPUT82), .ZN(n611) );
  INV_X1 U690 ( .A(KEYINPUT2), .ZN(n610) );
  NAND2_X1 U691 ( .A1(n628), .A2(n611), .ZN(n614) );
  AND2_X1 U692 ( .A1(KEYINPUT82), .A2(KEYINPUT2), .ZN(n612) );
  NAND2_X1 U693 ( .A1(n609), .A2(n612), .ZN(n613) );
  NAND2_X1 U694 ( .A1(n614), .A2(n613), .ZN(n615) );
  AND2_X1 U695 ( .A1(n616), .A2(n615), .ZN(n617) );
  NAND2_X1 U696 ( .A1(n350), .A2(n617), .ZN(n618) );
  INV_X1 U697 ( .A(n620), .ZN(n621) );
  BUF_X1 U698 ( .A(n646), .Z(n719) );
  NAND2_X1 U699 ( .A1(n719), .A2(G217), .ZN(n625) );
  XOR2_X1 U700 ( .A(n623), .B(KEYINPUT123), .Z(n624) );
  INV_X1 U701 ( .A(G952), .ZN(n626) );
  NOR2_X1 U702 ( .A1(n627), .A2(n727), .ZN(G66) );
  XOR2_X1 U703 ( .A(G134), .B(n628), .Z(G36) );
  XNOR2_X1 U704 ( .A(n629), .B(G131), .ZN(G33) );
  XNOR2_X1 U705 ( .A(n630), .B(G122), .ZN(G24) );
  XOR2_X1 U706 ( .A(n631), .B(G110), .Z(G12) );
  XOR2_X1 U707 ( .A(KEYINPUT120), .B(KEYINPUT59), .Z(n632) );
  XNOR2_X1 U708 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U709 ( .A(n635), .B(n634), .ZN(n636) );
  INV_X1 U710 ( .A(n727), .ZN(n650) );
  NAND2_X1 U711 ( .A1(n636), .A2(n650), .ZN(n638) );
  XNOR2_X1 U712 ( .A(KEYINPUT121), .B(KEYINPUT60), .ZN(n637) );
  XNOR2_X1 U713 ( .A(n638), .B(n637), .ZN(G60) );
  NAND2_X1 U714 ( .A1(n646), .A2(G210), .ZN(n642) );
  XOR2_X1 U715 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n639) );
  XNOR2_X1 U716 ( .A(n640), .B(n639), .ZN(n641) );
  XNOR2_X1 U717 ( .A(n642), .B(n641), .ZN(n643) );
  NAND2_X1 U718 ( .A1(n643), .A2(n650), .ZN(n645) );
  INV_X1 U719 ( .A(KEYINPUT56), .ZN(n644) );
  XNOR2_X1 U720 ( .A(n645), .B(n644), .ZN(G51) );
  NAND2_X1 U721 ( .A1(n646), .A2(G472), .ZN(n649) );
  XNOR2_X1 U722 ( .A(n649), .B(n648), .ZN(n651) );
  NAND2_X1 U723 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U724 ( .A(n652), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U725 ( .A(G101), .B(n653), .Z(G3) );
  NOR2_X1 U726 ( .A1(n666), .A2(n655), .ZN(n654) );
  XOR2_X1 U727 ( .A(G104), .B(n654), .Z(G6) );
  NOR2_X1 U728 ( .A1(n669), .A2(n655), .ZN(n657) );
  XNOR2_X1 U729 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n656) );
  XNOR2_X1 U730 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U731 ( .A(G107), .B(n658), .ZN(G9) );
  XOR2_X1 U732 ( .A(KEYINPUT112), .B(KEYINPUT29), .Z(n661) );
  NAND2_X1 U733 ( .A1(n663), .A2(n659), .ZN(n660) );
  XNOR2_X1 U734 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U735 ( .A(G128), .B(n662), .ZN(G30) );
  NAND2_X1 U736 ( .A1(n663), .A2(n577), .ZN(n664) );
  XNOR2_X1 U737 ( .A(n664), .B(G146), .ZN(G48) );
  NOR2_X1 U738 ( .A1(n666), .A2(n668), .ZN(n667) );
  XOR2_X1 U739 ( .A(G113), .B(n667), .Z(G15) );
  NOR2_X1 U740 ( .A1(n669), .A2(n668), .ZN(n670) );
  XOR2_X1 U741 ( .A(G116), .B(n670), .Z(G18) );
  XOR2_X1 U742 ( .A(n671), .B(G125), .Z(n672) );
  XNOR2_X1 U743 ( .A(n672), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U744 ( .A(G140), .B(n673), .ZN(n674) );
  XNOR2_X1 U745 ( .A(n674), .B(KEYINPUT113), .ZN(G42) );
  XNOR2_X1 U746 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n718) );
  INV_X1 U747 ( .A(KEYINPUT83), .ZN(n675) );
  XNOR2_X1 U748 ( .A(n676), .B(n675), .ZN(n679) );
  INV_X1 U749 ( .A(n677), .ZN(n709) );
  NAND2_X1 U750 ( .A1(n698), .A2(n709), .ZN(n678) );
  XNOR2_X1 U751 ( .A(KEYINPUT52), .B(KEYINPUT115), .ZN(n680) );
  XNOR2_X1 U752 ( .A(n680), .B(KEYINPUT116), .ZN(n713) );
  INV_X1 U753 ( .A(n682), .ZN(n685) );
  INV_X1 U754 ( .A(n683), .ZN(n684) );
  NAND2_X1 U755 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U756 ( .A(n686), .B(KEYINPUT50), .ZN(n694) );
  NAND2_X1 U757 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U758 ( .A(KEYINPUT49), .B(n689), .ZN(n691) );
  NOR2_X1 U759 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U760 ( .A(n692), .B(KEYINPUT114), .ZN(n693) );
  NAND2_X1 U761 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U762 ( .A1(n681), .A2(n695), .ZN(n696) );
  XOR2_X1 U763 ( .A(KEYINPUT51), .B(n696), .Z(n697) );
  NAND2_X1 U764 ( .A1(n698), .A2(n697), .ZN(n711) );
  NAND2_X1 U765 ( .A1(n700), .A2(n699), .ZN(n702) );
  NAND2_X1 U766 ( .A1(n702), .A2(n701), .ZN(n704) );
  NAND2_X1 U767 ( .A1(n704), .A2(n703), .ZN(n707) );
  INV_X1 U768 ( .A(n705), .ZN(n706) );
  NAND2_X1 U769 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U770 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U771 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U772 ( .A(n713), .B(n712), .ZN(n714) );
  NOR2_X1 U773 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U774 ( .A1(G953), .A2(n716), .ZN(n717) );
  NAND2_X1 U775 ( .A1(n719), .A2(G469), .ZN(n724) );
  XNOR2_X1 U776 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n720) );
  XNOR2_X1 U777 ( .A(n720), .B(KEYINPUT57), .ZN(n721) );
  XNOR2_X1 U778 ( .A(n722), .B(n721), .ZN(n723) );
  XNOR2_X1 U779 ( .A(n726), .B(n725), .ZN(n728) );
  NOR2_X1 U780 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U781 ( .A(KEYINPUT122), .B(n729), .ZN(G63) );
  NAND2_X1 U782 ( .A1(n350), .A2(n749), .ZN(n736) );
  NAND2_X1 U783 ( .A1(G224), .A2(G953), .ZN(n731) );
  XNOR2_X1 U784 ( .A(n731), .B(KEYINPUT124), .ZN(n732) );
  XNOR2_X1 U785 ( .A(KEYINPUT61), .B(n732), .ZN(n733) );
  NAND2_X1 U786 ( .A1(n733), .A2(G898), .ZN(n734) );
  XOR2_X1 U787 ( .A(KEYINPUT125), .B(n734), .Z(n735) );
  NAND2_X1 U788 ( .A1(n736), .A2(n735), .ZN(n741) );
  XOR2_X1 U789 ( .A(G110), .B(n737), .Z(n738) );
  NOR2_X1 U790 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U791 ( .A(n741), .B(n740), .ZN(G69) );
  XOR2_X1 U792 ( .A(n743), .B(n742), .Z(n747) );
  XOR2_X1 U793 ( .A(n747), .B(G227), .Z(n744) );
  XNOR2_X1 U794 ( .A(n744), .B(KEYINPUT127), .ZN(n745) );
  NAND2_X1 U795 ( .A1(G900), .A2(n745), .ZN(n746) );
  NAND2_X1 U796 ( .A1(n746), .A2(G953), .ZN(n752) );
  XNOR2_X1 U797 ( .A(n747), .B(KEYINPUT126), .ZN(n748) );
  NAND2_X1 U798 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U799 ( .A1(n752), .A2(n751), .ZN(G72) );
  XOR2_X1 U800 ( .A(G143), .B(n753), .Z(G45) );
  XOR2_X1 U801 ( .A(n754), .B(G119), .Z(G21) );
  XNOR2_X1 U802 ( .A(G137), .B(n755), .ZN(G39) );
endmodule

