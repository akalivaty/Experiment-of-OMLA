//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 1 0 0 0 0 1 0 0 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0 1 0 0 0 1 1 0 1 0 0 0 0 1 0 1 1 0 0 1 0 0 0 0 0 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n839, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n916, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1015, new_n1016;
  INV_X1    g000(.A(G15gat), .ZN(new_n202));
  INV_X1    g001(.A(G22gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G15gat), .A2(G22gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G1gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT16), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G8gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n204), .A2(new_n207), .A3(new_n205), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT93), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND4_X1  g013(.A1(new_n209), .A2(KEYINPUT93), .A3(new_n210), .A4(new_n211), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n209), .A2(KEYINPUT92), .A3(new_n211), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n217), .B(G8gat), .C1(KEYINPUT92), .C2(new_n209), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(G43gat), .B(G50gat), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G29gat), .ZN(new_n223));
  INV_X1    g022(.A(G36gat), .ZN(new_n224));
  AND3_X1   g023(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT14), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n224), .ZN(new_n226));
  NAND2_X1  g025(.A1(G29gat), .A2(G36gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT14), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n225), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT15), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT15), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n228), .A2(new_n226), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n231), .B1(new_n232), .B2(new_n225), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n222), .B1(new_n230), .B2(new_n233), .ZN(new_n234));
  NOR3_X1   g033(.A1(new_n232), .A2(new_n231), .A3(new_n225), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n235), .A2(new_n221), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT17), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n229), .A2(KEYINPUT15), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n221), .B1(new_n238), .B2(new_n235), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT17), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n230), .A2(new_n222), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n220), .A2(new_n237), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G229gat), .A2(G233gat), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n234), .A2(new_n236), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT94), .ZN(new_n246));
  AND3_X1   g045(.A1(new_n245), .A2(new_n219), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n246), .B1(new_n245), .B2(new_n219), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n243), .B(new_n244), .C1(new_n247), .C2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT95), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(KEYINPUT18), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n245), .A2(new_n219), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT94), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n245), .A2(new_n219), .A3(new_n246), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n257), .A2(new_n244), .A3(new_n251), .A4(new_n243), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n253), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n250), .A2(KEYINPUT18), .ZN(new_n260));
  OAI22_X1  g059(.A1(new_n247), .A2(new_n248), .B1(new_n219), .B2(new_n245), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n244), .B(KEYINPUT13), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n260), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G113gat), .B(G141gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(G197gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(KEYINPUT11), .ZN(new_n267));
  INV_X1    g066(.A(G169gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(KEYINPUT12), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n259), .A2(new_n264), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT96), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT96), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n259), .A2(new_n264), .A3(new_n273), .A4(new_n270), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n260), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n245), .A2(new_n219), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n277), .B1(new_n255), .B2(new_n256), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n276), .B1(new_n278), .B2(new_n262), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n279), .B1(new_n253), .B2(new_n258), .ZN(new_n280));
  OR2_X1    g079(.A1(new_n280), .A2(new_n270), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n284));
  INV_X1    g083(.A(G197gat), .ZN(new_n285));
  INV_X1    g084(.A(G204gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G197gat), .A2(G204gat), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n284), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n289), .A2(KEYINPUT74), .ZN(new_n290));
  OR2_X1    g089(.A1(G211gat), .A2(G218gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(G211gat), .A2(G218gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n290), .B(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT3), .ZN(new_n296));
  NOR2_X1   g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(G155gat), .A2(G162gat), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(G141gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(G148gat), .ZN(new_n301));
  INV_X1    g100(.A(G148gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G141gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT2), .ZN(new_n305));
  AOI211_X1 g104(.A(new_n297), .B(new_n299), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n301), .ZN(new_n308));
  XNOR2_X1  g107(.A(KEYINPUT77), .B(G148gat), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n308), .B1(new_n309), .B2(G141gat), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n299), .B1(new_n305), .B2(new_n297), .ZN(new_n311));
  NOR3_X1   g110(.A1(new_n310), .A2(new_n311), .A3(KEYINPUT78), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT78), .ZN(new_n313));
  AND2_X1   g112(.A1(KEYINPUT77), .A2(G148gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(KEYINPUT77), .A2(G148gat), .ZN(new_n315));
  OAI21_X1  g114(.A(G141gat), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(new_n301), .ZN(new_n317));
  INV_X1    g116(.A(new_n297), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n298), .B1(new_n318), .B2(KEYINPUT2), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n313), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n296), .B(new_n307), .C1(new_n312), .C2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT29), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n295), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n307), .B1(new_n312), .B2(new_n320), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT79), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT78), .B1(new_n310), .B2(new_n311), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n317), .A2(new_n313), .A3(new_n319), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n306), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT79), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n290), .B(new_n293), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n296), .B1(new_n332), .B2(KEYINPUT29), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n323), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G228gat), .A2(G233gat), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT81), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT29), .B1(new_n328), .B2(new_n296), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT80), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n287), .A2(new_n288), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n340), .B(new_n293), .C1(new_n341), .C2(new_n284), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n293), .A2(new_n340), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n291), .A2(KEYINPUT80), .A3(new_n292), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n343), .A2(new_n289), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n342), .A2(new_n345), .A3(new_n322), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n346), .A2(new_n296), .ZN(new_n347));
  OAI22_X1  g146(.A1(new_n339), .A2(new_n295), .B1(new_n328), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n338), .B1(new_n348), .B2(new_n335), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n326), .A2(new_n327), .ZN(new_n350));
  AOI22_X1  g149(.A1(new_n350), .A2(new_n307), .B1(new_n346), .B2(new_n296), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n338), .B(new_n335), .C1(new_n323), .C2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n337), .B1(new_n349), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT82), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT82), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n356), .B(new_n337), .C1(new_n349), .C2(new_n353), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n355), .A2(G22gat), .A3(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT83), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  XOR2_X1   g159(.A(G78gat), .B(G106gat), .Z(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(KEYINPUT31), .ZN(new_n362));
  XOR2_X1   g161(.A(new_n362), .B(G50gat), .Z(new_n363));
  NOR3_X1   g162(.A1(new_n354), .A2(KEYINPUT84), .A3(G22gat), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT84), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n335), .B1(new_n323), .B2(new_n351), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT81), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n367), .A2(new_n352), .B1(new_n336), .B2(new_n334), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n365), .B1(new_n368), .B2(new_n203), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n364), .A2(new_n369), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n355), .A2(KEYINPUT83), .A3(G22gat), .A4(new_n357), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n360), .A2(new_n363), .A3(new_n370), .A4(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n363), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n354), .A2(G22gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n368), .A2(new_n203), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n372), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT85), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT85), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n372), .A2(new_n379), .A3(new_n376), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(G227gat), .A2(G233gat), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(G169gat), .A2(G176gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n384), .B(KEYINPUT23), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G169gat), .A2(G176gat), .ZN(new_n387));
  NAND3_X1  g186(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n388), .B1(G183gat), .B2(G190gat), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT64), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n390), .B(new_n391), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n386), .B(new_n387), .C1(new_n389), .C2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT25), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT25), .B1(new_n389), .B2(new_n390), .ZN(new_n396));
  XOR2_X1   g195(.A(new_n387), .B(KEYINPUT65), .Z(new_n397));
  NOR3_X1   g196(.A1(new_n396), .A2(new_n397), .A3(new_n385), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT68), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT66), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT26), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n384), .A2(new_n405), .ZN(new_n406));
  OAI211_X1 g205(.A(KEYINPUT66), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n404), .A2(new_n387), .A3(new_n406), .A4(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(G183gat), .A2(G190gat), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT67), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n408), .A2(KEYINPUT67), .A3(new_n409), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT28), .ZN(new_n415));
  XNOR2_X1  g214(.A(KEYINPUT27), .B(G183gat), .ZN(new_n416));
  INV_X1    g215(.A(G190gat), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AND2_X1   g217(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n419));
  NOR2_X1   g218(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n415), .B(new_n417), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n401), .B1(new_n414), .B2(new_n423), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n408), .A2(KEYINPUT67), .A3(new_n409), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT67), .B1(new_n408), .B2(new_n409), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n401), .B(new_n423), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n400), .B1(new_n424), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT69), .ZN(new_n430));
  INV_X1    g229(.A(G127gat), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n431), .A2(G134gat), .ZN(new_n432));
  INV_X1    g231(.A(G134gat), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n433), .A2(G127gat), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n430), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(G120gat), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(G113gat), .ZN(new_n437));
  INV_X1    g236(.A(G113gat), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(G120gat), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT1), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n433), .A2(G127gat), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n431), .A2(G134gat), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n441), .A2(new_n442), .A3(KEYINPUT69), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n435), .A2(new_n440), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT70), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n432), .A2(new_n434), .ZN(new_n447));
  OR2_X1    g246(.A1(new_n447), .A2(new_n440), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n435), .A2(KEYINPUT70), .A3(new_n440), .A4(new_n443), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n446), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n429), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n398), .B1(new_n393), .B2(new_n394), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n423), .B1(new_n425), .B2(new_n426), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT68), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n452), .B1(new_n454), .B2(new_n427), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n446), .A2(new_n448), .A3(new_n449), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n383), .B1(new_n451), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT34), .ZN(new_n459));
  OR3_X1    g258(.A1(new_n458), .A2(KEYINPUT72), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n458), .A2(new_n459), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT72), .B1(new_n458), .B2(new_n459), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT32), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n451), .A2(new_n383), .A3(new_n457), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT71), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n451), .A2(new_n457), .A3(KEYINPUT71), .A4(new_n383), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n464), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT33), .B1(new_n467), .B2(new_n468), .ZN(new_n470));
  XNOR2_X1  g269(.A(G15gat), .B(G43gat), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n471), .B(G71gat), .ZN(new_n472));
  INV_X1    g271(.A(G99gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n472), .B(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NOR3_X1   g274(.A1(new_n469), .A2(new_n470), .A3(new_n475), .ZN(new_n476));
  AOI221_X4 g275(.A(new_n464), .B1(KEYINPUT33), .B2(new_n474), .C1(new_n467), .C2(new_n468), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n463), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT73), .ZN(new_n479));
  INV_X1    g278(.A(new_n469), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n467), .A2(new_n468), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT33), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n480), .A2(new_n483), .A3(new_n474), .ZN(new_n484));
  INV_X1    g283(.A(new_n477), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n478), .A2(new_n479), .A3(new_n487), .ZN(new_n488));
  OAI211_X1 g287(.A(KEYINPUT73), .B(new_n463), .C1(new_n476), .C2(new_n477), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT75), .ZN(new_n491));
  INV_X1    g290(.A(G226gat), .ZN(new_n492));
  INV_X1    g291(.A(G233gat), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n400), .A2(new_n453), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(KEYINPUT29), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n455), .A2(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n491), .B1(new_n497), .B2(new_n332), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n400), .B(new_n494), .C1(new_n424), .C2(new_n428), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n495), .A2(new_n496), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n501), .A2(KEYINPUT75), .A3(new_n295), .ZN(new_n502));
  INV_X1    g301(.A(new_n494), .ZN(new_n503));
  INV_X1    g302(.A(new_n496), .ZN(new_n504));
  OAI221_X1 g303(.A(new_n332), .B1(new_n495), .B2(new_n503), .C1(new_n455), .C2(new_n504), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n498), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G8gat), .B(G36gat), .ZN(new_n507));
  INV_X1    g306(.A(G64gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n507), .B(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(G92gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n509), .B(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n506), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n506), .A2(KEYINPUT76), .A3(KEYINPUT30), .A4(new_n512), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT76), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n498), .A2(new_n502), .A3(new_n505), .A4(new_n512), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT30), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n513), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(G1gat), .B(G29gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(KEYINPUT0), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(G57gat), .ZN(new_n522));
  INV_X1    g321(.A(G85gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n522), .B(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT4), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n450), .A2(new_n526), .A3(new_n328), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT4), .B1(new_n324), .B2(new_n456), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(G225gat), .A2(G233gat), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n296), .B1(new_n325), .B2(new_n330), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n321), .A2(new_n456), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n529), .B(new_n530), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT5), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n329), .B1(new_n350), .B2(new_n307), .ZN(new_n536));
  AOI211_X1 g335(.A(KEYINPUT79), .B(new_n306), .C1(new_n326), .C2(new_n327), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n456), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n324), .A2(new_n456), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n530), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(KEYINPUT3), .B1(new_n536), .B2(new_n537), .ZN(new_n542));
  INV_X1    g341(.A(new_n532), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n542), .A2(new_n543), .B1(new_n528), .B2(new_n527), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n541), .B1(new_n544), .B2(new_n530), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n525), .B(new_n535), .C1(new_n545), .C2(new_n534), .ZN(new_n546));
  INV_X1    g345(.A(new_n530), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n450), .B1(new_n325), .B2(new_n330), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n547), .B1(new_n548), .B2(new_n539), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n534), .B1(new_n533), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT5), .B1(new_n544), .B2(new_n530), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n524), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT6), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n546), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n550), .A2(new_n551), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n555), .A2(KEYINPUT6), .A3(new_n525), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n516), .A2(new_n517), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n519), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n381), .A2(new_n490), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT35), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n478), .A2(new_n487), .ZN(new_n563));
  OR2_X1    g362(.A1(KEYINPUT91), .A2(KEYINPUT35), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT35), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n519), .A2(new_n565), .A3(new_n557), .A4(new_n558), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT91), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n381), .A2(new_n563), .A3(new_n564), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n562), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n519), .A2(new_n558), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT86), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n571), .B1(new_n544), .B2(new_n530), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n529), .B1(new_n531), .B2(new_n532), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n573), .A2(KEYINPUT86), .A3(new_n547), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(KEYINPUT87), .B(KEYINPUT39), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n525), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n538), .A2(new_n530), .A3(new_n540), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n578), .A2(KEYINPUT88), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT39), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n580), .B1(new_n578), .B2(KEYINPUT88), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n572), .A2(new_n579), .A3(new_n574), .A4(new_n581), .ZN(new_n582));
  AND3_X1   g381(.A1(new_n577), .A2(KEYINPUT40), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(KEYINPUT40), .B1(new_n577), .B2(new_n582), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n570), .A2(new_n585), .A3(new_n546), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n554), .A2(new_n556), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT90), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n499), .A2(new_n500), .A3(new_n332), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT89), .ZN(new_n590));
  OAI22_X1  g389(.A1(new_n455), .A2(new_n504), .B1(new_n503), .B2(new_n495), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(new_n295), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT89), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n499), .A2(new_n500), .A3(new_n593), .A4(new_n332), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n590), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT37), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT38), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT37), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n498), .A2(new_n502), .A3(new_n505), .A4(new_n598), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n596), .A2(new_n597), .A3(new_n599), .A4(new_n511), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n587), .A2(new_n588), .A3(new_n516), .A4(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n554), .A2(new_n556), .A3(new_n516), .ZN(new_n602));
  INV_X1    g401(.A(new_n600), .ZN(new_n603));
  OAI21_X1  g402(.A(KEYINPUT90), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n506), .A2(new_n598), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n599), .A2(new_n511), .ZN(new_n606));
  OAI21_X1  g405(.A(KEYINPUT38), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n601), .A2(new_n604), .A3(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n381), .A2(new_n586), .A3(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT36), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n478), .A2(new_n610), .A3(new_n487), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n488), .A2(KEYINPUT36), .A3(new_n489), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n378), .A2(new_n380), .A3(new_n559), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n609), .A2(new_n611), .A3(new_n612), .A4(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n283), .B1(new_n569), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(G99gat), .A2(G106gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT8), .ZN(new_n617));
  XNOR2_X1  g416(.A(KEYINPUT103), .B(G92gat), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n617), .B1(new_n618), .B2(G85gat), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(G99gat), .B(G106gat), .Z(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  OR2_X1    g421(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n623));
  NAND2_X1  g422(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n623), .A2(G85gat), .A3(G92gat), .A4(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g425(.A1(G85gat), .A2(G92gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n620), .A2(new_n622), .A3(new_n625), .A4(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n625), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n621), .B1(new_n630), .B2(new_n619), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT104), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n629), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  OAI211_X1 g432(.A(KEYINPUT104), .B(new_n621), .C1(new_n630), .C2(new_n619), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n245), .ZN(new_n636));
  NAND2_X1  g435(.A1(G232gat), .A2(G233gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT101), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT41), .ZN(new_n639));
  OR2_X1    g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n242), .A2(new_n237), .ZN(new_n641));
  OAI211_X1 g440(.A(new_n636), .B(new_n640), .C1(new_n641), .C2(new_n635), .ZN(new_n642));
  XOR2_X1   g441(.A(G190gat), .B(G218gat), .Z(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT105), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(KEYINPUT106), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT107), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n638), .A2(new_n639), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(new_n433), .ZN(new_n649));
  INV_X1    g448(.A(G162gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n646), .A2(new_n647), .A3(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT106), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n653), .B1(new_n642), .B2(new_n644), .ZN(new_n654));
  INV_X1    g453(.A(new_n651), .ZN(new_n655));
  OAI21_X1  g454(.A(KEYINPUT107), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n642), .A2(new_n644), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n645), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n652), .A2(new_n656), .A3(new_n645), .A4(new_n658), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT108), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT100), .ZN(new_n664));
  NAND2_X1  g463(.A1(G71gat), .A2(G78gat), .ZN(new_n665));
  INV_X1    g464(.A(G71gat), .ZN(new_n666));
  INV_X1    g465(.A(G78gat), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(G57gat), .B(G64gat), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT9), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n665), .B(new_n668), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n665), .B1(new_n668), .B2(new_n670), .ZN(new_n672));
  INV_X1    g471(.A(G57gat), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n508), .B1(new_n673), .B2(KEYINPUT98), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT97), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n676), .A2(G57gat), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT98), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n676), .A2(new_n678), .A3(G57gat), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n508), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n671), .B1(new_n675), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(KEYINPUT21), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n220), .A2(new_n664), .A3(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n683), .ZN(new_n685));
  OAI21_X1  g484(.A(KEYINPUT100), .B1(new_n219), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT21), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n681), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g487(.A(G127gat), .B(G155gat), .Z(new_n689));
  XOR2_X1   g488(.A(new_n688), .B(new_n689), .Z(new_n690));
  NAND3_X1  g489(.A1(new_n684), .A2(new_n686), .A3(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n690), .B1(new_n686), .B2(new_n684), .ZN(new_n693));
  OAI211_X1 g492(.A(G231gat), .B(G233gat), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n693), .ZN(new_n695));
  NAND2_X1  g494(.A1(G231gat), .A2(G233gat), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n695), .A2(new_n696), .A3(new_n691), .ZN(new_n697));
  XNOR2_X1  g496(.A(G183gat), .B(G211gat), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT20), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT99), .B(KEYINPUT19), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n694), .A2(new_n697), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n701), .B1(new_n694), .B2(new_n697), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n662), .A2(new_n663), .A3(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n704), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n660), .A2(new_n661), .ZN(new_n707));
  OAI21_X1  g506(.A(KEYINPUT108), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(G230gat), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n710), .A2(new_n493), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n633), .A2(new_n681), .A3(new_n634), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n682), .A2(new_n629), .A3(new_n631), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n712), .B1(new_n715), .B2(KEYINPUT10), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT10), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n713), .A2(KEYINPUT109), .A3(new_n714), .A4(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n635), .A2(KEYINPUT10), .A3(new_n682), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n711), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n715), .A2(new_n711), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(G120gat), .B(G148gat), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT110), .ZN(new_n726));
  INV_X1    g525(.A(G176gat), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(new_n286), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n724), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n729), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n722), .A2(new_n723), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n709), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n615), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n735), .A2(new_n557), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(new_n207), .ZN(G1324gat));
  INV_X1    g536(.A(new_n735), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n210), .B1(new_n738), .B2(new_n570), .ZN(new_n739));
  INV_X1    g538(.A(new_n570), .ZN(new_n740));
  NOR2_X1   g539(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n741));
  AND2_X1   g540(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n742));
  NOR4_X1   g541(.A1(new_n735), .A2(new_n740), .A3(new_n741), .A4(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(KEYINPUT42), .B1(new_n739), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(KEYINPUT42), .B2(new_n743), .ZN(G1325gat));
  NAND2_X1  g544(.A1(new_n612), .A2(new_n611), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n612), .A2(KEYINPUT111), .A3(new_n611), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n735), .A2(new_n202), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n738), .A2(new_n563), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n751), .B1(new_n202), .B2(new_n752), .ZN(G1326gat));
  NOR2_X1   g552(.A1(new_n735), .A2(new_n381), .ZN(new_n754));
  XOR2_X1   g553(.A(KEYINPUT43), .B(G22gat), .Z(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(G1327gat));
  AOI21_X1  g555(.A(new_n662), .B1(new_n569), .B2(new_n614), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n283), .A2(new_n704), .A3(new_n733), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n760), .A2(new_n223), .A3(new_n587), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT45), .ZN(new_n762));
  AND3_X1   g561(.A1(new_n372), .A2(new_n379), .A3(new_n376), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n379), .B1(new_n372), .B2(new_n376), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n563), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n567), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI22_X1  g566(.A1(new_n767), .A2(new_n564), .B1(new_n561), .B2(KEYINPUT35), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n608), .A2(new_n586), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n763), .A2(new_n764), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n613), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n771), .A2(new_n746), .ZN(new_n772));
  OAI211_X1 g571(.A(KEYINPUT44), .B(new_n707), .C1(new_n768), .C2(new_n772), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n612), .A2(KEYINPUT111), .A3(new_n611), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT111), .B1(new_n612), .B2(new_n611), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n613), .B(new_n609), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n662), .B1(new_n776), .B2(new_n569), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n773), .B(new_n758), .C1(new_n777), .C2(KEYINPUT44), .ZN(new_n778));
  OAI21_X1  g577(.A(G29gat), .B1(new_n778), .B2(new_n557), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n762), .A2(new_n779), .ZN(G1328gat));
  NOR3_X1   g579(.A1(new_n759), .A2(G36gat), .A3(new_n740), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT46), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(G36gat), .B1(new_n778), .B2(new_n740), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n781), .A2(new_n782), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(G1329gat));
  NAND2_X1  g585(.A1(new_n776), .A2(new_n569), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT44), .B1(new_n787), .B2(new_n707), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT44), .ZN(new_n789));
  AOI211_X1 g588(.A(new_n789), .B(new_n662), .C1(new_n569), .C2(new_n614), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n792));
  INV_X1    g591(.A(new_n750), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n791), .A2(new_n792), .A3(new_n793), .A4(new_n758), .ZN(new_n794));
  OAI21_X1  g593(.A(KEYINPUT112), .B1(new_n778), .B2(new_n750), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n794), .A2(G43gat), .A3(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(new_n563), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n759), .A2(G43gat), .A3(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT47), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(G43gat), .ZN(new_n802));
  INV_X1    g601(.A(new_n778), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n802), .B1(new_n803), .B2(new_n793), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n799), .B1(new_n804), .B2(new_n798), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n801), .A2(new_n805), .ZN(G1330gat));
  INV_X1    g605(.A(KEYINPUT48), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n807), .A2(KEYINPUT114), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n807), .A2(KEYINPUT114), .ZN(new_n809));
  OAI21_X1  g608(.A(G50gat), .B1(new_n778), .B2(new_n381), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n381), .A2(G50gat), .ZN(new_n811));
  XOR2_X1   g610(.A(new_n811), .B(KEYINPUT113), .Z(new_n812));
  NAND2_X1  g611(.A1(new_n760), .A2(new_n812), .ZN(new_n813));
  AOI211_X1 g612(.A(new_n808), .B(new_n809), .C1(new_n810), .C2(new_n813), .ZN(new_n814));
  AND4_X1   g613(.A1(KEYINPUT114), .A2(new_n810), .A3(new_n807), .A4(new_n813), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n814), .A2(new_n815), .ZN(G1331gat));
  INV_X1    g615(.A(new_n733), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n709), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n771), .B1(new_n748), .B2(new_n749), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n818), .B(new_n283), .C1(new_n819), .C2(new_n768), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n787), .A2(KEYINPUT115), .A3(new_n283), .A4(new_n818), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n824), .A2(new_n557), .ZN(new_n825));
  XNOR2_X1  g624(.A(KEYINPUT97), .B(G57gat), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n825), .B(new_n826), .ZN(G1332gat));
  OAI22_X1  g626(.A1(new_n824), .A2(new_n740), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n828));
  XNOR2_X1  g627(.A(KEYINPUT49), .B(G64gat), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n822), .A2(new_n570), .A3(new_n823), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(G1333gat));
  OAI21_X1  g630(.A(new_n666), .B1(new_n824), .B2(new_n797), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n822), .A2(G71gat), .A3(new_n793), .A4(new_n823), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT50), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n832), .A2(new_n836), .A3(new_n833), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(G1334gat));
  NOR2_X1   g637(.A1(new_n824), .A2(new_n381), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(new_n667), .ZN(G1335gat));
  NAND2_X1  g639(.A1(new_n283), .A2(new_n706), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(KEYINPUT116), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n777), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT51), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT51), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n777), .A2(new_n845), .A3(new_n842), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n844), .A2(new_n587), .A3(new_n733), .A4(new_n846), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n773), .B(new_n733), .C1(new_n777), .C2(KEYINPUT44), .ZN(new_n848));
  INV_X1    g647(.A(new_n842), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n557), .A2(new_n523), .ZN(new_n851));
  AOI22_X1  g650(.A1(new_n847), .A2(new_n523), .B1(new_n850), .B2(new_n851), .ZN(G1336gat));
  NOR2_X1   g651(.A1(new_n740), .A2(G92gat), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n844), .A2(new_n733), .A3(new_n846), .A4(new_n853), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n848), .A2(new_n740), .A3(new_n849), .ZN(new_n855));
  XOR2_X1   g654(.A(KEYINPUT103), .B(G92gat), .Z(new_n856));
  OAI21_X1  g655(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(KEYINPUT52), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT52), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n859), .B(new_n854), .C1(new_n855), .C2(new_n856), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(new_n860), .ZN(G1337gat));
  NOR2_X1   g660(.A1(new_n797), .A2(G99gat), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n844), .A2(new_n733), .A3(new_n846), .A4(new_n862), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n848), .A2(new_n750), .A3(new_n849), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n863), .B1(new_n864), .B2(new_n473), .ZN(G1338gat));
  NOR2_X1   g664(.A1(new_n381), .A2(G106gat), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n844), .A2(new_n733), .A3(new_n846), .A4(new_n866), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n848), .A2(new_n381), .A3(new_n849), .ZN(new_n868));
  INV_X1    g667(.A(G106gat), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  XNOR2_X1  g669(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n871), .B(new_n867), .C1(new_n868), .C2(new_n869), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(G1339gat));
  NOR2_X1   g674(.A1(new_n261), .A2(new_n263), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n244), .B1(new_n257), .B2(new_n243), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n269), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n273), .B1(new_n280), .B2(new_n270), .ZN(new_n879));
  INV_X1    g678(.A(new_n274), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n707), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n275), .A2(new_n661), .A3(new_n660), .A4(new_n281), .ZN(new_n883));
  INV_X1    g682(.A(new_n711), .ZN(new_n884));
  INV_X1    g683(.A(new_n720), .ZN(new_n885));
  AOI211_X1 g684(.A(new_n884), .B(new_n885), .C1(new_n716), .C2(new_n718), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n721), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n719), .A2(new_n720), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(new_n887), .A3(new_n884), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n729), .ZN(new_n891));
  OAI21_X1  g690(.A(KEYINPUT55), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n731), .B1(new_n721), .B2(new_n887), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT55), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT54), .B1(new_n889), .B2(new_n884), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n893), .B(new_n894), .C1(new_n721), .C2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n882), .A2(new_n732), .A3(new_n883), .A4(new_n897), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n662), .A2(new_n733), .A3(new_n275), .A4(new_n878), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n704), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  AND4_X1   g700(.A1(new_n708), .A2(new_n705), .A3(new_n817), .A4(new_n283), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n570), .A2(new_n557), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n906), .A2(new_n563), .A3(new_n381), .ZN(new_n907));
  OAI21_X1  g706(.A(G113gat), .B1(new_n907), .B2(new_n283), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n381), .A2(new_n490), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n282), .A2(new_n438), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(G1340gat));
  OAI21_X1  g711(.A(G120gat), .B1(new_n907), .B2(new_n817), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n733), .A2(new_n436), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n913), .B1(new_n910), .B2(new_n914), .ZN(G1341gat));
  INV_X1    g714(.A(new_n910), .ZN(new_n916));
  AOI21_X1  g715(.A(G127gat), .B1(new_n916), .B2(new_n704), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n907), .A2(new_n431), .A3(new_n706), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n917), .A2(new_n918), .ZN(G1342gat));
  NAND3_X1  g718(.A1(new_n916), .A2(new_n433), .A3(new_n707), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n920), .A2(KEYINPUT56), .ZN(new_n921));
  OAI21_X1  g720(.A(G134gat), .B1(new_n907), .B2(new_n662), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(KEYINPUT56), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(G1343gat));
  OAI21_X1  g723(.A(new_n770), .B1(new_n900), .B2(new_n902), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT57), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n925), .B(new_n926), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n750), .A2(new_n905), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n927), .A2(new_n282), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(G141gat), .ZN(new_n930));
  NAND2_X1  g729(.A1(KEYINPUT119), .A2(KEYINPUT58), .ZN(new_n931));
  INV_X1    g730(.A(new_n925), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n282), .A2(new_n300), .ZN(new_n934));
  XOR2_X1   g733(.A(new_n934), .B(KEYINPUT118), .Z(new_n935));
  OAI211_X1 g734(.A(new_n930), .B(new_n931), .C1(new_n933), .C2(new_n935), .ZN(new_n936));
  OR2_X1    g735(.A1(KEYINPUT119), .A2(KEYINPUT58), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n936), .B(new_n937), .ZN(G1344gat));
  INV_X1    g737(.A(new_n933), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n939), .A2(new_n309), .A3(new_n733), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT59), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n927), .A2(new_n928), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(new_n733), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n941), .B1(new_n943), .B2(G148gat), .ZN(new_n944));
  AOI211_X1 g743(.A(KEYINPUT59), .B(new_n309), .C1(new_n942), .C2(new_n733), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n940), .B1(new_n944), .B2(new_n945), .ZN(G1345gat));
  NAND2_X1  g745(.A1(new_n939), .A2(new_n704), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT120), .ZN(new_n948));
  INV_X1    g747(.A(G155gat), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n706), .A2(new_n949), .ZN(new_n950));
  AOI22_X1  g749(.A1(new_n948), .A2(new_n949), .B1(new_n942), .B2(new_n950), .ZN(G1346gat));
  NAND3_X1  g750(.A1(new_n939), .A2(new_n650), .A3(new_n707), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n942), .A2(new_n707), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n952), .B1(new_n953), .B2(new_n650), .ZN(G1347gat));
  NAND2_X1  g753(.A1(new_n909), .A2(new_n570), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT121), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n909), .A2(KEYINPUT121), .A3(new_n570), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n957), .A2(new_n557), .A3(new_n904), .A4(new_n958), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT122), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n960), .A2(new_n268), .A3(new_n282), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n740), .A2(new_n587), .ZN(new_n962));
  AOI21_X1  g761(.A(KEYINPUT123), .B1(new_n962), .B2(new_n563), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n963), .B1(new_n378), .B2(new_n380), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n962), .A2(KEYINPUT123), .A3(new_n563), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n964), .A2(new_n904), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g765(.A(G169gat), .B1(new_n966), .B2(new_n283), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n961), .A2(new_n967), .ZN(G1348gat));
  NOR3_X1   g767(.A1(new_n966), .A2(new_n727), .A3(new_n817), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n960), .A2(new_n733), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n969), .B1(new_n970), .B2(new_n727), .ZN(G1349gat));
  OAI21_X1  g770(.A(G183gat), .B1(new_n966), .B2(new_n706), .ZN(new_n972));
  INV_X1    g771(.A(new_n416), .ZN(new_n973));
  OR2_X1    g772(.A1(new_n959), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n972), .B1(new_n974), .B2(new_n706), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n975), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g775(.A1(new_n960), .A2(new_n417), .A3(new_n707), .ZN(new_n977));
  OAI21_X1  g776(.A(G190gat), .B1(new_n966), .B2(new_n662), .ZN(new_n978));
  XNOR2_X1  g777(.A(new_n978), .B(KEYINPUT61), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n977), .A2(new_n979), .ZN(G1351gat));
  OAI21_X1  g779(.A(new_n962), .B1(new_n774), .B2(new_n775), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(KEYINPUT124), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT124), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n750), .A2(new_n983), .A3(new_n962), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  INV_X1    g784(.A(new_n985), .ZN(new_n986));
  AND2_X1   g785(.A1(new_n986), .A2(new_n927), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n987), .A2(KEYINPUT125), .A3(new_n282), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n986), .A2(new_n282), .A3(new_n927), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT125), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n988), .A2(G197gat), .A3(new_n991), .ZN(new_n992));
  INV_X1    g791(.A(new_n981), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n993), .A2(new_n932), .ZN(new_n994));
  INV_X1    g793(.A(new_n994), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n995), .A2(new_n285), .A3(new_n282), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n992), .A2(new_n996), .ZN(G1352gat));
  NOR3_X1   g796(.A1(new_n994), .A2(G204gat), .A3(new_n817), .ZN(new_n998));
  XNOR2_X1  g797(.A(new_n998), .B(KEYINPUT62), .ZN(new_n999));
  AND2_X1   g798(.A1(new_n987), .A2(new_n733), .ZN(new_n1000));
  OAI21_X1  g799(.A(new_n999), .B1(new_n1000), .B2(new_n286), .ZN(G1353gat));
  NAND4_X1  g800(.A1(new_n927), .A2(new_n704), .A3(new_n982), .A4(new_n984), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1002), .A2(G211gat), .ZN(new_n1003));
  INV_X1    g802(.A(KEYINPUT63), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g804(.A(KEYINPUT127), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g806(.A1(new_n1002), .A2(KEYINPUT126), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n1008));
  INV_X1    g807(.A(KEYINPUT126), .ZN(new_n1009));
  OAI21_X1  g808(.A(new_n1009), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n1003), .A2(KEYINPUT127), .A3(new_n1004), .ZN(new_n1011));
  NAND4_X1  g810(.A1(new_n1007), .A2(new_n1008), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  OR3_X1    g811(.A1(new_n994), .A2(G211gat), .A3(new_n706), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n1012), .A2(new_n1013), .ZN(G1354gat));
  AOI21_X1  g813(.A(G218gat), .B1(new_n995), .B2(new_n707), .ZN(new_n1015));
  AND2_X1   g814(.A1(new_n707), .A2(G218gat), .ZN(new_n1016));
  AOI21_X1  g815(.A(new_n1015), .B1(new_n987), .B2(new_n1016), .ZN(G1355gat));
endmodule


