//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 0 1 1 1 1 1 0 1 1 1 0 1 1 0 1 0 0 0 0 1 1 1 0 0 0 1 1 0 0 0 0 0 0 1 0 0 0 0 1 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967;
  INV_X1    g000(.A(KEYINPUT23), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G128), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT23), .A3(G119), .ZN(new_n191));
  OAI211_X1 g005(.A(new_n189), .B(new_n191), .C1(G119), .C2(new_n190), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G110), .ZN(new_n193));
  XOR2_X1   g007(.A(G119), .B(G128), .Z(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT24), .B(G110), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT16), .ZN(new_n196));
  INV_X1    g010(.A(G140), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n197), .A3(G125), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(G125), .ZN(new_n199));
  INV_X1    g013(.A(G125), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G140), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n198), .B1(new_n202), .B2(new_n196), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(G125), .B(G140), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT16), .ZN(new_n207));
  AOI21_X1  g021(.A(G146), .B1(new_n207), .B2(new_n198), .ZN(new_n208));
  OAI221_X1 g022(.A(new_n193), .B1(new_n194), .B2(new_n195), .C1(new_n205), .C2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT71), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n210), .B1(new_n202), .B2(G146), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n206), .A2(KEYINPUT71), .A3(new_n204), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n207), .A2(G146), .A3(new_n198), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT72), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n194), .A2(new_n195), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n217), .B1(new_n192), .B2(G110), .ZN(new_n218));
  AND3_X1   g032(.A1(new_n215), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n216), .B1(new_n215), .B2(new_n218), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n209), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT22), .B(G137), .ZN(new_n222));
  INV_X1    g036(.A(G953), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n223), .A2(G221), .A3(G234), .ZN(new_n224));
  XOR2_X1   g038(.A(new_n222), .B(new_n224), .Z(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n221), .A2(new_n226), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n209), .B(new_n225), .C1(new_n219), .C2(new_n220), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(KEYINPUT25), .B1(new_n229), .B2(G902), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT25), .ZN(new_n231));
  INV_X1    g045(.A(G902), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n227), .A2(new_n231), .A3(new_n232), .A4(new_n228), .ZN(new_n233));
  INV_X1    g047(.A(G217), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n234), .B1(G234), .B2(new_n232), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n235), .B(KEYINPUT70), .ZN(new_n236));
  AND3_X1   g050(.A1(new_n230), .A2(new_n233), .A3(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n235), .A2(G902), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n227), .A2(new_n228), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT73), .ZN(new_n240));
  XNOR2_X1  g054(.A(new_n239), .B(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n237), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT28), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n204), .A2(G143), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT64), .ZN(new_n246));
  INV_X1    g060(.A(G143), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n246), .B1(new_n247), .B2(G146), .ZN(new_n248));
  NOR3_X1   g062(.A1(new_n204), .A2(KEYINPUT64), .A3(G143), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n245), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  AND2_X1   g064(.A1(KEYINPUT0), .A2(G128), .ZN(new_n251));
  NOR2_X1   g065(.A1(KEYINPUT0), .A2(G128), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n247), .A2(G146), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n245), .A2(new_n254), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n250), .A2(new_n253), .B1(new_n255), .B2(new_n251), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT11), .ZN(new_n257));
  INV_X1    g071(.A(G134), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n257), .B1(new_n258), .B2(G137), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(G137), .ZN(new_n260));
  INV_X1    g074(.A(G137), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n261), .A2(KEYINPUT11), .A3(G134), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n259), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G131), .ZN(new_n264));
  INV_X1    g078(.A(G131), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n259), .A2(new_n262), .A3(new_n265), .A4(new_n260), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n256), .A2(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n190), .A2(KEYINPUT1), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n255), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n245), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n254), .A2(KEYINPUT64), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n246), .A2(new_n247), .A3(G146), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n190), .B1(new_n245), .B2(KEYINPUT1), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n270), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n261), .A2(G134), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n258), .A2(G137), .ZN(new_n278));
  OAI21_X1  g092(.A(G131), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n266), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n268), .A2(new_n281), .ZN(new_n282));
  XOR2_X1   g096(.A(KEYINPUT2), .B(G113), .Z(new_n283));
  XNOR2_X1  g097(.A(G116), .B(G119), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n188), .A2(G116), .ZN(new_n286));
  INV_X1    g100(.A(G116), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G119), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(KEYINPUT2), .B(G113), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n285), .A2(KEYINPUT65), .A3(new_n291), .ZN(new_n292));
  OR3_X1    g106(.A1(new_n283), .A2(KEYINPUT65), .A3(new_n284), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n244), .B1(new_n282), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n282), .A2(new_n295), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT66), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n256), .A2(new_n298), .A3(new_n267), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n298), .B1(new_n256), .B2(new_n267), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n294), .B(new_n281), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n296), .B(new_n297), .C1(new_n301), .C2(new_n244), .ZN(new_n302));
  NOR2_X1   g116(.A1(G237), .A2(G953), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G210), .ZN(new_n304));
  XOR2_X1   g118(.A(new_n304), .B(KEYINPUT27), .Z(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT26), .B(G101), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n305), .B(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT69), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n308), .B(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n307), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT30), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n268), .A2(new_n281), .A3(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n281), .B1(new_n299), .B2(new_n300), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n313), .B1(new_n314), .B2(KEYINPUT30), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT67), .ZN(new_n316));
  NOR3_X1   g130(.A1(new_n315), .A2(new_n316), .A3(new_n294), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n301), .A2(new_n316), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n268), .A2(new_n281), .A3(new_n312), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n264), .A2(new_n266), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n255), .A2(new_n251), .ZN(new_n321));
  INV_X1    g135(.A(new_n253), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n321), .B1(new_n274), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT66), .B1(new_n320), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n256), .A2(new_n298), .A3(new_n267), .ZN(new_n325));
  AOI22_X1  g139(.A1(new_n324), .A2(new_n325), .B1(new_n276), .B2(new_n280), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n319), .B1(new_n326), .B2(new_n312), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n318), .B1(new_n327), .B2(new_n295), .ZN(new_n328));
  OAI211_X1 g142(.A(KEYINPUT68), .B(new_n311), .C1(new_n317), .C2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT31), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(KEYINPUT67), .B1(new_n326), .B2(new_n294), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n332), .B1(new_n315), .B2(new_n294), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n327), .A2(KEYINPUT67), .A3(new_n295), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n307), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(KEYINPUT68), .A3(KEYINPUT31), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n310), .B1(new_n331), .B2(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(G472), .A2(G902), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(KEYINPUT32), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n310), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n333), .A2(new_n334), .ZN(new_n342));
  AND4_X1   g156(.A1(KEYINPUT68), .A2(new_n342), .A3(KEYINPUT31), .A4(new_n311), .ZN(new_n343));
  AOI21_X1  g157(.A(KEYINPUT31), .B1(new_n335), .B2(KEYINPUT68), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n341), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT32), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(new_n346), .A3(new_n338), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n340), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G472), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n314), .A2(new_n295), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n301), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(KEYINPUT28), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n352), .A2(new_n296), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT29), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n307), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(G902), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n333), .A2(new_n334), .A3(new_n307), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n357), .B(new_n354), .C1(new_n307), .C2(new_n302), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n349), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n243), .B1(new_n348), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G101), .ZN(new_n362));
  INV_X1    g176(.A(G107), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n363), .A2(G104), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(G104), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n362), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT77), .ZN(new_n368));
  INV_X1    g182(.A(G104), .ZN(new_n369));
  OAI21_X1  g183(.A(KEYINPUT3), .B1(new_n369), .B2(G107), .ZN(new_n370));
  XNOR2_X1  g184(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n368), .B(new_n370), .C1(new_n371), .C2(new_n366), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT3), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT76), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT76), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT3), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n366), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(KEYINPUT77), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n372), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n364), .A2(G101), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n367), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(G113), .B1(new_n286), .B2(KEYINPUT5), .ZN(new_n383));
  OR2_X1    g197(.A1(new_n383), .A2(KEYINPUT85), .ZN(new_n384));
  AOI22_X1  g198(.A1(new_n383), .A2(KEYINPUT85), .B1(new_n284), .B2(KEYINPUT5), .ZN(new_n385));
  AOI22_X1  g199(.A1(new_n384), .A2(new_n385), .B1(new_n284), .B2(new_n283), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(KEYINPUT86), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT86), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n382), .A2(new_n389), .A3(new_n386), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n383), .B1(KEYINPUT5), .B2(new_n284), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n391), .B1(new_n284), .B2(new_n283), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n388), .B(new_n390), .C1(new_n382), .C2(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(G110), .B(G122), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n394), .B(KEYINPUT8), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n366), .B1(new_n374), .B2(new_n376), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n370), .A2(new_n368), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NOR3_X1   g212(.A1(new_n371), .A2(new_n368), .A3(new_n366), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n365), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n362), .A2(KEYINPUT4), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n294), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n381), .B1(new_n398), .B2(new_n399), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n364), .B1(new_n372), .B2(new_n379), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n403), .B(KEYINPUT4), .C1(new_n404), .C2(new_n362), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n402), .A2(new_n405), .B1(new_n382), .B2(new_n392), .ZN(new_n406));
  AOI22_X1  g220(.A1(new_n393), .A2(new_n395), .B1(new_n394), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(KEYINPUT84), .B1(new_n256), .B2(new_n200), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n270), .B(new_n200), .C1(new_n274), .C2(new_n275), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT84), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n323), .A2(new_n410), .A3(G125), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n408), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G224), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n413), .A2(G953), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT87), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(KEYINPUT7), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n417), .B(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(G902), .B1(new_n407), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT6), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n421), .B1(new_n406), .B2(new_n394), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n402), .A2(new_n405), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n382), .A2(new_n392), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n394), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n425), .A2(new_n421), .A3(new_n426), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n412), .B(new_n414), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n420), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(G210), .B1(G237), .B2(G902), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n420), .A2(new_n431), .A3(new_n433), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(G214), .B1(G237), .B2(G902), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT89), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n441), .B1(new_n205), .B2(new_n208), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n303), .A2(G214), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n247), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n303), .A2(G143), .A3(G214), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n265), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT17), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n444), .A2(new_n265), .A3(new_n445), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n203), .A2(new_n204), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(KEYINPUT89), .A3(new_n214), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n446), .A2(KEYINPUT17), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n442), .A2(new_n450), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(G113), .B(G122), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(new_n369), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n444), .A2(new_n445), .ZN(new_n457));
  AND2_X1   g271(.A1(KEYINPUT18), .A2(G131), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(KEYINPUT18), .A2(G131), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n444), .A2(new_n445), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n211), .A2(new_n212), .B1(G146), .B2(new_n202), .ZN(new_n463));
  OR2_X1    g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n454), .A2(new_n456), .A3(new_n464), .ZN(new_n465));
  AND2_X1   g279(.A1(KEYINPUT88), .A2(KEYINPUT19), .ZN(new_n466));
  NOR2_X1   g280(.A1(KEYINPUT88), .A2(KEYINPUT19), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n206), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n468), .B1(new_n206), .B2(new_n467), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n214), .B1(new_n469), .B2(G146), .ZN(new_n470));
  INV_X1    g284(.A(new_n449), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n471), .A2(new_n446), .ZN(new_n472));
  OAI22_X1  g286(.A1(new_n470), .A2(new_n472), .B1(new_n463), .B2(new_n462), .ZN(new_n473));
  INV_X1    g287(.A(new_n456), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n465), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT20), .ZN(new_n477));
  INV_X1    g291(.A(G475), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n476), .A2(new_n477), .A3(new_n478), .A4(new_n232), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n465), .A2(new_n475), .A3(KEYINPUT90), .ZN(new_n480));
  AOI21_X1  g294(.A(KEYINPUT90), .B1(new_n465), .B2(new_n475), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n478), .A2(new_n232), .ZN(new_n482));
  NOR3_X1   g296(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n479), .B1(new_n483), .B2(new_n477), .ZN(new_n484));
  INV_X1    g298(.A(new_n465), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n456), .B1(new_n454), .B2(new_n464), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n232), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT92), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(KEYINPUT91), .B(G475), .ZN(new_n490));
  OAI211_X1 g304(.A(KEYINPUT92), .B(new_n232), .C1(new_n485), .C2(new_n486), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n484), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(G478), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n494), .A2(KEYINPUT15), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n247), .A2(G128), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n190), .A2(G143), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G134), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n496), .A2(new_n497), .A3(new_n258), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT93), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT93), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n499), .A2(new_n503), .A3(new_n500), .ZN(new_n504));
  OR2_X1    g318(.A1(new_n287), .A2(G122), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n287), .A2(G122), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n505), .B(new_n506), .C1(KEYINPUT14), .C2(new_n363), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n506), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n505), .A2(KEYINPUT14), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(new_n509), .A3(G107), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n502), .A2(new_n504), .A3(new_n507), .A4(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT13), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n496), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n497), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n496), .A2(new_n512), .ZN(new_n515));
  OAI21_X1  g329(.A(G134), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n508), .A2(new_n363), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n505), .A2(new_n506), .A3(G107), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n516), .A2(new_n517), .A3(new_n518), .A4(new_n500), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT9), .B(G234), .ZN(new_n520));
  NOR3_X1   g334(.A1(new_n520), .A2(new_n234), .A3(G953), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n511), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n521), .B1(new_n511), .B2(new_n519), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n232), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT94), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n495), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n525), .A2(new_n526), .ZN(new_n528));
  INV_X1    g342(.A(new_n524), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n522), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n530), .A2(KEYINPUT94), .A3(new_n232), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n527), .B1(new_n532), .B2(new_n495), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(G234), .A2(G237), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n535), .A2(G952), .A3(new_n223), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n535), .A2(G902), .A3(G953), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT21), .B(G898), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR3_X1   g353(.A1(new_n493), .A2(new_n534), .A3(new_n539), .ZN(new_n540));
  AND2_X1   g354(.A1(new_n440), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n245), .A2(KEYINPUT79), .A3(KEYINPUT1), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(G128), .ZN(new_n543));
  AOI21_X1  g357(.A(KEYINPUT79), .B1(new_n245), .B2(KEYINPUT1), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n270), .B1(new_n545), .B2(new_n255), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n382), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT10), .ZN(new_n548));
  AND2_X1   g362(.A1(new_n276), .A2(KEYINPUT10), .ZN(new_n549));
  AOI22_X1  g363(.A1(new_n547), .A2(new_n548), .B1(new_n549), .B2(new_n382), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT78), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n323), .B1(new_n400), .B2(new_n401), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n405), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n551), .B1(new_n405), .B2(new_n552), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n320), .B(new_n550), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT80), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n405), .A2(new_n552), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT78), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n405), .A2(new_n552), .A3(new_n551), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT80), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n560), .A2(new_n561), .A3(new_n320), .A4(new_n550), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n556), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n320), .B1(new_n560), .B2(new_n550), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(G110), .B(G140), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n223), .A2(G227), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n567), .B(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n569), .B(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n566), .A2(KEYINPUT82), .A3(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT82), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n564), .B1(new_n562), .B2(new_n556), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n574), .B1(new_n575), .B2(new_n571), .ZN(new_n576));
  OR2_X1    g390(.A1(new_n382), .A2(new_n276), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n320), .B1(new_n577), .B2(new_n547), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(KEYINPUT12), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n563), .A2(new_n571), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n573), .A2(new_n576), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(G469), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(new_n582), .A3(new_n232), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n582), .A2(new_n232), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT81), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n563), .A2(new_n571), .A3(new_n565), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n571), .B1(new_n563), .B2(new_n579), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n563), .A2(new_n571), .A3(new_n565), .ZN(new_n590));
  OR2_X1    g404(.A1(new_n578), .A2(KEYINPUT12), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n578), .A2(KEYINPUT12), .ZN(new_n592));
  AOI22_X1  g406(.A1(new_n556), .A2(new_n562), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n590), .B(KEYINPUT81), .C1(new_n571), .C2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n589), .A2(G469), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n583), .A2(new_n585), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(G221), .ZN(new_n597));
  INV_X1    g411(.A(new_n520), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n597), .B1(new_n598), .B2(new_n232), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n596), .A2(KEYINPUT83), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(KEYINPUT83), .B1(new_n596), .B2(new_n600), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n361), .B(new_n541), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(G101), .ZN(G3));
  NAND2_X1  g418(.A1(new_n525), .A2(new_n494), .ZN(new_n605));
  OR2_X1    g419(.A1(new_n523), .A2(KEYINPUT96), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n523), .A2(KEYINPUT96), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n606), .A2(KEYINPUT33), .A3(new_n607), .ZN(new_n608));
  XOR2_X1   g422(.A(new_n524), .B(KEYINPUT95), .Z(new_n609));
  INV_X1    g423(.A(new_n530), .ZN(new_n610));
  OAI22_X1  g424(.A1(new_n608), .A2(new_n609), .B1(KEYINPUT33), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n232), .A2(G478), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n605), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n493), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n349), .B1(new_n345), .B2(new_n232), .ZN(new_n616));
  INV_X1    g430(.A(new_n539), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n437), .A2(new_n438), .A3(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n337), .A2(new_n339), .ZN(new_n619));
  NOR4_X1   g433(.A1(new_n616), .A2(new_n618), .A3(new_n619), .A4(new_n243), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n615), .B(new_n620), .C1(new_n601), .C2(new_n602), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT34), .B(G104), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT97), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n621), .B(new_n623), .ZN(G6));
  OR2_X1    g438(.A1(new_n601), .A2(new_n602), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n483), .B(new_n477), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n626), .A2(new_n492), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n625), .A2(new_n534), .A3(new_n620), .A4(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT35), .B(G107), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G9));
  XNOR2_X1  g444(.A(new_n221), .B(KEYINPUT98), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n226), .A2(KEYINPUT36), .ZN(new_n632));
  XOR2_X1   g446(.A(new_n631), .B(new_n632), .Z(new_n633));
  AOI21_X1  g447(.A(new_n237), .B1(new_n633), .B2(new_n238), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n616), .A2(new_n619), .A3(new_n634), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n635), .B(new_n541), .C1(new_n601), .C2(new_n602), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT37), .B(G110), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G12));
  AOI21_X1  g452(.A(new_n359), .B1(new_n340), .B2(new_n347), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n639), .A2(new_n439), .A3(new_n634), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n625), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n627), .A2(new_n534), .ZN(new_n642));
  INV_X1    g456(.A(G900), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n537), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n536), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n641), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G128), .ZN(G30));
  XNOR2_X1  g464(.A(new_n646), .B(KEYINPUT39), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n625), .A2(new_n651), .ZN(new_n652));
  OR2_X1    g466(.A1(new_n652), .A2(KEYINPUT40), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(KEYINPUT40), .ZN(new_n654));
  INV_X1    g468(.A(new_n348), .ZN(new_n655));
  INV_X1    g469(.A(new_n335), .ZN(new_n656));
  INV_X1    g470(.A(new_n351), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n656), .B1(new_n311), .B2(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n349), .B1(new_n658), .B2(new_n232), .ZN(new_n659));
  OR2_X1    g473(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n634), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n437), .B(KEYINPUT38), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n533), .B1(new_n484), .B2(new_n492), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n663), .A2(new_n438), .A3(new_n664), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n661), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n653), .A2(new_n654), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G143), .ZN(G45));
  NOR2_X1   g482(.A1(new_n614), .A2(new_n647), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n641), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT99), .B(G146), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G48));
  INV_X1    g486(.A(new_n361), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n581), .A2(new_n582), .A3(new_n232), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n582), .B1(new_n581), .B2(new_n232), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n674), .A2(new_n675), .A3(new_n599), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n618), .A2(new_n614), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT41), .B(G113), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G15));
  NOR2_X1   g496(.A1(new_n642), .A2(new_n618), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n678), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(new_n287), .ZN(G18));
  NAND2_X1  g499(.A1(new_n348), .A2(new_n360), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n540), .A3(new_n662), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n674), .A2(new_n675), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT100), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n688), .A2(new_n689), .A3(new_n600), .A4(new_n440), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n581), .A2(new_n232), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(G469), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n692), .A2(new_n600), .A3(new_n583), .A4(new_n440), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(KEYINPUT100), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n687), .B1(new_n690), .B2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(new_n188), .ZN(G21));
  OAI21_X1  g510(.A(G472), .B1(new_n337), .B2(G902), .ZN(new_n697));
  OAI21_X1  g511(.A(KEYINPUT101), .B1(new_n237), .B2(new_n241), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n239), .B(KEYINPUT73), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n230), .A2(new_n233), .A3(new_n236), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT101), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n343), .A2(new_n344), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n353), .A2(new_n311), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n338), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n697), .A2(new_n703), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT102), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT102), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n697), .A2(new_n703), .A3(new_n706), .A4(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n437), .A2(new_n438), .A3(new_n617), .A4(new_n664), .ZN(new_n712));
  NOR4_X1   g526(.A1(new_n674), .A2(new_n675), .A3(new_n712), .A4(new_n599), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G122), .ZN(G24));
  NAND2_X1  g529(.A1(new_n690), .A2(new_n694), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n697), .A2(new_n706), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n662), .ZN(new_n718));
  INV_X1    g532(.A(new_n669), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  XOR2_X1   g535(.A(KEYINPUT103), .B(G125), .Z(new_n722));
  XNOR2_X1  g536(.A(new_n721), .B(new_n722), .ZN(G27));
  NOR2_X1   g537(.A1(new_n587), .A2(new_n588), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n584), .B1(new_n724), .B2(G469), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n583), .A2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n438), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n599), .A2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n437), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT42), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n731), .A2(new_n732), .A3(new_n719), .ZN(new_n733));
  AOI21_X1  g547(.A(KEYINPUT104), .B1(new_n686), .B2(new_n703), .ZN(new_n734));
  INV_X1    g548(.A(new_n703), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT104), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n639), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n733), .B1(new_n734), .B2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n730), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n739), .B1(new_n583), .B2(new_n725), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n361), .A2(new_n740), .A3(new_n669), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n732), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G131), .ZN(G33));
  AND3_X1   g558(.A1(new_n361), .A2(new_n740), .A3(new_n648), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n258), .ZN(G36));
  AOI21_X1  g560(.A(KEYINPUT45), .B1(new_n589), .B2(new_n594), .ZN(new_n747));
  AOI211_X1 g561(.A(new_n582), .B(new_n747), .C1(KEYINPUT45), .C2(new_n724), .ZN(new_n748));
  OR2_X1    g562(.A1(new_n748), .A2(new_n584), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT46), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n674), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n751), .B1(new_n750), .B2(new_n749), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n600), .A3(new_n651), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n613), .A2(new_n484), .A3(new_n492), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT105), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XOR2_X1   g570(.A(new_n756), .B(KEYINPUT43), .Z(new_n757));
  NOR2_X1   g571(.A1(new_n616), .A2(new_n619), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n757), .A2(new_n758), .A3(new_n634), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n759), .A2(KEYINPUT44), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n753), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n437), .A2(new_n727), .ZN(new_n762));
  INV_X1    g576(.A(new_n759), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT44), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  XOR2_X1   g579(.A(new_n765), .B(KEYINPUT106), .Z(new_n766));
  OR2_X1    g580(.A1(new_n761), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G137), .ZN(G39));
  NAND4_X1  g582(.A1(new_n639), .A2(new_n243), .A3(new_n669), .A4(new_n762), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(KEYINPUT107), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n752), .A2(KEYINPUT47), .A3(new_n600), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(KEYINPUT47), .B1(new_n752), .B2(new_n600), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n770), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G140), .ZN(G42));
  XNOR2_X1  g589(.A(new_n688), .B(KEYINPUT49), .ZN(new_n776));
  NOR4_X1   g590(.A1(new_n663), .A2(new_n735), .A3(new_n729), .A4(new_n754), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n776), .A2(new_n661), .A3(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n688), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(new_n739), .ZN(new_n780));
  AND4_X1   g594(.A1(new_n242), .A2(new_n661), .A3(new_n536), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n615), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n782), .A2(G952), .A3(new_n223), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n757), .A2(new_n645), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n784), .A2(new_n780), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n734), .A2(new_n737), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  XOR2_X1   g602(.A(new_n788), .B(KEYINPUT48), .Z(new_n789));
  AND2_X1   g603(.A1(new_n784), .A2(new_n711), .ZN(new_n790));
  AOI211_X1 g604(.A(new_n783), .B(new_n789), .C1(new_n716), .C2(new_n790), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n677), .A2(new_n438), .A3(new_n663), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  XOR2_X1   g607(.A(new_n793), .B(KEYINPUT50), .Z(new_n794));
  NOR2_X1   g608(.A1(new_n493), .A2(new_n613), .ZN(new_n795));
  INV_X1    g609(.A(new_n718), .ZN(new_n796));
  AOI22_X1  g610(.A1(new_n781), .A2(new_n795), .B1(new_n785), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n773), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n799), .B(new_n771), .C1(new_n600), .C2(new_n779), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n790), .A2(new_n762), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n798), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n791), .B1(new_n803), .B2(KEYINPUT51), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n805));
  OAI221_X1 g619(.A(new_n640), .B1(new_n648), .B2(new_n669), .C1(new_n601), .C2(new_n602), .ZN(new_n806));
  INV_X1    g620(.A(new_n664), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n439), .A2(new_n807), .ZN(new_n808));
  AND4_X1   g622(.A1(new_n600), .A2(new_n726), .A3(new_n646), .A4(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n660), .A2(new_n809), .A3(new_n634), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n806), .A2(new_n721), .A3(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n806), .A2(new_n721), .A3(KEYINPUT52), .A4(new_n810), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(KEYINPUT53), .B1(new_n815), .B2(KEYINPUT110), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n493), .A2(new_n533), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n620), .B(new_n817), .C1(new_n601), .C2(new_n602), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT109), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n636), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n819), .B1(new_n636), .B2(new_n818), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n603), .A2(new_n621), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n687), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n716), .A2(new_n824), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n361), .B(new_n676), .C1(new_n679), .C2(new_n683), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n825), .A2(KEYINPUT108), .A3(new_n714), .A4(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT108), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n714), .A2(new_n826), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n828), .B1(new_n829), .B2(new_n695), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n745), .B1(new_n738), .B2(new_n742), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n762), .A2(new_n533), .A3(new_n627), .A4(new_n646), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n639), .A2(new_n833), .A3(new_n634), .ZN(new_n834));
  AOI22_X1  g648(.A1(new_n625), .A2(new_n834), .B1(new_n720), .B2(new_n740), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n815), .A2(new_n823), .A3(new_n831), .A4(new_n836), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n816), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n816), .A2(new_n837), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n805), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT53), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n829), .A2(new_n695), .A3(new_n842), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n823), .A2(new_n836), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(KEYINPUT54), .B1(new_n844), .B2(new_n815), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n827), .A2(new_n830), .A3(new_n832), .A4(new_n835), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n636), .A2(new_n818), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT109), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n636), .A2(new_n818), .A3(new_n819), .ZN(new_n849));
  INV_X1    g663(.A(new_n822), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n846), .A2(new_n851), .ZN(new_n852));
  AOI211_X1 g666(.A(KEYINPUT111), .B(KEYINPUT53), .C1(new_n852), .C2(new_n815), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT111), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n854), .B1(new_n837), .B2(new_n842), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n845), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n841), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n803), .A2(KEYINPUT51), .ZN(new_n858));
  OR2_X1    g672(.A1(new_n858), .A2(KEYINPUT112), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(KEYINPUT112), .ZN(new_n860));
  AOI211_X1 g674(.A(new_n804), .B(new_n857), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(G952), .A2(G953), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n778), .B1(new_n861), .B2(new_n862), .ZN(G75));
  NAND2_X1  g677(.A1(new_n844), .A2(new_n815), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n864), .B1(new_n853), .B2(new_n855), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n865), .A2(G210), .A3(G902), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT56), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n866), .A2(KEYINPUT114), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n428), .A2(new_n429), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(new_n430), .ZN(new_n870));
  XNOR2_X1  g684(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n870), .B(new_n871), .Z(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n868), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n866), .A2(KEYINPUT114), .A3(new_n867), .A4(new_n872), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n223), .A2(G952), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n874), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT115), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n874), .A2(KEYINPUT115), .A3(new_n875), .A4(new_n877), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(G51));
  INV_X1    g696(.A(KEYINPUT116), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n856), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n865), .A2(KEYINPUT54), .ZN(new_n885));
  OAI211_X1 g699(.A(KEYINPUT116), .B(new_n845), .C1(new_n853), .C2(new_n855), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n584), .B(KEYINPUT57), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT117), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n887), .A2(KEYINPUT117), .A3(new_n888), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n891), .A2(new_n581), .A3(new_n892), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n865), .A2(G902), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n748), .B(KEYINPUT118), .Z(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n876), .B1(new_n893), .B2(new_n896), .ZN(G54));
  NAND3_X1  g711(.A1(new_n894), .A2(KEYINPUT58), .A3(G475), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n480), .A2(new_n481), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n898), .A2(new_n900), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n901), .A2(new_n902), .A3(new_n876), .ZN(G60));
  NAND2_X1  g717(.A1(G478), .A2(G902), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT59), .Z(new_n905));
  NOR2_X1   g719(.A1(new_n611), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n876), .B1(new_n887), .B2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT119), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n841), .A2(new_n856), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n611), .B1(new_n910), .B2(new_n905), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n911), .B1(new_n907), .B2(new_n908), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n909), .A2(new_n912), .ZN(G63));
  NAND2_X1  g727(.A1(G217), .A2(G902), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT60), .Z(new_n915));
  NAND2_X1  g729(.A1(new_n865), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n876), .B1(new_n916), .B2(new_n229), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT120), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT61), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n865), .A2(new_n633), .A3(new_n915), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n919), .B(new_n921), .ZN(G66));
  OAI21_X1  g736(.A(G953), .B1(new_n538), .B2(new_n413), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n823), .A2(new_n831), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n923), .B1(new_n924), .B2(G953), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n869), .B1(G898), .B2(new_n223), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT122), .Z(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT121), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n925), .B(new_n928), .ZN(G69));
  AOI21_X1  g743(.A(new_n223), .B1(G227), .B2(G900), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n315), .B(new_n469), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n762), .B1(new_n817), .B2(new_n615), .ZN(new_n932));
  OR3_X1    g746(.A1(new_n652), .A2(new_n673), .A3(new_n932), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n767), .A2(new_n774), .A3(new_n933), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n806), .A2(new_n721), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n667), .A2(new_n935), .ZN(new_n936));
  OR2_X1    g750(.A1(new_n936), .A2(KEYINPUT62), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(KEYINPUT62), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n934), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n931), .B1(new_n939), .B2(new_n223), .ZN(new_n940));
  NAND2_X1  g754(.A1(G900), .A2(G953), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n931), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n787), .A2(new_n808), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n767), .B1(new_n753), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n774), .A2(new_n935), .A3(new_n832), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n942), .B1(new_n946), .B2(new_n223), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n930), .B1(new_n940), .B2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n947), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n930), .B(KEYINPUT124), .Z(new_n950));
  OAI211_X1 g764(.A(new_n949), .B(new_n950), .C1(new_n940), .C2(KEYINPUT123), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n940), .A2(KEYINPUT123), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n948), .B1(new_n951), .B2(new_n952), .ZN(G72));
  XOR2_X1   g767(.A(new_n342), .B(KEYINPUT125), .Z(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n934), .A2(new_n924), .A3(new_n937), .A4(new_n938), .ZN(new_n956));
  NAND2_X1  g770(.A1(G472), .A2(G902), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT63), .Z(new_n958));
  AOI211_X1 g772(.A(new_n307), .B(new_n955), .C1(new_n956), .C2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n958), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n946), .B2(new_n924), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n955), .A2(new_n307), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT126), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n877), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n960), .B1(new_n656), .B2(new_n357), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT127), .Z(new_n966));
  AOI21_X1  g780(.A(new_n966), .B1(new_n838), .B2(new_n839), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n959), .A2(new_n964), .A3(new_n967), .ZN(G57));
endmodule


