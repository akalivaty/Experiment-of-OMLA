//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 0 0 0 1 0 0 1 1 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 1 1 1 0 0 1 1 1 1 0 0 0 0 1 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n559, new_n561, new_n562, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n581, new_n582,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n622, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1233, new_n1234, new_n1235;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT65), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT66), .Z(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n462), .A2(G137), .A3(new_n461), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n465), .A2(new_n470), .ZN(G160));
  NAND2_X1  g046(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(new_n461), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n461), .A2(G112), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n475), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n481), .A2(KEYINPUT67), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n481), .A2(KEYINPUT67), .ZN(new_n483));
  OAI221_X1 g058(.A(new_n477), .B1(new_n478), .B2(new_n479), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  XOR2_X1   g059(.A(new_n484), .B(KEYINPUT68), .Z(G162));
  NAND4_X1  g060(.A1(new_n472), .A2(new_n474), .A3(G138), .A4(new_n461), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT4), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n462), .A2(new_n488), .A3(G138), .A4(new_n461), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  AND4_X1   g065(.A1(G126), .A2(new_n472), .A3(new_n474), .A4(G2105), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n493), .B1(new_n461), .B2(G114), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n495), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n492), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n491), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n490), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(new_n507), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n505), .A2(new_n512), .A3(G88), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(G50), .A3(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT70), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n513), .A2(new_n514), .A3(KEYINPUT70), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n508), .B1(new_n517), .B2(new_n518), .ZN(G166));
  INV_X1    g094(.A(new_n504), .ZN(new_n520));
  NOR2_X1   g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(G63), .A2(G651), .ZN(new_n523));
  OR3_X1    g098(.A1(new_n522), .A2(KEYINPUT71), .A3(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n503), .A2(new_n504), .B1(new_n510), .B2(new_n511), .ZN(new_n525));
  XOR2_X1   g100(.A(KEYINPUT74), .B(G89), .Z(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g102(.A(KEYINPUT71), .B1(new_n522), .B2(new_n523), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n524), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT73), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT7), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n512), .A2(G543), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT72), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n502), .B1(new_n510), .B2(new_n511), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(KEYINPUT72), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  AOI211_X1 g114(.A(new_n529), .B(new_n533), .C1(G51), .C2(new_n539), .ZN(G168));
  XNOR2_X1  g115(.A(KEYINPUT75), .B(G52), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(G77), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G64), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n522), .B2(new_n544), .ZN(new_n545));
  XNOR2_X1  g120(.A(KEYINPUT76), .B(G90), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n545), .A2(G651), .B1(new_n525), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n542), .A2(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  NAND2_X1  g124(.A1(new_n539), .A2(G43), .ZN(new_n550));
  NAND2_X1  g125(.A1(G68), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G56), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n522), .B2(new_n552), .ZN(new_n553));
  XOR2_X1   g128(.A(KEYINPUT77), .B(G81), .Z(new_n554));
  AOI22_X1  g129(.A1(new_n553), .A2(G651), .B1(new_n525), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  AND3_X1   g133(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G36), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n562), .ZN(G188));
  INV_X1    g138(.A(KEYINPUT78), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n505), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n565), .B2(new_n507), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n522), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n569), .A2(KEYINPUT78), .A3(G651), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT9), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n537), .A2(new_n572), .A3(G53), .ZN(new_n573));
  INV_X1    g148(.A(new_n511), .ZN(new_n574));
  NOR2_X1   g149(.A1(KEYINPUT6), .A2(G651), .ZN(new_n575));
  OAI211_X1 g150(.A(G53), .B(G543), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(KEYINPUT9), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n573), .A2(new_n577), .B1(new_n525), .B2(G91), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n571), .A2(new_n578), .ZN(G299));
  INV_X1    g154(.A(G168), .ZN(G286));
  INV_X1    g155(.A(new_n518), .ZN(new_n581));
  AOI21_X1  g156(.A(KEYINPUT70), .B1(new_n513), .B2(new_n514), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n581), .A2(new_n582), .B1(new_n507), .B2(new_n506), .ZN(G303));
  OAI21_X1  g158(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n537), .A2(G49), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n505), .A2(new_n512), .A3(G87), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT79), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n584), .A2(new_n585), .A3(new_n586), .A4(KEYINPUT79), .ZN(new_n590));
  AND2_X1   g165(.A1(new_n589), .A2(new_n590), .ZN(G288));
  AOI22_X1  g166(.A1(new_n525), .A2(G86), .B1(new_n537), .B2(G48), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n593), .B(KEYINPUT80), .ZN(new_n594));
  INV_X1    g169(.A(G61), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n595), .B1(new_n503), .B2(new_n504), .ZN(new_n596));
  OAI21_X1  g171(.A(G651), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n592), .A2(new_n597), .ZN(G305));
  NAND2_X1  g173(.A1(G72), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G60), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n522), .B2(new_n600), .ZN(new_n601));
  XNOR2_X1  g176(.A(KEYINPUT81), .B(G85), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n601), .A2(G651), .B1(new_n525), .B2(new_n602), .ZN(new_n603));
  AND2_X1   g178(.A1(new_n536), .A2(new_n538), .ZN(new_n604));
  INV_X1    g179(.A(G47), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(G301), .A2(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(G79), .A2(G543), .ZN(new_n608));
  INV_X1    g183(.A(G66), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n522), .B2(new_n609), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n539), .A2(G54), .B1(G651), .B2(new_n610), .ZN(new_n611));
  AND3_X1   g186(.A1(new_n505), .A2(new_n512), .A3(G92), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT10), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n607), .B1(new_n615), .B2(G868), .ZN(G284));
  XOR2_X1   g191(.A(G284), .B(KEYINPUT82), .Z(G321));
  NAND2_X1  g192(.A1(G286), .A2(G868), .ZN(new_n618));
  INV_X1    g193(.A(G299), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(G868), .B2(new_n619), .ZN(G297));
  OAI21_X1  g195(.A(new_n618), .B1(G868), .B2(new_n619), .ZN(G280));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n615), .B1(new_n622), .B2(G860), .ZN(G148));
  NAND2_X1  g198(.A1(new_n615), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G868), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G868), .B2(new_n557), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n476), .A2(G123), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT83), .Z(new_n629));
  OR2_X1    g204(.A1(G99), .A2(G2105), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n630), .B(G2104), .C1(G111), .C2(new_n461), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n480), .A2(G135), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n629), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(G2096), .Z(new_n634));
  NAND2_X1  g209(.A1(new_n480), .A2(G2104), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT13), .Z(new_n637));
  OR2_X1    g212(.A1(new_n637), .A2(G2100), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(G2100), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n634), .A2(new_n638), .A3(new_n639), .ZN(G156));
  XNOR2_X1  g215(.A(G2427), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(KEYINPUT14), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT84), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(G1341), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n647), .A2(G1341), .ZN(new_n650));
  OAI21_X1  g225(.A(G1348), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2451), .B(G2454), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n653), .B(new_n654), .Z(new_n655));
  OR2_X1    g230(.A1(new_n647), .A2(G1341), .ZN(new_n656));
  INV_X1    g231(.A(G1348), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n656), .A2(new_n657), .A3(new_n648), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n651), .A2(new_n655), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(G14), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n655), .B1(new_n651), .B2(new_n658), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(G401));
  XNOR2_X1  g237(.A(G2084), .B(G2090), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT85), .Z(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2072), .B(G2078), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n664), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n667), .A2(KEYINPUT86), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(KEYINPUT86), .ZN(new_n669));
  INV_X1    g244(.A(new_n665), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n666), .B(KEYINPUT17), .Z(new_n671));
  OAI211_X1 g246(.A(new_n668), .B(new_n669), .C1(new_n670), .C2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n663), .B(KEYINPUT85), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n673), .A2(new_n665), .A3(new_n666), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT18), .Z(new_n675));
  NAND3_X1  g250(.A1(new_n671), .A2(new_n673), .A3(new_n670), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n672), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2100), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT87), .B(G2096), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n677), .A2(G2100), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n677), .A2(G2100), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n682), .A2(new_n679), .A3(new_n683), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n681), .A2(new_n684), .ZN(G227));
  XNOR2_X1  g260(.A(G1971), .B(G1976), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1956), .B(G2474), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1961), .B(G1966), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT20), .ZN(new_n693));
  INV_X1    g268(.A(new_n688), .ZN(new_n694));
  INV_X1    g269(.A(new_n691), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n689), .A2(new_n690), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n693), .B(new_n697), .C1(new_n694), .C2(new_n696), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(G1991), .B(G1996), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1981), .B(G1986), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(G229));
  XNOR2_X1  g280(.A(KEYINPUT90), .B(KEYINPUT91), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(new_n592), .B2(new_n597), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT32), .B(G1981), .ZN(new_n710));
  INV_X1    g285(.A(G6), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n711), .A2(G16), .ZN(new_n712));
  NOR3_X1   g287(.A1(new_n709), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n710), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n537), .A2(G48), .ZN(new_n715));
  INV_X1    g290(.A(G86), .ZN(new_n716));
  OAI22_X1  g291(.A1(new_n521), .A2(new_n520), .B1(new_n574), .B2(new_n575), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n715), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n505), .A2(G61), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT80), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n593), .B(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n507), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(G16), .B1(new_n718), .B2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n712), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n714), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n707), .B1(new_n713), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n708), .A2(G22), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G166), .B2(new_n708), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT92), .B(G1971), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT93), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(G303), .A2(G16), .ZN(new_n732));
  INV_X1    g307(.A(new_n730), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n732), .A2(new_n727), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n710), .B1(new_n709), .B2(new_n712), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n723), .A2(new_n714), .A3(new_n724), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n735), .A2(new_n736), .A3(new_n706), .ZN(new_n737));
  NAND4_X1  g312(.A1(new_n726), .A2(new_n731), .A3(new_n734), .A4(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G1976), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n708), .A2(G23), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n587), .B2(G16), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT33), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n739), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n741), .A2(new_n742), .ZN(new_n746));
  AOI211_X1 g321(.A(KEYINPUT33), .B(new_n740), .C1(new_n587), .C2(G16), .ZN(new_n747));
  NOR3_X1   g322(.A1(new_n746), .A2(new_n747), .A3(G1976), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  NOR3_X1   g324(.A1(new_n738), .A2(new_n749), .A3(KEYINPUT34), .ZN(new_n750));
  INV_X1    g325(.A(G29), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G25), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n480), .A2(G131), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n476), .A2(G119), .ZN(new_n754));
  OR2_X1    g329(.A1(G95), .A2(G2105), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n755), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n753), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n752), .B1(new_n758), .B2(new_n751), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT35), .B(G1991), .Z(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  OAI211_X1 g336(.A(G16), .B(new_n603), .C1(new_n604), .C2(new_n605), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT89), .ZN(new_n763));
  NOR2_X1   g338(.A1(G16), .A2(G24), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n762), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n763), .B1(new_n762), .B2(new_n765), .ZN(new_n768));
  NOR3_X1   g343(.A1(new_n767), .A2(new_n768), .A3(G1986), .ZN(new_n769));
  INV_X1    g344(.A(G1986), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n762), .A2(new_n765), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n771), .A2(KEYINPUT89), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n770), .B1(new_n772), .B2(new_n766), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n761), .B1(new_n769), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(KEYINPUT94), .B1(new_n750), .B2(new_n774), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n726), .A2(new_n737), .ZN(new_n776));
  AND2_X1   g351(.A1(new_n731), .A2(new_n734), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT34), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n743), .A2(new_n739), .A3(new_n744), .ZN(new_n779));
  OAI21_X1  g354(.A(G1976), .B1(new_n746), .B2(new_n747), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n776), .A2(new_n777), .A3(new_n778), .A4(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT94), .ZN(new_n783));
  INV_X1    g358(.A(new_n760), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n759), .B(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(G1986), .B1(new_n767), .B2(new_n768), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n772), .A2(new_n766), .A3(new_n770), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n785), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n782), .A2(new_n783), .A3(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(KEYINPUT34), .B1(new_n738), .B2(new_n749), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n790), .A2(KEYINPUT95), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT95), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n792), .B(KEYINPUT34), .C1(new_n738), .C2(new_n749), .ZN(new_n793));
  AOI22_X1  g368(.A1(new_n775), .A2(new_n789), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT36), .ZN(new_n795));
  OAI21_X1  g370(.A(KEYINPUT96), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n791), .A2(new_n793), .ZN(new_n797));
  NOR3_X1   g372(.A1(new_n750), .A2(new_n774), .A3(KEYINPUT94), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n783), .B1(new_n782), .B2(new_n788), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT96), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n800), .A2(new_n801), .A3(KEYINPUT36), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n796), .A2(new_n802), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n797), .B(new_n795), .C1(new_n798), .C2(new_n799), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(KEYINPUT97), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n775), .A2(new_n789), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT97), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n806), .A2(new_n807), .A3(new_n795), .A4(new_n797), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n803), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n708), .A2(G19), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n557), .B2(new_n708), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n812), .A2(G1341), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n476), .A2(G129), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT98), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n468), .A2(G105), .ZN(new_n816));
  NAND3_X1  g391(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT26), .ZN(new_n818));
  AOI211_X1 g393(.A(new_n816), .B(new_n818), .C1(G141), .C2(new_n480), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  MUX2_X1   g395(.A(G32), .B(new_n820), .S(G29), .Z(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT27), .B(G1996), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n813), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(G1961), .ZN(new_n825));
  NOR2_X1   g400(.A1(G5), .A2(G16), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT100), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(G301), .B2(new_n708), .ZN(new_n828));
  OAI221_X1 g403(.A(new_n824), .B1(new_n825), .B2(new_n828), .C1(new_n821), .C2(new_n823), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT31), .B(G11), .ZN(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT99), .B(G28), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n831), .A2(KEYINPUT30), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(KEYINPUT30), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(new_n751), .ZN(new_n834));
  OAI221_X1 g409(.A(new_n830), .B1(new_n832), .B2(new_n834), .C1(new_n633), .C2(new_n751), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT24), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n751), .B1(new_n836), .B2(G34), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(new_n836), .B2(G34), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(G160), .B2(G29), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n835), .B1(G2084), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n812), .A2(G1341), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n480), .A2(G140), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n476), .A2(G128), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n461), .A2(G116), .ZN(new_n844));
  OAI21_X1  g419(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n842), .B(new_n843), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(G29), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n751), .A2(G26), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT28), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(G2067), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n828), .A2(new_n825), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n840), .A2(new_n841), .A3(new_n852), .A4(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n829), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n708), .A2(G21), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n856), .B1(G168), .B2(new_n708), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(G1966), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n708), .A2(G20), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(KEYINPUT23), .Z(new_n860));
  AOI21_X1  g435(.A(new_n860), .B1(G299), .B2(G16), .ZN(new_n861));
  INV_X1    g436(.A(G1956), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n858), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n751), .A2(G35), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n865), .B1(G162), .B2(new_n751), .ZN(new_n866));
  XOR2_X1   g441(.A(KEYINPUT29), .B(G2090), .Z(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n751), .A2(G27), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n869), .B1(G164), .B2(new_n751), .ZN(new_n870));
  INV_X1    g445(.A(G2078), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n870), .B(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(G4), .A2(G16), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n873), .B1(new_n615), .B2(G16), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n657), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n839), .A2(G2084), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n751), .A2(G33), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n480), .A2(G139), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n879), .B(KEYINPUT25), .Z(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  AOI22_X1  g456(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n882), .A2(new_n461), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n877), .B1(new_n884), .B2(new_n751), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(G2072), .Z(new_n886));
  AND4_X1   g461(.A1(new_n872), .A2(new_n875), .A3(new_n876), .A4(new_n886), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n855), .A2(new_n864), .A3(new_n868), .A4(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(KEYINPUT101), .B1(new_n810), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT101), .ZN(new_n891));
  AOI211_X1 g466(.A(new_n891), .B(new_n888), .C1(new_n803), .C2(new_n809), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n890), .A2(new_n892), .ZN(G311));
  NAND2_X1  g468(.A1(new_n810), .A2(new_n889), .ZN(G150));
  AOI22_X1  g469(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n895));
  INV_X1    g470(.A(G93), .ZN(new_n896));
  OAI22_X1  g471(.A1(new_n895), .A2(new_n507), .B1(new_n896), .B2(new_n717), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n897), .B1(G55), .B2(new_n539), .ZN(new_n898));
  INV_X1    g473(.A(G860), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT37), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n614), .A2(new_n622), .ZN(new_n902));
  XNOR2_X1  g477(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n902), .B(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n898), .A2(new_n550), .A3(new_n555), .ZN(new_n905));
  INV_X1    g480(.A(new_n897), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n539), .A2(G55), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(new_n556), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n904), .B(new_n910), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n911), .A2(KEYINPUT39), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n899), .B1(new_n911), .B2(KEYINPUT39), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n901), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  XOR2_X1   g489(.A(new_n914), .B(KEYINPUT103), .Z(G145));
  INV_X1    g490(.A(G37), .ZN(new_n916));
  XNOR2_X1  g491(.A(G162), .B(G160), .ZN(new_n917));
  INV_X1    g492(.A(new_n633), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n918), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n476), .A2(G130), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n461), .A2(G118), .ZN(new_n923));
  OAI21_X1  g498(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n925), .B1(G142), .B2(new_n480), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(new_n636), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(new_n758), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  NOR3_X1   g504(.A1(new_n881), .A2(KEYINPUT104), .A3(new_n883), .ZN(new_n930));
  XOR2_X1   g505(.A(new_n820), .B(new_n930), .Z(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n846), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n931), .A2(new_n846), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n499), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OR2_X1    g510(.A1(new_n931), .A2(new_n846), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n936), .A2(G164), .A3(new_n932), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n929), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n935), .A2(new_n937), .A3(new_n929), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n921), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n940), .ZN(new_n942));
  NOR3_X1   g517(.A1(new_n942), .A2(new_n938), .A3(KEYINPUT105), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n919), .B(new_n920), .C1(new_n940), .C2(new_n944), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n916), .B(new_n941), .C1(new_n943), .C2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n946), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g522(.A1(new_n908), .A2(G868), .ZN(new_n948));
  XNOR2_X1  g523(.A(G290), .B(G166), .ZN(new_n949));
  XNOR2_X1  g524(.A(G305), .B(new_n587), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n949), .B(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT42), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n953), .B(KEYINPUT106), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n624), .B(new_n910), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n615), .A2(new_n619), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT41), .ZN(new_n957));
  AOI22_X1  g532(.A1(new_n611), .A2(new_n613), .B1(new_n571), .B2(new_n578), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n956), .A2(new_n957), .A3(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n614), .A2(G299), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT41), .B1(new_n961), .B2(new_n958), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n955), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n956), .A2(new_n959), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n963), .B1(new_n955), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT108), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT42), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n951), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(KEYINPUT107), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n954), .A2(new_n968), .A3(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n966), .A2(new_n967), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n972), .B(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n948), .B1(new_n974), .B2(G868), .ZN(G295));
  AOI21_X1  g550(.A(new_n948), .B1(new_n974), .B2(G868), .ZN(G331));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n905), .A2(new_n909), .A3(G301), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(G301), .B1(new_n905), .B2(new_n909), .ZN(new_n980));
  NOR3_X1   g555(.A1(new_n979), .A2(new_n980), .A3(G286), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n910), .A2(G171), .ZN(new_n982));
  AOI21_X1  g557(.A(G168), .B1(new_n982), .B2(new_n978), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n965), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(G286), .B1(new_n979), .B2(new_n980), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n960), .A2(new_n962), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n982), .A2(G168), .A3(new_n978), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n984), .A2(new_n952), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(G37), .B1(new_n989), .B2(KEYINPUT109), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT109), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n984), .A2(new_n988), .A3(new_n991), .A4(new_n952), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n964), .A2(KEYINPUT110), .A3(KEYINPUT41), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n985), .A2(new_n993), .A3(new_n987), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n986), .A2(KEYINPUT110), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n964), .B1(new_n985), .B2(new_n987), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n951), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n990), .A2(new_n992), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n977), .B1(new_n999), .B2(KEYINPUT43), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n989), .A2(KEYINPUT109), .ZN(new_n1001));
  INV_X1    g576(.A(new_n988), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n951), .B1(new_n1002), .B2(new_n997), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n1001), .A2(new_n916), .A3(new_n992), .A4(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1000), .B1(KEYINPUT43), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT111), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(KEYINPUT43), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT43), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n990), .A2(new_n1008), .A3(new_n992), .A4(new_n998), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1006), .B1(new_n1010), .B2(new_n977), .ZN(new_n1011));
  AOI211_X1 g586(.A(KEYINPUT111), .B(KEYINPUT44), .C1(new_n1007), .C2(new_n1009), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1005), .B1(new_n1011), .B2(new_n1012), .ZN(G397));
  INV_X1    g588(.A(KEYINPUT45), .ZN(new_n1014));
  AOI21_X1  g589(.A(G1384), .B1(new_n490), .B2(new_n498), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1014), .B1(new_n1015), .B2(KEYINPUT112), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT112), .ZN(new_n1017));
  AOI211_X1 g592(.A(new_n1017), .B(G1384), .C1(new_n490), .C2(new_n498), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G40), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n465), .A2(new_n470), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1023), .A2(G1996), .A3(new_n820), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT113), .ZN(new_n1025));
  OR2_X1    g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n846), .B(new_n851), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1028), .B1(G1996), .B2(new_n820), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1023), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1026), .A2(new_n1027), .A3(new_n1030), .ZN(new_n1031));
  OR2_X1    g606(.A1(G290), .A2(G1986), .ZN(new_n1032));
  NAND2_X1  g607(.A1(G290), .A2(G1986), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1022), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n757), .A2(new_n784), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n758), .A2(new_n760), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1022), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NOR3_X1   g612(.A1(new_n1031), .A2(new_n1034), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G8), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1039), .B1(new_n1021), .B2(new_n1015), .ZN(new_n1040));
  OR2_X1    g615(.A1(new_n587), .A2(new_n739), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT52), .ZN(new_n1043));
  NAND2_X1  g618(.A1(G305), .A2(G1981), .ZN(new_n1044));
  INV_X1    g619(.A(G1981), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n592), .A2(new_n1045), .A3(new_n597), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1044), .B(new_n1046), .C1(KEYINPUT115), .C2(KEYINPUT49), .ZN(new_n1047));
  NOR2_X1   g622(.A1(KEYINPUT115), .A2(KEYINPUT49), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1046), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1045), .B1(new_n592), .B2(new_n597), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1048), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1047), .A2(new_n1051), .A3(new_n1040), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT52), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n589), .A2(new_n739), .A3(new_n590), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1040), .A2(new_n1053), .A3(new_n1041), .A4(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1043), .A2(new_n1052), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT118), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT118), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1043), .A2(new_n1052), .A3(new_n1058), .A4(new_n1055), .ZN(new_n1059));
  NOR2_X1   g634(.A1(G166), .A2(new_n1039), .ZN(new_n1060));
  XNOR2_X1  g635(.A(new_n1060), .B(KEYINPUT55), .ZN(new_n1061));
  INV_X1    g636(.A(G1384), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n499), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n1014), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1015), .A2(KEYINPUT45), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1064), .A2(new_n1021), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G1971), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1063), .A2(KEYINPUT50), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT50), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1015), .A2(new_n1070), .ZN(new_n1071));
  XOR2_X1   g646(.A(KEYINPUT114), .B(G2090), .Z(new_n1072));
  NAND4_X1  g647(.A1(new_n1069), .A2(new_n1071), .A3(new_n1021), .A4(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1039), .B1(new_n1068), .B2(new_n1073), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1057), .A2(new_n1059), .B1(new_n1061), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1021), .B1(new_n1015), .B2(new_n1070), .ZN(new_n1077));
  AOI211_X1 g652(.A(KEYINPUT50), .B(G1384), .C1(new_n490), .C2(new_n498), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1076), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1069), .A2(KEYINPUT116), .A3(new_n1071), .A4(new_n1021), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1079), .A2(new_n1080), .A3(new_n1072), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT117), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1081), .A2(new_n1082), .A3(new_n1068), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1082), .B1(new_n1081), .B2(new_n1068), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n1083), .A2(new_n1084), .A3(new_n1039), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1075), .B1(new_n1085), .B2(new_n1061), .ZN(new_n1086));
  INV_X1    g661(.A(G1966), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1021), .B1(new_n1015), .B2(KEYINPUT45), .ZN(new_n1088));
  AOI211_X1 g663(.A(new_n1014), .B(G1384), .C1(new_n490), .C2(new_n498), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1087), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(G2084), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1069), .A2(new_n1091), .A3(new_n1071), .A4(new_n1021), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1090), .A2(new_n1092), .A3(G168), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(G8), .ZN(new_n1094));
  AOI21_X1  g669(.A(G168), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT51), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT51), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1093), .A2(new_n1097), .A3(G8), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1065), .A2(KEYINPUT53), .A3(new_n871), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1021), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT122), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1100), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  OAI211_X1 g678(.A(KEYINPUT122), .B(new_n1021), .C1(new_n1016), .C2(new_n1018), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1069), .A2(new_n1071), .A3(new_n1021), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1103), .A2(new_n1104), .B1(new_n825), .B2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1064), .A2(new_n871), .A3(new_n1021), .A4(new_n1065), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT53), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(G301), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1110));
  NOR3_X1   g685(.A1(new_n1088), .A2(G2078), .A3(new_n1089), .ZN(new_n1111));
  AOI22_X1  g686(.A1(new_n1111), .A2(KEYINPUT53), .B1(new_n1105), .B2(new_n825), .ZN(new_n1112));
  AOI21_X1  g687(.A(G171), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT54), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1099), .B1(new_n1110), .B2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1086), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(G301), .B1(new_n1112), .B2(new_n1109), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1100), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1119), .A2(new_n1104), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1105), .A2(new_n825), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1121), .A2(new_n1122), .A3(new_n1113), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1118), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1121), .A2(KEYINPUT123), .A3(new_n1122), .A4(new_n1113), .ZN(new_n1126));
  AOI211_X1 g701(.A(KEYINPUT124), .B(KEYINPUT54), .C1(new_n1125), .C2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT124), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1118), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1129), .A2(new_n1126), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT54), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1128), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1117), .B1(new_n1127), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n862), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1136));
  XNOR2_X1  g711(.A(KEYINPUT56), .B(G2072), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1064), .A2(new_n1021), .A3(new_n1065), .A4(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT57), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n571), .A2(new_n1140), .A3(new_n578), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1140), .B1(new_n571), .B2(new_n578), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1139), .A2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1144), .A2(new_n1136), .A3(new_n1138), .A4(KEYINPUT119), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1146), .A2(KEYINPUT61), .A3(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1144), .A2(new_n1136), .A3(new_n1138), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT119), .ZN(new_n1150));
  AND2_X1   g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1135), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1144), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT61), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1155), .A2(KEYINPUT120), .A3(new_n1156), .A4(new_n1147), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1152), .A2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(KEYINPUT61), .B1(new_n1146), .B2(new_n1149), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1066), .A2(G1996), .ZN(new_n1160));
  AND2_X1   g735(.A1(new_n1021), .A2(new_n1015), .ZN(new_n1161));
  XNOR2_X1  g736(.A(KEYINPUT58), .B(G1341), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n557), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(KEYINPUT59), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT59), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1166), .B(new_n557), .C1(new_n1160), .C2(new_n1163), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1159), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1158), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(KEYINPUT121), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT121), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1158), .A2(new_n1171), .A3(new_n1168), .ZN(new_n1172));
  AOI22_X1  g747(.A1(new_n1105), .A2(new_n657), .B1(new_n851), .B2(new_n1161), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(KEYINPUT60), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n1174), .B(new_n615), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1175), .B1(KEYINPUT60), .B2(new_n1173), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1170), .A2(new_n1172), .A3(new_n1176), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1173), .A2(new_n614), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1153), .B1(new_n1178), .B2(new_n1149), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1134), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  AND3_X1   g755(.A1(new_n1096), .A2(KEYINPUT62), .A3(new_n1098), .ZN(new_n1181));
  AOI21_X1  g756(.A(KEYINPUT62), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  OAI211_X1 g758(.A(new_n1118), .B(new_n1075), .C1(new_n1085), .C2(new_n1061), .ZN(new_n1184));
  OAI21_X1  g759(.A(KEYINPUT125), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1081), .A2(new_n1068), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1039), .B1(new_n1186), .B2(KEYINPUT117), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1081), .A2(new_n1082), .A3(new_n1068), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1061), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1074), .A2(new_n1061), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NOR3_X1   g767(.A1(new_n1189), .A2(new_n1192), .A3(new_n1130), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT62), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1099), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1096), .A2(KEYINPUT62), .A3(new_n1098), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT125), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1193), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1185), .A2(new_n1199), .ZN(new_n1200));
  AOI211_X1 g775(.A(G1976), .B(G288), .C1(new_n1047), .C2(new_n1051), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1040), .B1(new_n1201), .B2(new_n1049), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1202), .B1(new_n1191), .B2(new_n1056), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT63), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1205), .A2(G8), .A3(G168), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1204), .B1(new_n1086), .B2(new_n1206), .ZN(new_n1207));
  NOR3_X1   g782(.A1(new_n1206), .A2(new_n1056), .A3(new_n1204), .ZN(new_n1208));
  OR2_X1    g783(.A1(new_n1074), .A2(new_n1061), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1208), .A2(new_n1209), .A3(new_n1191), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1203), .B1(new_n1207), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1200), .A2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1038), .B1(new_n1180), .B2(new_n1212), .ZN(new_n1213));
  NOR2_X1   g788(.A1(new_n1031), .A2(new_n1037), .ZN(new_n1214));
  OR2_X1    g789(.A1(new_n1214), .A2(KEYINPUT126), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1214), .A2(KEYINPUT126), .ZN(new_n1216));
  NOR2_X1   g791(.A1(new_n1022), .A2(new_n1032), .ZN(new_n1217));
  XOR2_X1   g792(.A(new_n1217), .B(KEYINPUT48), .Z(new_n1218));
  NAND3_X1  g793(.A1(new_n1215), .A2(new_n1216), .A3(new_n1218), .ZN(new_n1219));
  INV_X1    g794(.A(new_n1028), .ZN(new_n1220));
  OAI21_X1  g795(.A(new_n1023), .B1(new_n820), .B2(new_n1220), .ZN(new_n1221));
  INV_X1    g796(.A(KEYINPUT46), .ZN(new_n1222));
  INV_X1    g797(.A(G1996), .ZN(new_n1223));
  AOI21_X1  g798(.A(new_n1222), .B1(new_n1023), .B2(new_n1223), .ZN(new_n1224));
  NOR3_X1   g799(.A1(new_n1022), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1225));
  OAI21_X1  g800(.A(new_n1221), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  XNOR2_X1  g801(.A(new_n1226), .B(KEYINPUT47), .ZN(new_n1227));
  OAI22_X1  g802(.A1(new_n1031), .A2(new_n1036), .B1(G2067), .B2(new_n846), .ZN(new_n1228));
  NAND2_X1  g803(.A1(new_n1228), .A2(new_n1023), .ZN(new_n1229));
  AND3_X1   g804(.A1(new_n1219), .A2(new_n1227), .A3(new_n1229), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1213), .A2(new_n1230), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g806(.A(new_n459), .B1(new_n681), .B2(new_n684), .ZN(new_n1233));
  OAI21_X1  g807(.A(new_n1233), .B1(new_n660), .B2(new_n661), .ZN(new_n1234));
  XNOR2_X1  g808(.A(new_n1234), .B(KEYINPUT127), .ZN(new_n1235));
  NAND4_X1  g809(.A1(new_n1235), .A2(new_n704), .A3(new_n946), .A4(new_n1010), .ZN(G225));
  INV_X1    g810(.A(G225), .ZN(G308));
endmodule


