

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U554 ( .A(G2104), .ZN(n624) );
  OR2_X1 U555 ( .A1(n764), .A2(n763), .ZN(n777) );
  AND2_X1 U556 ( .A1(n530), .A2(n527), .ZN(n526) );
  XNOR2_X1 U557 ( .A(n703), .B(n702), .ZN(n531) );
  NOR2_X1 U558 ( .A1(n989), .A2(n657), .ZN(n673) );
  BUF_X1 U559 ( .A(n652), .Z(n696) );
  XNOR2_X1 U560 ( .A(KEYINPUT97), .B(n652), .ZN(n677) );
  NAND2_X1 U561 ( .A1(n635), .A2(n731), .ZN(n652) );
  NOR2_X1 U562 ( .A1(G164), .A2(G1384), .ZN(n731) );
  XNOR2_X1 U563 ( .A(n634), .B(KEYINPUT90), .ZN(G164) );
  NAND2_X2 U564 ( .A1(n535), .A2(n532), .ZN(n918) );
  NOR2_X2 U565 ( .A1(G2105), .A2(n624), .ZN(n917) );
  NOR2_X1 U566 ( .A1(G2104), .A2(KEYINPUT17), .ZN(n537) );
  BUF_X1 U567 ( .A(n627), .Z(n520) );
  XNOR2_X1 U568 ( .A(n619), .B(KEYINPUT65), .ZN(n627) );
  NOR2_X1 U569 ( .A1(n539), .A2(n521), .ZN(n636) );
  INV_X1 U570 ( .A(KEYINPUT32), .ZN(n529) );
  AND2_X1 U571 ( .A1(n1005), .A2(n549), .ZN(n711) );
  NOR2_X1 U572 ( .A1(n641), .A2(n640), .ZN(n642) );
  AND2_X1 U573 ( .A1(n709), .A2(n528), .ZN(n527) );
  NAND2_X1 U574 ( .A1(n529), .A2(n540), .ZN(n528) );
  INV_X1 U575 ( .A(n727), .ZN(n714) );
  INV_X1 U576 ( .A(n993), .ZN(n719) );
  AND2_X1 U577 ( .A1(n534), .A2(n533), .ZN(n532) );
  NAND2_X1 U578 ( .A1(n537), .A2(n536), .ZN(n535) );
  NAND2_X1 U579 ( .A1(G2104), .A2(KEYINPUT17), .ZN(n534) );
  XNOR2_X1 U580 ( .A(KEYINPUT64), .B(n558), .ZN(n818) );
  NOR2_X1 U581 ( .A1(n563), .A2(G543), .ZN(n555) );
  NOR2_X1 U582 ( .A1(n652), .A2(n970), .ZN(n654) );
  NOR2_X1 U583 ( .A1(n696), .A2(G2084), .ZN(n538) );
  XNOR2_X1 U584 ( .A(n642), .B(n546), .ZN(n545) );
  XNOR2_X1 U585 ( .A(KEYINPUT31), .B(KEYINPUT103), .ZN(n546) );
  NAND2_X1 U586 ( .A1(n526), .A2(n524), .ZN(n725) );
  NAND2_X1 U587 ( .A1(n525), .A2(n529), .ZN(n524) );
  INV_X1 U588 ( .A(G2105), .ZN(n536) );
  NAND2_X1 U589 ( .A1(G2105), .A2(KEYINPUT17), .ZN(n533) );
  XNOR2_X1 U590 ( .A(n541), .B(KEYINPUT109), .ZN(n764) );
  NAND2_X1 U591 ( .A1(n544), .A2(n553), .ZN(n543) );
  OR2_X1 U592 ( .A1(n762), .A2(n552), .ZN(n763) );
  NOR2_X1 U593 ( .A1(n550), .A2(n623), .ZN(n780) );
  XNOR2_X1 U594 ( .A(KEYINPUT70), .B(n581), .ZN(G171) );
  XNOR2_X1 U595 ( .A(n572), .B(n571), .ZN(G168) );
  XNOR2_X2 U596 ( .A(KEYINPUT68), .B(n556), .ZN(n658) );
  NAND2_X1 U597 ( .A1(n547), .A2(n545), .ZN(n707) );
  XOR2_X1 U598 ( .A(n538), .B(KEYINPUT95), .Z(n521) );
  OR2_X1 U599 ( .A1(n727), .A2(n722), .ZN(n522) );
  AND2_X1 U600 ( .A1(KEYINPUT32), .A2(G8), .ZN(n523) );
  INV_X1 U601 ( .A(n531), .ZN(n525) );
  NAND2_X1 U602 ( .A1(n531), .A2(n523), .ZN(n530) );
  OR2_X1 U603 ( .A1(n706), .A2(n540), .ZN(n539) );
  INV_X1 U604 ( .A(G8), .ZN(n540) );
  NAND2_X1 U605 ( .A1(n543), .A2(n542), .ZN(n541) );
  AND2_X1 U606 ( .A1(n729), .A2(n522), .ZN(n542) );
  NAND2_X1 U607 ( .A1(n717), .A2(n716), .ZN(n544) );
  NAND2_X1 U608 ( .A1(n707), .A2(G286), .ZN(n701) );
  XNOR2_X1 U609 ( .A(n548), .B(KEYINPUT102), .ZN(n547) );
  NAND2_X1 U610 ( .A1(n694), .A2(n693), .ZN(n548) );
  NAND2_X1 U611 ( .A1(n715), .A2(n714), .ZN(n717) );
  OR2_X1 U612 ( .A1(G1971), .A2(G303), .ZN(n549) );
  AND2_X1 U613 ( .A1(n520), .A2(G125), .ZN(n550) );
  XNOR2_X1 U614 ( .A(n568), .B(KEYINPUT5), .ZN(n551) );
  AND2_X1 U615 ( .A1(n1000), .A2(n774), .ZN(n552) );
  AND2_X1 U616 ( .A1(n720), .A2(n719), .ZN(n553) );
  INV_X1 U617 ( .A(KEYINPUT26), .ZN(n653) );
  INV_X1 U618 ( .A(KEYINPUT98), .ZN(n679) );
  INV_X1 U619 ( .A(KEYINPUT101), .ZN(n671) );
  INV_X1 U620 ( .A(KEYINPUT29), .ZN(n690) );
  XNOR2_X1 U621 ( .A(n691), .B(n690), .ZN(n694) );
  INV_X1 U622 ( .A(KEYINPUT105), .ZN(n702) );
  INV_X1 U623 ( .A(KEYINPUT1), .ZN(n554) );
  INV_X1 U624 ( .A(KEYINPUT0), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n555), .B(n554), .ZN(n556) );
  INV_X1 U626 ( .A(KEYINPUT6), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n557), .B(G543), .ZN(n598) );
  AND2_X1 U628 ( .A1(G2104), .A2(G2105), .ZN(n912) );
  XNOR2_X1 U629 ( .A(n570), .B(KEYINPUT75), .ZN(n572) );
  XNOR2_X1 U630 ( .A(G651), .B(KEYINPUT67), .ZN(n563) );
  NAND2_X1 U631 ( .A1(G63), .A2(n658), .ZN(n560) );
  NOR2_X1 U632 ( .A1(G651), .A2(n598), .ZN(n558) );
  NAND2_X1 U633 ( .A1(G51), .A2(n818), .ZN(n559) );
  NAND2_X1 U634 ( .A1(n560), .A2(n559), .ZN(n562) );
  XNOR2_X1 U635 ( .A(n562), .B(n561), .ZN(n569) );
  NOR2_X1 U636 ( .A1(n598), .A2(n563), .ZN(n817) );
  NAND2_X1 U637 ( .A1(n817), .A2(G76), .ZN(n564) );
  XNOR2_X1 U638 ( .A(n564), .B(KEYINPUT74), .ZN(n567) );
  NOR2_X1 U639 ( .A1(G651), .A2(G543), .ZN(n814) );
  NAND2_X1 U640 ( .A1(n814), .A2(G89), .ZN(n565) );
  XNOR2_X1 U641 ( .A(KEYINPUT4), .B(n565), .ZN(n566) );
  NAND2_X1 U642 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U643 ( .A1(n569), .A2(n551), .ZN(n570) );
  XOR2_X1 U644 ( .A(KEYINPUT76), .B(KEYINPUT7), .Z(n571) );
  XOR2_X1 U645 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U646 ( .A1(G64), .A2(n658), .ZN(n574) );
  NAND2_X1 U647 ( .A1(G52), .A2(n818), .ZN(n573) );
  NAND2_X1 U648 ( .A1(n574), .A2(n573), .ZN(n580) );
  NAND2_X1 U649 ( .A1(n817), .A2(G77), .ZN(n575) );
  XOR2_X1 U650 ( .A(KEYINPUT69), .B(n575), .Z(n577) );
  NAND2_X1 U651 ( .A1(n814), .A2(G90), .ZN(n576) );
  NAND2_X1 U652 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U653 ( .A(KEYINPUT9), .B(n578), .Z(n579) );
  NOR2_X1 U654 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U655 ( .A1(G78), .A2(n817), .ZN(n583) );
  NAND2_X1 U656 ( .A1(G53), .A2(n818), .ZN(n582) );
  NAND2_X1 U657 ( .A1(n583), .A2(n582), .ZN(n587) );
  NAND2_X1 U658 ( .A1(n814), .A2(G91), .ZN(n585) );
  NAND2_X1 U659 ( .A1(G65), .A2(n658), .ZN(n584) );
  NAND2_X1 U660 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U661 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U662 ( .A(n588), .B(KEYINPUT71), .ZN(G299) );
  NAND2_X1 U663 ( .A1(G88), .A2(n814), .ZN(n590) );
  NAND2_X1 U664 ( .A1(G75), .A2(n817), .ZN(n589) );
  NAND2_X1 U665 ( .A1(n590), .A2(n589), .ZN(n594) );
  NAND2_X1 U666 ( .A1(G62), .A2(n658), .ZN(n592) );
  NAND2_X1 U667 ( .A1(G50), .A2(n818), .ZN(n591) );
  NAND2_X1 U668 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U669 ( .A1(n594), .A2(n593), .ZN(G166) );
  INV_X1 U670 ( .A(G166), .ZN(G303) );
  NAND2_X1 U671 ( .A1(G651), .A2(G74), .ZN(n596) );
  NAND2_X1 U672 ( .A1(G49), .A2(n818), .ZN(n595) );
  NAND2_X1 U673 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U674 ( .A(n597), .B(KEYINPUT81), .ZN(n600) );
  NAND2_X1 U675 ( .A1(G87), .A2(n598), .ZN(n599) );
  NAND2_X1 U676 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U677 ( .A1(n658), .A2(n601), .ZN(n602) );
  XOR2_X1 U678 ( .A(KEYINPUT82), .B(n602), .Z(G288) );
  NAND2_X1 U679 ( .A1(n814), .A2(G86), .ZN(n604) );
  NAND2_X1 U680 ( .A1(G61), .A2(n658), .ZN(n603) );
  NAND2_X1 U681 ( .A1(n604), .A2(n603), .ZN(n609) );
  XOR2_X1 U682 ( .A(KEYINPUT84), .B(KEYINPUT2), .Z(n606) );
  NAND2_X1 U683 ( .A1(G73), .A2(n817), .ZN(n605) );
  XNOR2_X1 U684 ( .A(n606), .B(n605), .ZN(n607) );
  XOR2_X1 U685 ( .A(KEYINPUT83), .B(n607), .Z(n608) );
  NOR2_X1 U686 ( .A1(n609), .A2(n608), .ZN(n610) );
  XOR2_X1 U687 ( .A(KEYINPUT85), .B(n610), .Z(n612) );
  NAND2_X1 U688 ( .A1(G48), .A2(n818), .ZN(n611) );
  NAND2_X1 U689 ( .A1(n612), .A2(n611), .ZN(G305) );
  AND2_X1 U690 ( .A1(n814), .A2(G85), .ZN(n616) );
  NAND2_X1 U691 ( .A1(G60), .A2(n658), .ZN(n614) );
  NAND2_X1 U692 ( .A1(G47), .A2(n818), .ZN(n613) );
  NAND2_X1 U693 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U694 ( .A1(n616), .A2(n615), .ZN(n618) );
  NAND2_X1 U695 ( .A1(n817), .A2(G72), .ZN(n617) );
  NAND2_X1 U696 ( .A1(n618), .A2(n617), .ZN(G290) );
  NAND2_X1 U697 ( .A1(n624), .A2(G2105), .ZN(n619) );
  NAND2_X1 U698 ( .A1(G113), .A2(n912), .ZN(n621) );
  NAND2_X1 U699 ( .A1(G137), .A2(n918), .ZN(n620) );
  NAND2_X1 U700 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U701 ( .A(n622), .B(KEYINPUT66), .ZN(n623) );
  NAND2_X1 U702 ( .A1(G101), .A2(n917), .ZN(n625) );
  XOR2_X1 U703 ( .A(KEYINPUT23), .B(n625), .Z(n779) );
  AND2_X1 U704 ( .A1(n779), .A2(G40), .ZN(n626) );
  NAND2_X1 U705 ( .A1(n780), .A2(n626), .ZN(n730) );
  INV_X1 U706 ( .A(n730), .ZN(n635) );
  NAND2_X1 U707 ( .A1(G126), .A2(n627), .ZN(n629) );
  NAND2_X1 U708 ( .A1(G138), .A2(n918), .ZN(n628) );
  NAND2_X1 U709 ( .A1(n629), .A2(n628), .ZN(n633) );
  NAND2_X1 U710 ( .A1(G114), .A2(n912), .ZN(n631) );
  NAND2_X1 U711 ( .A1(G102), .A2(n917), .ZN(n630) );
  NAND2_X1 U712 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U713 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U714 ( .A1(G8), .A2(n652), .ZN(n727) );
  NOR2_X1 U715 ( .A1(G1966), .A2(n727), .ZN(n706) );
  XOR2_X1 U716 ( .A(KEYINPUT30), .B(n636), .Z(n637) );
  NOR2_X1 U717 ( .A1(G168), .A2(n637), .ZN(n641) );
  INV_X1 U718 ( .A(G1961), .ZN(n1021) );
  NAND2_X1 U719 ( .A1(n1021), .A2(n696), .ZN(n639) );
  XNOR2_X1 U720 ( .A(G2078), .B(KEYINPUT25), .ZN(n969) );
  NAND2_X1 U721 ( .A1(n677), .A2(n969), .ZN(n638) );
  NAND2_X1 U722 ( .A1(n639), .A2(n638), .ZN(n692) );
  NOR2_X1 U723 ( .A1(G171), .A2(n692), .ZN(n640) );
  NAND2_X1 U724 ( .A1(n658), .A2(G56), .ZN(n643) );
  XOR2_X1 U725 ( .A(KEYINPUT14), .B(n643), .Z(n649) );
  NAND2_X1 U726 ( .A1(n814), .A2(G81), .ZN(n644) );
  XNOR2_X1 U727 ( .A(n644), .B(KEYINPUT12), .ZN(n646) );
  NAND2_X1 U728 ( .A1(G68), .A2(n817), .ZN(n645) );
  NAND2_X1 U729 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U730 ( .A(KEYINPUT13), .B(n647), .Z(n648) );
  NOR2_X1 U731 ( .A1(n649), .A2(n648), .ZN(n651) );
  NAND2_X1 U732 ( .A1(G43), .A2(n818), .ZN(n650) );
  NAND2_X1 U733 ( .A1(n651), .A2(n650), .ZN(n989) );
  INV_X1 U734 ( .A(G1996), .ZN(n970) );
  XNOR2_X1 U735 ( .A(n654), .B(n653), .ZN(n656) );
  NAND2_X1 U736 ( .A1(n696), .A2(G1341), .ZN(n655) );
  NAND2_X1 U737 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U738 ( .A1(n814), .A2(G92), .ZN(n660) );
  NAND2_X1 U739 ( .A1(G66), .A2(n658), .ZN(n659) );
  NAND2_X1 U740 ( .A1(n660), .A2(n659), .ZN(n664) );
  NAND2_X1 U741 ( .A1(G79), .A2(n817), .ZN(n662) );
  NAND2_X1 U742 ( .A1(G54), .A2(n818), .ZN(n661) );
  NAND2_X1 U743 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U744 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X2 U745 ( .A(KEYINPUT15), .B(n665), .Z(n988) );
  NAND2_X1 U746 ( .A1(n673), .A2(n988), .ZN(n670) );
  NAND2_X1 U747 ( .A1(G1348), .A2(n696), .ZN(n666) );
  XNOR2_X1 U748 ( .A(n666), .B(KEYINPUT100), .ZN(n668) );
  NAND2_X1 U749 ( .A1(n677), .A2(G2067), .ZN(n667) );
  NAND2_X1 U750 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U751 ( .A1(n670), .A2(n669), .ZN(n672) );
  XNOR2_X1 U752 ( .A(n672), .B(n671), .ZN(n675) );
  OR2_X1 U753 ( .A1(n988), .A2(n673), .ZN(n674) );
  NAND2_X1 U754 ( .A1(n675), .A2(n674), .ZN(n684) );
  NAND2_X1 U755 ( .A1(n677), .A2(G2072), .ZN(n676) );
  XNOR2_X1 U756 ( .A(KEYINPUT27), .B(n676), .ZN(n682) );
  INV_X1 U757 ( .A(n677), .ZN(n678) );
  NAND2_X1 U758 ( .A1(G1956), .A2(n678), .ZN(n680) );
  XNOR2_X1 U759 ( .A(n680), .B(n679), .ZN(n681) );
  NOR2_X1 U760 ( .A1(n682), .A2(n681), .ZN(n685) );
  INV_X1 U761 ( .A(G299), .ZN(n827) );
  NAND2_X1 U762 ( .A1(n685), .A2(n827), .ZN(n683) );
  NAND2_X1 U763 ( .A1(n684), .A2(n683), .ZN(n689) );
  NOR2_X1 U764 ( .A1(n685), .A2(n827), .ZN(n687) );
  XNOR2_X1 U765 ( .A(KEYINPUT99), .B(KEYINPUT28), .ZN(n686) );
  XNOR2_X1 U766 ( .A(n687), .B(n686), .ZN(n688) );
  NAND2_X1 U767 ( .A1(n689), .A2(n688), .ZN(n691) );
  NAND2_X1 U768 ( .A1(G171), .A2(n692), .ZN(n693) );
  NOR2_X1 U769 ( .A1(G1971), .A2(n727), .ZN(n695) );
  XNOR2_X1 U770 ( .A(n695), .B(KEYINPUT104), .ZN(n698) );
  NOR2_X1 U771 ( .A1(n696), .A2(G2090), .ZN(n697) );
  NOR2_X1 U772 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U773 ( .A1(n699), .A2(G303), .ZN(n700) );
  NAND2_X1 U774 ( .A1(n701), .A2(n700), .ZN(n703) );
  NAND2_X1 U775 ( .A1(G8), .A2(n521), .ZN(n704) );
  XOR2_X1 U776 ( .A(KEYINPUT96), .B(n704), .Z(n705) );
  NOR2_X1 U777 ( .A1(n706), .A2(n705), .ZN(n708) );
  NAND2_X1 U778 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U779 ( .A1(G1976), .A2(G288), .ZN(n710) );
  XOR2_X1 U780 ( .A(KEYINPUT106), .B(n710), .Z(n1005) );
  NAND2_X1 U781 ( .A1(n725), .A2(n711), .ZN(n712) );
  NAND2_X1 U782 ( .A1(G1976), .A2(G288), .ZN(n1001) );
  NAND2_X1 U783 ( .A1(n712), .A2(n1001), .ZN(n713) );
  XNOR2_X1 U784 ( .A(n713), .B(KEYINPUT107), .ZN(n715) );
  INV_X1 U785 ( .A(KEYINPUT33), .ZN(n716) );
  NOR2_X1 U786 ( .A1(n727), .A2(n1005), .ZN(n718) );
  NAND2_X1 U787 ( .A1(KEYINPUT33), .A2(n718), .ZN(n720) );
  XNOR2_X1 U788 ( .A(G1981), .B(G305), .ZN(n993) );
  NOR2_X1 U789 ( .A1(G1981), .A2(G305), .ZN(n721) );
  XOR2_X1 U790 ( .A(n721), .B(KEYINPUT24), .Z(n722) );
  NOR2_X1 U791 ( .A1(G2090), .A2(G303), .ZN(n723) );
  NAND2_X1 U792 ( .A1(G8), .A2(n723), .ZN(n724) );
  NAND2_X1 U793 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U794 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U795 ( .A(KEYINPUT108), .B(n728), .ZN(n729) );
  NOR2_X1 U796 ( .A1(n731), .A2(n730), .ZN(n774) );
  XNOR2_X1 U797 ( .A(KEYINPUT37), .B(G2067), .ZN(n772) );
  NAND2_X1 U798 ( .A1(n912), .A2(G116), .ZN(n732) );
  XNOR2_X1 U799 ( .A(n732), .B(KEYINPUT92), .ZN(n734) );
  NAND2_X1 U800 ( .A1(G128), .A2(n520), .ZN(n733) );
  NAND2_X1 U801 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U802 ( .A(n735), .B(KEYINPUT35), .ZN(n741) );
  XNOR2_X1 U803 ( .A(KEYINPUT34), .B(KEYINPUT91), .ZN(n739) );
  NAND2_X1 U804 ( .A1(G104), .A2(n917), .ZN(n737) );
  NAND2_X1 U805 ( .A1(G140), .A2(n918), .ZN(n736) );
  NAND2_X1 U806 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U807 ( .A(n739), .B(n738), .ZN(n740) );
  NAND2_X1 U808 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U809 ( .A(KEYINPUT36), .B(n742), .Z(n906) );
  OR2_X1 U810 ( .A1(n772), .A2(n906), .ZN(n743) );
  XNOR2_X1 U811 ( .A(KEYINPUT93), .B(n743), .ZN(n947) );
  NAND2_X1 U812 ( .A1(n774), .A2(n947), .ZN(n770) );
  NAND2_X1 U813 ( .A1(G95), .A2(n917), .ZN(n745) );
  NAND2_X1 U814 ( .A1(G131), .A2(n918), .ZN(n744) );
  NAND2_X1 U815 ( .A1(n745), .A2(n744), .ZN(n749) );
  NAND2_X1 U816 ( .A1(G107), .A2(n912), .ZN(n747) );
  NAND2_X1 U817 ( .A1(G119), .A2(n520), .ZN(n746) );
  NAND2_X1 U818 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U819 ( .A1(n749), .A2(n748), .ZN(n904) );
  INV_X1 U820 ( .A(G1991), .ZN(n967) );
  NOR2_X1 U821 ( .A1(n904), .A2(n967), .ZN(n759) );
  NAND2_X1 U822 ( .A1(G117), .A2(n912), .ZN(n751) );
  NAND2_X1 U823 ( .A1(G129), .A2(n520), .ZN(n750) );
  NAND2_X1 U824 ( .A1(n751), .A2(n750), .ZN(n754) );
  NAND2_X1 U825 ( .A1(n917), .A2(G105), .ZN(n752) );
  XOR2_X1 U826 ( .A(KEYINPUT38), .B(n752), .Z(n753) );
  NOR2_X1 U827 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U828 ( .A(n755), .B(KEYINPUT94), .ZN(n757) );
  NAND2_X1 U829 ( .A1(G141), .A2(n918), .ZN(n756) );
  NAND2_X1 U830 ( .A1(n757), .A2(n756), .ZN(n900) );
  AND2_X1 U831 ( .A1(G1996), .A2(n900), .ZN(n758) );
  NOR2_X1 U832 ( .A1(n759), .A2(n758), .ZN(n945) );
  INV_X1 U833 ( .A(n774), .ZN(n760) );
  NOR2_X1 U834 ( .A1(n945), .A2(n760), .ZN(n767) );
  INV_X1 U835 ( .A(n767), .ZN(n761) );
  NAND2_X1 U836 ( .A1(n770), .A2(n761), .ZN(n762) );
  XNOR2_X1 U837 ( .A(G1986), .B(G290), .ZN(n1000) );
  NOR2_X1 U838 ( .A1(G1996), .A2(n900), .ZN(n955) );
  AND2_X1 U839 ( .A1(n967), .A2(n904), .ZN(n940) );
  NOR2_X1 U840 ( .A1(G1986), .A2(G290), .ZN(n765) );
  NOR2_X1 U841 ( .A1(n940), .A2(n765), .ZN(n766) );
  NOR2_X1 U842 ( .A1(n767), .A2(n766), .ZN(n768) );
  NOR2_X1 U843 ( .A1(n955), .A2(n768), .ZN(n769) );
  XNOR2_X1 U844 ( .A(n769), .B(KEYINPUT39), .ZN(n771) );
  NAND2_X1 U845 ( .A1(n771), .A2(n770), .ZN(n773) );
  NAND2_X1 U846 ( .A1(n772), .A2(n906), .ZN(n944) );
  NAND2_X1 U847 ( .A1(n773), .A2(n944), .ZN(n775) );
  NAND2_X1 U848 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U849 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U850 ( .A(n778), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U851 ( .A1(n780), .A2(n779), .ZN(G160) );
  XOR2_X1 U852 ( .A(G2443), .B(G2446), .Z(n782) );
  XNOR2_X1 U853 ( .A(G2427), .B(G2451), .ZN(n781) );
  XNOR2_X1 U854 ( .A(n782), .B(n781), .ZN(n788) );
  XOR2_X1 U855 ( .A(G2430), .B(G2454), .Z(n784) );
  XNOR2_X1 U856 ( .A(G1348), .B(G1341), .ZN(n783) );
  XNOR2_X1 U857 ( .A(n784), .B(n783), .ZN(n786) );
  XOR2_X1 U858 ( .A(G2435), .B(G2438), .Z(n785) );
  XNOR2_X1 U859 ( .A(n786), .B(n785), .ZN(n787) );
  XOR2_X1 U860 ( .A(n788), .B(n787), .Z(n789) );
  AND2_X1 U861 ( .A1(G14), .A2(n789), .ZN(G401) );
  INV_X1 U862 ( .A(G57), .ZN(G237) );
  AND2_X1 U863 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U864 ( .A(G108), .ZN(G238) );
  INV_X1 U865 ( .A(G120), .ZN(G236) );
  INV_X1 U866 ( .A(G82), .ZN(G220) );
  NAND2_X1 U867 ( .A1(G7), .A2(G661), .ZN(n791) );
  XNOR2_X1 U868 ( .A(n791), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U869 ( .A(G567), .ZN(n848) );
  NOR2_X1 U870 ( .A1(n848), .A2(G223), .ZN(n792) );
  XNOR2_X1 U871 ( .A(n792), .B(KEYINPUT11), .ZN(G234) );
  INV_X1 U872 ( .A(G860), .ZN(n862) );
  OR2_X1 U873 ( .A1(n989), .A2(n862), .ZN(G153) );
  XNOR2_X1 U874 ( .A(KEYINPUT73), .B(G171), .ZN(G301) );
  NAND2_X1 U875 ( .A1(G868), .A2(G301), .ZN(n794) );
  OR2_X1 U876 ( .A1(n988), .A2(G868), .ZN(n793) );
  NAND2_X1 U877 ( .A1(n794), .A2(n793), .ZN(G284) );
  XNOR2_X1 U878 ( .A(KEYINPUT77), .B(G868), .ZN(n795) );
  NOR2_X1 U879 ( .A1(G286), .A2(n795), .ZN(n797) );
  NOR2_X1 U880 ( .A1(G868), .A2(G299), .ZN(n796) );
  NOR2_X1 U881 ( .A1(n797), .A2(n796), .ZN(G297) );
  NAND2_X1 U882 ( .A1(n862), .A2(G559), .ZN(n798) );
  NAND2_X1 U883 ( .A1(n798), .A2(n988), .ZN(n799) );
  XNOR2_X1 U884 ( .A(n799), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U885 ( .A1(G868), .A2(n989), .ZN(n802) );
  NAND2_X1 U886 ( .A1(G868), .A2(n988), .ZN(n800) );
  NOR2_X1 U887 ( .A1(G559), .A2(n800), .ZN(n801) );
  NOR2_X1 U888 ( .A1(n802), .A2(n801), .ZN(G282) );
  NAND2_X1 U889 ( .A1(G111), .A2(n912), .ZN(n804) );
  NAND2_X1 U890 ( .A1(G99), .A2(n917), .ZN(n803) );
  NAND2_X1 U891 ( .A1(n804), .A2(n803), .ZN(n811) );
  NAND2_X1 U892 ( .A1(G123), .A2(n520), .ZN(n805) );
  XNOR2_X1 U893 ( .A(n805), .B(KEYINPUT78), .ZN(n806) );
  XNOR2_X1 U894 ( .A(n806), .B(KEYINPUT18), .ZN(n808) );
  NAND2_X1 U895 ( .A1(G135), .A2(n918), .ZN(n807) );
  NAND2_X1 U896 ( .A1(n808), .A2(n807), .ZN(n809) );
  XOR2_X1 U897 ( .A(KEYINPUT79), .B(n809), .Z(n810) );
  NOR2_X1 U898 ( .A1(n811), .A2(n810), .ZN(n939) );
  XNOR2_X1 U899 ( .A(n939), .B(G2096), .ZN(n813) );
  INV_X1 U900 ( .A(G2100), .ZN(n812) );
  NAND2_X1 U901 ( .A1(n813), .A2(n812), .ZN(G156) );
  XOR2_X1 U902 ( .A(KEYINPUT86), .B(KEYINPUT19), .Z(n825) );
  NAND2_X1 U903 ( .A1(n814), .A2(G93), .ZN(n816) );
  NAND2_X1 U904 ( .A1(G67), .A2(n658), .ZN(n815) );
  NAND2_X1 U905 ( .A1(n816), .A2(n815), .ZN(n822) );
  NAND2_X1 U906 ( .A1(G80), .A2(n817), .ZN(n820) );
  NAND2_X1 U907 ( .A1(G55), .A2(n818), .ZN(n819) );
  NAND2_X1 U908 ( .A1(n820), .A2(n819), .ZN(n821) );
  NOR2_X1 U909 ( .A1(n822), .A2(n821), .ZN(n823) );
  XOR2_X1 U910 ( .A(KEYINPUT80), .B(n823), .Z(n863) );
  XNOR2_X1 U911 ( .A(G166), .B(n863), .ZN(n824) );
  XNOR2_X1 U912 ( .A(n825), .B(n824), .ZN(n826) );
  XNOR2_X1 U913 ( .A(n827), .B(n826), .ZN(n829) );
  XNOR2_X1 U914 ( .A(G290), .B(G288), .ZN(n828) );
  XNOR2_X1 U915 ( .A(n829), .B(n828), .ZN(n830) );
  XOR2_X1 U916 ( .A(n830), .B(G305), .Z(n928) );
  NAND2_X1 U917 ( .A1(G559), .A2(n988), .ZN(n831) );
  XOR2_X1 U918 ( .A(n989), .B(n831), .Z(n861) );
  XNOR2_X1 U919 ( .A(n928), .B(n861), .ZN(n832) );
  NAND2_X1 U920 ( .A1(n832), .A2(G868), .ZN(n835) );
  INV_X1 U921 ( .A(G868), .ZN(n833) );
  NAND2_X1 U922 ( .A1(n833), .A2(n863), .ZN(n834) );
  NAND2_X1 U923 ( .A1(n835), .A2(n834), .ZN(G295) );
  NAND2_X1 U924 ( .A1(G2084), .A2(G2078), .ZN(n836) );
  XOR2_X1 U925 ( .A(KEYINPUT20), .B(n836), .Z(n837) );
  NAND2_X1 U926 ( .A1(G2090), .A2(n837), .ZN(n838) );
  XNOR2_X1 U927 ( .A(KEYINPUT21), .B(n838), .ZN(n839) );
  NAND2_X1 U928 ( .A1(n839), .A2(G2072), .ZN(G158) );
  XOR2_X1 U929 ( .A(KEYINPUT72), .B(G132), .Z(G219) );
  XNOR2_X1 U930 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U931 ( .A1(G219), .A2(G220), .ZN(n841) );
  XNOR2_X1 U932 ( .A(KEYINPUT87), .B(KEYINPUT22), .ZN(n840) );
  XNOR2_X1 U933 ( .A(n841), .B(n840), .ZN(n842) );
  NOR2_X1 U934 ( .A1(n842), .A2(G218), .ZN(n843) );
  NAND2_X1 U935 ( .A1(G96), .A2(n843), .ZN(n844) );
  XNOR2_X1 U936 ( .A(KEYINPUT88), .B(n844), .ZN(n860) );
  NAND2_X1 U937 ( .A1(n860), .A2(G2106), .ZN(n845) );
  XNOR2_X1 U938 ( .A(n845), .B(KEYINPUT89), .ZN(n850) );
  NOR2_X1 U939 ( .A1(G236), .A2(G238), .ZN(n846) );
  NAND2_X1 U940 ( .A1(G69), .A2(n846), .ZN(n847) );
  NOR2_X1 U941 ( .A1(G237), .A2(n847), .ZN(n858) );
  NOR2_X1 U942 ( .A1(n848), .A2(n858), .ZN(n849) );
  NOR2_X1 U943 ( .A1(n850), .A2(n849), .ZN(G319) );
  INV_X1 U944 ( .A(G319), .ZN(n852) );
  NAND2_X1 U945 ( .A1(G483), .A2(G661), .ZN(n851) );
  NOR2_X1 U946 ( .A1(n852), .A2(n851), .ZN(n855) );
  NAND2_X1 U947 ( .A1(n855), .A2(G36), .ZN(G176) );
  INV_X1 U948 ( .A(G223), .ZN(n853) );
  NAND2_X1 U949 ( .A1(G2106), .A2(n853), .ZN(G217) );
  AND2_X1 U950 ( .A1(G15), .A2(G2), .ZN(n854) );
  NAND2_X1 U951 ( .A1(G661), .A2(n854), .ZN(G259) );
  NAND2_X1 U952 ( .A1(G1), .A2(G3), .ZN(n856) );
  NAND2_X1 U953 ( .A1(n856), .A2(n855), .ZN(n857) );
  XNOR2_X1 U954 ( .A(n857), .B(KEYINPUT110), .ZN(G188) );
  INV_X1 U955 ( .A(n858), .ZN(n859) );
  NOR2_X1 U956 ( .A1(n860), .A2(n859), .ZN(G325) );
  XNOR2_X1 U957 ( .A(KEYINPUT111), .B(G325), .ZN(G261) );
  NAND2_X1 U959 ( .A1(n862), .A2(n861), .ZN(n864) );
  XNOR2_X1 U960 ( .A(n864), .B(n863), .ZN(G145) );
  INV_X1 U961 ( .A(G96), .ZN(G221) );
  XNOR2_X1 U962 ( .A(G1961), .B(KEYINPUT41), .ZN(n874) );
  XOR2_X1 U963 ( .A(G1956), .B(G1966), .Z(n866) );
  XNOR2_X1 U964 ( .A(G1986), .B(G1981), .ZN(n865) );
  XNOR2_X1 U965 ( .A(n866), .B(n865), .ZN(n870) );
  XOR2_X1 U966 ( .A(G1971), .B(G1976), .Z(n868) );
  XNOR2_X1 U967 ( .A(G1996), .B(G1991), .ZN(n867) );
  XNOR2_X1 U968 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U969 ( .A(n870), .B(n869), .Z(n872) );
  XNOR2_X1 U970 ( .A(KEYINPUT114), .B(G2474), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n872), .B(n871), .ZN(n873) );
  XNOR2_X1 U972 ( .A(n874), .B(n873), .ZN(G229) );
  XOR2_X1 U973 ( .A(G2100), .B(KEYINPUT42), .Z(n876) );
  XNOR2_X1 U974 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n875) );
  XNOR2_X1 U975 ( .A(n876), .B(n875), .ZN(n880) );
  XOR2_X1 U976 ( .A(KEYINPUT43), .B(G2090), .Z(n878) );
  XNOR2_X1 U977 ( .A(G2067), .B(G2072), .ZN(n877) );
  XNOR2_X1 U978 ( .A(n878), .B(n877), .ZN(n879) );
  XOR2_X1 U979 ( .A(n880), .B(n879), .Z(n882) );
  XNOR2_X1 U980 ( .A(G2678), .B(G2096), .ZN(n881) );
  XNOR2_X1 U981 ( .A(n882), .B(n881), .ZN(n884) );
  XOR2_X1 U982 ( .A(G2084), .B(G2078), .Z(n883) );
  XNOR2_X1 U983 ( .A(n884), .B(n883), .ZN(G227) );
  NAND2_X1 U984 ( .A1(G112), .A2(n912), .ZN(n886) );
  NAND2_X1 U985 ( .A1(G100), .A2(n917), .ZN(n885) );
  NAND2_X1 U986 ( .A1(n886), .A2(n885), .ZN(n891) );
  NAND2_X1 U987 ( .A1(n520), .A2(G124), .ZN(n887) );
  XNOR2_X1 U988 ( .A(n887), .B(KEYINPUT44), .ZN(n889) );
  NAND2_X1 U989 ( .A1(G136), .A2(n918), .ZN(n888) );
  NAND2_X1 U990 ( .A1(n889), .A2(n888), .ZN(n890) );
  NOR2_X1 U991 ( .A1(n891), .A2(n890), .ZN(G162) );
  NAND2_X1 U992 ( .A1(G118), .A2(n912), .ZN(n893) );
  NAND2_X1 U993 ( .A1(G130), .A2(n520), .ZN(n892) );
  NAND2_X1 U994 ( .A1(n893), .A2(n892), .ZN(n899) );
  NAND2_X1 U995 ( .A1(n917), .A2(G106), .ZN(n894) );
  XOR2_X1 U996 ( .A(KEYINPUT115), .B(n894), .Z(n896) );
  NAND2_X1 U997 ( .A1(n918), .A2(G142), .ZN(n895) );
  NAND2_X1 U998 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U999 ( .A(n897), .B(KEYINPUT45), .Z(n898) );
  NOR2_X1 U1000 ( .A1(n899), .A2(n898), .ZN(n901) );
  XNOR2_X1 U1001 ( .A(n901), .B(n900), .ZN(n910) );
  XOR2_X1 U1002 ( .A(KEYINPUT116), .B(KEYINPUT46), .Z(n903) );
  XNOR2_X1 U1003 ( .A(n939), .B(KEYINPUT48), .ZN(n902) );
  XNOR2_X1 U1004 ( .A(n903), .B(n902), .ZN(n905) );
  XOR2_X1 U1005 ( .A(n905), .B(n904), .Z(n908) );
  XOR2_X1 U1006 ( .A(G160), .B(n906), .Z(n907) );
  XNOR2_X1 U1007 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1008 ( .A(n910), .B(n909), .Z(n926) );
  XNOR2_X1 U1009 ( .A(KEYINPUT119), .B(KEYINPUT47), .ZN(n916) );
  NAND2_X1 U1010 ( .A1(n520), .A2(G127), .ZN(n911) );
  XNOR2_X1 U1011 ( .A(n911), .B(KEYINPUT118), .ZN(n914) );
  NAND2_X1 U1012 ( .A1(G115), .A2(n912), .ZN(n913) );
  NAND2_X1 U1013 ( .A1(n914), .A2(n913), .ZN(n915) );
  XNOR2_X1 U1014 ( .A(n916), .B(n915), .ZN(n923) );
  NAND2_X1 U1015 ( .A1(G103), .A2(n917), .ZN(n920) );
  NAND2_X1 U1016 ( .A1(G139), .A2(n918), .ZN(n919) );
  NAND2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1018 ( .A(KEYINPUT117), .B(n921), .Z(n922) );
  NOR2_X1 U1019 ( .A1(n923), .A2(n922), .ZN(n950) );
  XNOR2_X1 U1020 ( .A(n950), .B(G162), .ZN(n924) );
  XNOR2_X1 U1021 ( .A(n924), .B(G164), .ZN(n925) );
  XOR2_X1 U1022 ( .A(n926), .B(n925), .Z(n927) );
  NOR2_X1 U1023 ( .A1(G37), .A2(n927), .ZN(G395) );
  XNOR2_X1 U1024 ( .A(n988), .B(n989), .ZN(n929) );
  XNOR2_X1 U1025 ( .A(n929), .B(n928), .ZN(n930) );
  XNOR2_X1 U1026 ( .A(n930), .B(G171), .ZN(n931) );
  XNOR2_X1 U1027 ( .A(n931), .B(G286), .ZN(n932) );
  NOR2_X1 U1028 ( .A1(G37), .A2(n932), .ZN(G397) );
  NOR2_X1 U1029 ( .A1(G229), .A2(G227), .ZN(n933) );
  XNOR2_X1 U1030 ( .A(KEYINPUT49), .B(n933), .ZN(n934) );
  NOR2_X1 U1031 ( .A1(G401), .A2(n934), .ZN(n935) );
  AND2_X1 U1032 ( .A1(G319), .A2(n935), .ZN(n937) );
  NOR2_X1 U1033 ( .A1(G395), .A2(G397), .ZN(n936) );
  NAND2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(G225) );
  INV_X1 U1035 ( .A(G225), .ZN(G308) );
  INV_X1 U1036 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1037 ( .A(G160), .B(G2084), .ZN(n938) );
  XNOR2_X1 U1038 ( .A(n938), .B(KEYINPUT120), .ZN(n942) );
  NOR2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1041 ( .A(KEYINPUT121), .B(n943), .ZN(n949) );
  NAND2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1044 ( .A1(n949), .A2(n948), .ZN(n960) );
  XOR2_X1 U1045 ( .A(G2072), .B(n950), .Z(n952) );
  XOR2_X1 U1046 ( .A(G164), .B(G2078), .Z(n951) );
  NOR2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1048 ( .A(KEYINPUT50), .B(n953), .ZN(n958) );
  XOR2_X1 U1049 ( .A(G2090), .B(G162), .Z(n954) );
  NOR2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n956) );
  XOR2_X1 U1051 ( .A(KEYINPUT51), .B(n956), .Z(n957) );
  NAND2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1054 ( .A(KEYINPUT52), .B(n961), .ZN(n962) );
  XOR2_X1 U1055 ( .A(KEYINPUT55), .B(KEYINPUT122), .Z(n984) );
  NAND2_X1 U1056 ( .A1(n962), .A2(n984), .ZN(n963) );
  NAND2_X1 U1057 ( .A1(n963), .A2(G29), .ZN(n964) );
  XOR2_X1 U1058 ( .A(KEYINPUT123), .B(n964), .Z(n1042) );
  XNOR2_X1 U1059 ( .A(G2067), .B(G26), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(G33), .B(G2072), .ZN(n965) );
  NOR2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n976) );
  XNOR2_X1 U1062 ( .A(G25), .B(n967), .ZN(n968) );
  NAND2_X1 U1063 ( .A1(n968), .A2(G28), .ZN(n974) );
  XNOR2_X1 U1064 ( .A(n969), .B(G27), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(n970), .B(G32), .ZN(n971) );
  NAND2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n973) );
  NOR2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1069 ( .A(n977), .B(KEYINPUT53), .ZN(n980) );
  XOR2_X1 U1070 ( .A(G2084), .B(KEYINPUT54), .Z(n978) );
  XNOR2_X1 U1071 ( .A(G34), .B(n978), .ZN(n979) );
  NAND2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(G35), .B(G2090), .ZN(n981) );
  NOR2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n983) );
  XOR2_X1 U1075 ( .A(n984), .B(n983), .Z(n986) );
  INV_X1 U1076 ( .A(G29), .ZN(n985) );
  NAND2_X1 U1077 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1078 ( .A1(n987), .A2(G11), .ZN(n1040) );
  XNOR2_X1 U1079 ( .A(G16), .B(KEYINPUT56), .ZN(n1012) );
  XOR2_X1 U1080 ( .A(G1348), .B(n988), .Z(n991) );
  XNOR2_X1 U1081 ( .A(n989), .B(G1341), .ZN(n990) );
  NOR2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n998) );
  XOR2_X1 U1083 ( .A(G171), .B(G1961), .Z(n996) );
  XOR2_X1 U1084 ( .A(G1966), .B(G168), .Z(n992) );
  NOR2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1086 ( .A(KEYINPUT57), .B(n994), .ZN(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n1009) );
  XNOR2_X1 U1089 ( .A(G1971), .B(G303), .ZN(n999) );
  NOR2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1002) );
  NAND2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  XNOR2_X1 U1092 ( .A(G1956), .B(G299), .ZN(n1003) );
  NOR2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1006) );
  NAND2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(KEYINPUT124), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(KEYINPUT125), .B(n1010), .ZN(n1011) );
  NAND2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1038) );
  INV_X1 U1099 ( .A(G16), .ZN(n1036) );
  XNOR2_X1 U1100 ( .A(G1348), .B(KEYINPUT59), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(n1013), .B(G4), .ZN(n1017) );
  XNOR2_X1 U1102 ( .A(G1981), .B(G6), .ZN(n1015) );
  XNOR2_X1 U1103 ( .A(G1341), .B(G19), .ZN(n1014) );
  NOR2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1019) );
  XNOR2_X1 U1106 ( .A(G20), .B(G1956), .ZN(n1018) );
  NOR2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1108 ( .A(KEYINPUT60), .B(n1020), .ZN(n1023) );
  XNOR2_X1 U1109 ( .A(n1021), .B(G5), .ZN(n1022) );
  NAND2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1025) );
  XNOR2_X1 U1111 ( .A(G21), .B(G1966), .ZN(n1024) );
  NOR2_X1 U1112 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1113 ( .A(KEYINPUT126), .B(n1026), .Z(n1033) );
  XOR2_X1 U1114 ( .A(G1976), .B(G23), .Z(n1028) );
  XOR2_X1 U1115 ( .A(G1971), .B(G22), .Z(n1027) );
  NAND2_X1 U1116 ( .A1(n1028), .A2(n1027), .ZN(n1030) );
  XNOR2_X1 U1117 ( .A(G24), .B(G1986), .ZN(n1029) );
  NOR2_X1 U1118 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1119 ( .A(KEYINPUT58), .B(n1031), .Z(n1032) );
  NOR2_X1 U1120 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XNOR2_X1 U1121 ( .A(KEYINPUT61), .B(n1034), .ZN(n1035) );
  NAND2_X1 U1122 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NAND2_X1 U1123 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  NOR2_X1 U1124 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  NAND2_X1 U1125 ( .A1(n1042), .A2(n1041), .ZN(n1043) );
  XNOR2_X1 U1126 ( .A(n1043), .B(KEYINPUT127), .ZN(n1044) );
  XNOR2_X1 U1127 ( .A(KEYINPUT62), .B(n1044), .ZN(G311) );
  INV_X1 U1128 ( .A(G311), .ZN(G150) );
endmodule

